VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_rom_krom
   CLASS BLOCK ;
   SIZE 84.33 BY 87.06 ;
   SYMMETRY X Y R90 ;
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 6.83 -7.1 7.21 ;
      END
   END clk0
   PIN cs0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  15.895 -7.48 16.275 -7.1 ;
      END
   END cs0
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  19.71 -7.48 20.09 -7.1 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  21.75 -7.48 22.13 -7.1 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 23.69 -7.1 24.07 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 24.435 -7.1 24.815 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 25.125 -7.1 25.505 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 22.22 -7.1 22.6 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 25.815 -7.1 26.195 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 21.53 -7.1 21.91 ;
      END
   END addr0[7]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  49.105 -7.48 49.485 -7.1 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  52.285 -7.48 52.665 -7.1 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  53.715 -7.48 54.095 -7.1 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  55.255 -7.48 55.635 -7.1 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  56.795 -7.48 57.175 -7.1 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  58.335 -7.48 58.715 -7.1 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  59.875 -7.48 60.255 -7.1 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  61.415 -7.48 61.795 -7.1 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  62.955 -7.48 63.335 -7.1 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  64.495 -7.48 64.875 -7.1 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  66.035 -7.48 66.415 -7.1 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  67.575 -7.48 67.955 -7.1 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  69.86 -7.48 70.24 -7.1 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  71.52 -7.48 71.9 -7.1 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  72.21 -7.48 72.59 -7.1 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  72.9 -7.48 73.28 -7.1 ;
      END
   END dout0[15]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  -7.48 92.8 91.81 94.54 ;
         LAYER met4 ;
         RECT  -7.48 -7.48 -5.74 94.54 ;
         LAYER met3 ;
         RECT  -7.48 -7.48 91.81 -5.74 ;
         LAYER met4 ;
         RECT  90.07 -7.48 91.81 94.54 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  -4.0 -4.0 -2.26 91.06 ;
         LAYER met4 ;
         RECT  86.59 -4.0 88.33 91.06 ;
         LAYER met3 ;
         RECT  -4.0 -4.0 88.33 -2.26 ;
         LAYER met3 ;
         RECT  -4.0 89.32 88.33 91.06 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 83.71 86.44 ;
   LAYER  met2 ;
      RECT  0.62 0.62 83.71 86.44 ;
   LAYER  met3 ;
      RECT  0.62 0.62 83.71 86.44 ;
   LAYER  met4 ;
      RECT  0.62 0.62 83.71 86.44 ;
   END
END    sky130_rom_krom
END    LIBRARY
