magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1296 -1277 1988 3436
<< nwell >>
rect -36 1017 728 2176
<< pwell >>
rect 28 159 554 329
rect 28 25 658 159
<< scnmos >>
rect 114 51 144 303
rect 222 51 252 303
rect 330 51 360 303
rect 438 51 468 303
<< scpmos >>
rect 114 1668 144 2068
rect 222 1668 252 2068
rect 330 1668 360 2068
rect 438 1668 468 2068
<< ndiff >>
rect 54 194 114 303
rect 54 160 62 194
rect 96 160 114 194
rect 54 51 114 160
rect 144 194 222 303
rect 144 160 166 194
rect 200 160 222 194
rect 144 51 222 160
rect 252 194 330 303
rect 252 160 274 194
rect 308 160 330 194
rect 252 51 330 160
rect 360 194 438 303
rect 360 160 382 194
rect 416 160 438 194
rect 360 51 438 160
rect 468 194 528 303
rect 468 160 486 194
rect 520 160 528 194
rect 468 51 528 160
<< pdiff >>
rect 54 1885 114 2068
rect 54 1851 62 1885
rect 96 1851 114 1885
rect 54 1668 114 1851
rect 144 1885 222 2068
rect 144 1851 166 1885
rect 200 1851 222 1885
rect 144 1668 222 1851
rect 252 1885 330 2068
rect 252 1851 274 1885
rect 308 1851 330 1885
rect 252 1668 330 1851
rect 360 1885 438 2068
rect 360 1851 382 1885
rect 416 1851 438 1885
rect 360 1668 438 1851
rect 468 1885 528 2068
rect 468 1851 486 1885
rect 520 1851 528 1885
rect 468 1668 528 1851
<< ndiffc >>
rect 62 160 96 194
rect 166 160 200 194
rect 274 160 308 194
rect 382 160 416 194
rect 486 160 520 194
<< pdiffc >>
rect 62 1851 96 1885
rect 166 1851 200 1885
rect 274 1851 308 1885
rect 382 1851 416 1885
rect 486 1851 520 1885
<< psubdiff >>
rect 582 109 632 133
rect 582 75 590 109
rect 624 75 632 109
rect 582 51 632 75
<< nsubdiff >>
rect 582 2031 632 2055
rect 582 1997 590 2031
rect 624 1997 632 2031
rect 582 1973 632 1997
<< psubdiffcont >>
rect 590 75 624 109
<< nsubdiffcont >>
rect 590 1997 624 2031
<< poly >>
rect 114 2068 144 2094
rect 222 2068 252 2094
rect 330 2068 360 2094
rect 438 2068 468 2094
rect 114 1642 144 1668
rect 222 1642 252 1668
rect 330 1642 360 1668
rect 438 1642 468 1668
rect 114 1612 468 1642
rect 114 1056 144 1612
rect 48 1040 144 1056
rect 48 1006 64 1040
rect 98 1006 144 1040
rect 48 990 144 1006
rect 114 359 144 990
rect 114 329 468 359
rect 114 303 144 329
rect 222 303 252 329
rect 330 303 360 329
rect 438 303 468 329
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
rect 438 25 468 51
<< polycont >>
rect 64 1006 98 1040
<< locali >>
rect 0 2102 692 2136
rect 62 1885 96 2102
rect 62 1835 96 1851
rect 166 1885 200 1901
rect 166 1801 200 1851
rect 274 1885 308 2102
rect 274 1835 308 1851
rect 382 1885 416 1901
rect 382 1801 416 1851
rect 486 1885 520 2102
rect 590 2031 624 2102
rect 590 1981 624 1997
rect 486 1835 520 1851
rect 166 1767 416 1801
rect 64 1040 98 1056
rect 64 990 98 1006
rect 274 1040 308 1767
rect 274 1006 325 1040
rect 274 278 308 1006
rect 166 244 416 278
rect 62 194 96 210
rect 62 17 96 160
rect 166 194 200 244
rect 166 144 200 160
rect 274 194 308 210
rect 274 17 308 160
rect 382 194 416 244
rect 382 144 416 160
rect 486 194 520 210
rect 486 17 520 160
rect 590 109 624 125
rect 590 17 624 75
rect 0 -17 692 17
<< labels >>
rlabel locali s 81 1023 81 1023 4 A
port 1 nsew
rlabel locali s 308 1023 308 1023 4 Z
port 2 nsew
rlabel locali s 346 0 346 0 4 gnd
port 3 nsew
rlabel locali s 346 2119 346 2119 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 692 1784
<< end >>
