magic
tech sky130A
magscale 1 2
timestamp 1581479693
<< checkpaint >>
rect -1296 -1277 1988 3946
<< nwell >>
rect -36 1262 728 2686
<< pwell >>
rect 28 159 554 477
rect 28 25 658 159
<< scnmos >>
rect 114 51 144 451
rect 222 51 252 451
rect 330 51 360 451
rect 438 51 468 451
<< scpmos >>
rect 114 1978 144 2578
rect 222 1978 252 2578
rect 330 1978 360 2578
rect 438 1978 468 2578
<< ndiff >>
rect 54 268 114 451
rect 54 234 62 268
rect 96 234 114 268
rect 54 51 114 234
rect 144 268 222 451
rect 144 234 166 268
rect 200 234 222 268
rect 144 51 222 234
rect 252 268 330 451
rect 252 234 274 268
rect 308 234 330 268
rect 252 51 330 234
rect 360 268 438 451
rect 360 234 382 268
rect 416 234 438 268
rect 360 51 438 234
rect 468 268 528 451
rect 468 234 486 268
rect 520 234 528 268
rect 468 51 528 234
<< pdiff >>
rect 54 2295 114 2578
rect 54 2261 62 2295
rect 96 2261 114 2295
rect 54 1978 114 2261
rect 144 2295 222 2578
rect 144 2261 166 2295
rect 200 2261 222 2295
rect 144 1978 222 2261
rect 252 2295 330 2578
rect 252 2261 274 2295
rect 308 2261 330 2295
rect 252 1978 330 2261
rect 360 2295 438 2578
rect 360 2261 382 2295
rect 416 2261 438 2295
rect 360 1978 438 2261
rect 468 2295 528 2578
rect 468 2261 486 2295
rect 520 2261 528 2295
rect 468 1978 528 2261
<< ndiffc >>
rect 62 234 96 268
rect 166 234 200 268
rect 274 234 308 268
rect 382 234 416 268
rect 486 234 520 268
<< pdiffc >>
rect 62 2261 96 2295
rect 166 2261 200 2295
rect 274 2261 308 2295
rect 382 2261 416 2295
rect 486 2261 520 2295
<< psubdiff >>
rect 582 109 632 133
rect 582 75 590 109
rect 624 75 632 109
rect 582 51 632 75
<< nsubdiff >>
rect 582 2541 632 2565
rect 582 2507 590 2541
rect 624 2507 632 2541
rect 582 2483 632 2507
<< psubdiffcont >>
rect 590 75 624 109
<< nsubdiffcont >>
rect 590 2507 624 2541
<< poly >>
rect 114 2578 144 2604
rect 222 2578 252 2604
rect 330 2578 360 2604
rect 438 2578 468 2604
rect 114 1952 144 1978
rect 222 1952 252 1978
rect 330 1952 360 1978
rect 438 1952 468 1978
rect 114 1922 468 1952
rect 114 1298 144 1922
rect 48 1282 144 1298
rect 48 1248 64 1282
rect 98 1248 144 1282
rect 48 1232 144 1248
rect 114 507 144 1232
rect 114 477 468 507
rect 114 451 144 477
rect 222 451 252 477
rect 330 451 360 477
rect 438 451 468 477
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
rect 438 25 468 51
<< polycont >>
rect 64 1248 98 1282
<< locali >>
rect 0 2612 692 2646
rect 62 2295 96 2612
rect 62 2245 96 2261
rect 166 2295 200 2311
rect 166 2211 200 2261
rect 274 2295 308 2612
rect 274 2245 308 2261
rect 382 2295 416 2311
rect 382 2211 416 2261
rect 486 2295 520 2612
rect 590 2541 624 2612
rect 590 2491 624 2507
rect 486 2245 520 2261
rect 166 2177 416 2211
rect 64 1282 98 1298
rect 64 1232 98 1248
rect 274 1282 308 2177
rect 274 1248 325 1282
rect 274 352 308 1248
rect 166 318 416 352
rect 62 268 96 284
rect 62 17 96 234
rect 166 268 200 318
rect 166 218 200 234
rect 274 268 308 284
rect 274 17 308 234
rect 382 268 416 318
rect 382 218 416 234
rect 486 268 520 284
rect 486 17 520 234
rect 590 109 624 125
rect 590 17 624 75
rect 0 -17 692 17
<< labels >>
rlabel locali s 81 1265 81 1265 4 A
port 1 nsew
rlabel locali s 308 1265 308 1265 4 Z
port 2 nsew
rlabel locali s 346 0 346 0 4 gnd
port 3 nsew
rlabel locali s 346 2629 346 2629 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 692 2194
<< end >>
