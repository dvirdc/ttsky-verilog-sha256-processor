magic
tech sky130A
magscale 1 2
timestamp 1581582910
<< checkpaint >>
rect -1266 -1344 3325 3572
<< poly >>
rect 0 2164 66 2180
rect 0 2130 16 2164
rect 50 2162 66 2164
rect 1736 2164 1802 2180
rect 1736 2162 1752 2164
rect 50 2132 1752 2162
rect 50 2130 66 2132
rect 0 2114 66 2130
rect 1736 2130 1752 2132
rect 1786 2130 1802 2164
rect 1736 2114 1802 2130
rect 0 1960 66 1976
rect 0 1926 16 1960
rect 50 1958 66 1960
rect 1736 1960 1802 1976
rect 1736 1958 1752 1960
rect 50 1928 1752 1958
rect 50 1926 66 1928
rect 0 1910 66 1926
rect 1736 1926 1752 1928
rect 1786 1926 1802 1960
rect 1736 1910 1802 1926
rect 0 1756 66 1772
rect 0 1722 16 1756
rect 50 1754 66 1756
rect 1736 1756 1802 1772
rect 1736 1754 1752 1756
rect 50 1724 1752 1754
rect 50 1722 66 1724
rect 0 1706 66 1722
rect 1736 1722 1752 1724
rect 1786 1722 1802 1756
rect 1736 1706 1802 1722
rect 0 1552 66 1568
rect 0 1518 16 1552
rect 50 1550 66 1552
rect 1736 1552 1802 1568
rect 1736 1550 1752 1552
rect 50 1520 1752 1550
rect 50 1518 66 1520
rect 0 1502 66 1518
rect 1736 1518 1752 1520
rect 1786 1518 1802 1552
rect 1736 1502 1802 1518
rect 0 1348 66 1364
rect 0 1314 16 1348
rect 50 1346 66 1348
rect 1736 1348 1802 1364
rect 1736 1346 1752 1348
rect 50 1316 1752 1346
rect 50 1314 66 1316
rect 0 1298 66 1314
rect 1736 1314 1752 1316
rect 1786 1314 1802 1348
rect 1736 1298 1802 1314
rect 0 1144 66 1160
rect 0 1110 16 1144
rect 50 1142 66 1144
rect 1736 1144 1802 1160
rect 1736 1142 1752 1144
rect 50 1112 1752 1142
rect 50 1110 66 1112
rect 0 1094 66 1110
rect 1736 1110 1752 1112
rect 1786 1110 1802 1144
rect 1736 1094 1802 1110
rect 0 940 66 956
rect 0 906 16 940
rect 50 938 66 940
rect 1736 940 1802 956
rect 1736 938 1752 940
rect 50 908 1752 938
rect 50 906 66 908
rect 0 890 66 906
rect 1736 906 1752 908
rect 1786 906 1802 940
rect 1736 890 1802 906
<< polycont >>
rect 16 2130 50 2164
rect 1752 2130 1786 2164
rect 16 1926 50 1960
rect 1752 1926 1786 1960
rect 16 1722 50 1756
rect 1752 1722 1786 1756
rect 16 1518 50 1552
rect 1752 1518 1786 1552
rect 16 1314 50 1348
rect 1752 1314 1786 1348
rect 16 1110 50 1144
rect 1752 1110 1786 1144
rect 16 906 50 940
rect 1752 906 1786 940
<< locali >>
rect 16 2164 50 2180
rect 16 2114 50 2130
rect 1752 2164 1786 2180
rect 1752 2114 1786 2130
rect 28 2028 44 2062
rect 78 2028 94 2062
rect 1764 2028 1780 2062
rect 1814 2028 1830 2062
rect 16 1960 50 1976
rect 16 1910 50 1926
rect 1752 1960 1786 1976
rect 1752 1910 1786 1926
rect 28 1824 44 1858
rect 78 1824 94 1858
rect 1764 1824 1780 1858
rect 1814 1824 1830 1858
rect 16 1756 50 1772
rect 16 1706 50 1722
rect 1752 1756 1786 1772
rect 1752 1706 1786 1722
rect 28 1620 44 1654
rect 78 1620 94 1654
rect 1764 1620 1780 1654
rect 1814 1620 1830 1654
rect 16 1552 50 1568
rect 16 1502 50 1518
rect 1752 1552 1786 1568
rect 1752 1502 1786 1518
rect 28 1416 44 1450
rect 78 1416 94 1450
rect 1764 1416 1780 1450
rect 1814 1416 1830 1450
rect 16 1348 50 1364
rect 16 1298 50 1314
rect 1752 1348 1786 1364
rect 1752 1298 1786 1314
rect 28 1212 44 1246
rect 78 1212 94 1246
rect 1764 1212 1780 1246
rect 1814 1212 1830 1246
rect 16 1144 50 1160
rect 16 1094 50 1110
rect 1752 1144 1786 1160
rect 1752 1094 1786 1110
rect 28 1008 44 1042
rect 78 1008 94 1042
rect 1764 1008 1780 1042
rect 1814 1008 1830 1042
rect 16 940 50 956
rect 16 890 50 906
rect 1752 940 1786 956
rect 1752 890 1786 906
<< viali >>
rect 16 2130 50 2164
rect 1752 2130 1786 2164
rect 44 2028 78 2062
rect 1780 2028 1814 2062
rect 16 1926 50 1960
rect 1752 1926 1786 1960
rect 44 1824 78 1858
rect 1780 1824 1814 1858
rect 16 1722 50 1756
rect 1752 1722 1786 1756
rect 44 1620 78 1654
rect 1780 1620 1814 1654
rect 16 1518 50 1552
rect 1752 1518 1786 1552
rect 44 1416 78 1450
rect 1780 1416 1814 1450
rect 16 1314 50 1348
rect 1752 1314 1786 1348
rect 44 1212 78 1246
rect 1780 1212 1814 1246
rect 16 1110 50 1144
rect 1752 1110 1786 1144
rect 44 1008 78 1042
rect 1780 1008 1814 1042
rect 16 906 50 940
rect 1752 906 1786 940
<< metal1 >>
rect 29 2248 35 2300
rect 87 2288 93 2300
rect 1765 2288 1771 2300
rect 87 2260 1771 2288
rect 87 2248 93 2260
rect 1765 2248 1771 2260
rect 1823 2248 1829 2300
rect 8 2173 59 2180
rect 1744 2173 1795 2180
rect 1 2121 7 2173
rect 59 2121 65 2173
rect 1737 2121 1743 2173
rect 1795 2161 1801 2173
rect 1795 2133 2065 2161
rect 1795 2121 1801 2133
rect 8 2114 59 2121
rect 1744 2114 1795 2121
rect 35 2071 87 2077
rect 35 2013 87 2019
rect 1771 2071 1823 2077
rect 1771 2013 1823 2019
rect 8 1969 59 1976
rect 1744 1969 1795 1976
rect 1 1917 7 1969
rect 59 1917 65 1969
rect 1737 1917 1743 1969
rect 1795 1917 1801 1969
rect 8 1910 59 1917
rect 1744 1910 1795 1917
rect 35 1867 87 1873
rect 35 1809 87 1815
rect 1771 1867 1823 1873
rect 1771 1809 1823 1815
rect 8 1765 59 1772
rect 1744 1765 1795 1772
rect 1 1713 7 1765
rect 59 1713 65 1765
rect 1737 1713 1743 1765
rect 1795 1713 1801 1765
rect 8 1706 59 1713
rect 1744 1706 1795 1713
rect 35 1663 87 1669
rect 35 1605 87 1611
rect 1771 1663 1823 1669
rect 1771 1605 1823 1611
rect 8 1561 59 1568
rect 1744 1561 1795 1568
rect 1 1509 7 1561
rect 59 1509 65 1561
rect 1737 1509 1743 1561
rect 1795 1509 1801 1561
rect 8 1502 59 1509
rect 1744 1502 1795 1509
rect 35 1459 87 1465
rect 35 1401 87 1407
rect 1771 1459 1823 1465
rect 1771 1401 1823 1407
rect 8 1357 59 1364
rect 1744 1357 1795 1364
rect 1 1305 7 1357
rect 59 1305 65 1357
rect 1737 1305 1743 1357
rect 1795 1305 1801 1357
rect 8 1298 59 1305
rect 1744 1298 1795 1305
rect 35 1255 87 1261
rect 35 1197 87 1203
rect 1771 1255 1823 1261
rect 1771 1197 1823 1203
rect 8 1153 59 1160
rect 1744 1153 1795 1160
rect 1 1101 7 1153
rect 59 1101 65 1153
rect 1737 1101 1743 1153
rect 1795 1101 1801 1153
rect 8 1094 59 1101
rect 1744 1094 1795 1101
rect 35 1051 87 1057
rect 35 993 87 999
rect 1771 1051 1823 1057
rect 1771 993 1823 999
rect 8 949 59 956
rect 1744 949 1795 956
rect 1 897 7 949
rect 59 897 65 949
rect 1737 897 1743 949
rect 1795 897 1801 949
rect 8 890 59 897
rect 1744 890 1795 897
rect 232 -14 260 873
rect 436 -14 464 873
rect 640 -14 668 873
rect 844 -14 872 873
rect 1048 -14 1076 873
rect 1252 -14 1280 873
rect 1456 -14 1484 873
rect 1660 -14 1688 873
rect 2037 396 2065 2133
rect 1811 368 2065 396
<< via1 >>
rect 35 2248 87 2300
rect 1771 2248 1823 2300
rect 7 2164 59 2173
rect 7 2130 16 2164
rect 16 2130 50 2164
rect 50 2130 59 2164
rect 7 2121 59 2130
rect 1743 2164 1795 2173
rect 1743 2130 1752 2164
rect 1752 2130 1786 2164
rect 1786 2130 1795 2164
rect 1743 2121 1795 2130
rect 35 2062 87 2071
rect 35 2028 44 2062
rect 44 2028 78 2062
rect 78 2028 87 2062
rect 35 2019 87 2028
rect 1771 2062 1823 2071
rect 1771 2028 1780 2062
rect 1780 2028 1814 2062
rect 1814 2028 1823 2062
rect 1771 2019 1823 2028
rect 7 1960 59 1969
rect 7 1926 16 1960
rect 16 1926 50 1960
rect 50 1926 59 1960
rect 7 1917 59 1926
rect 1743 1960 1795 1969
rect 1743 1926 1752 1960
rect 1752 1926 1786 1960
rect 1786 1926 1795 1960
rect 1743 1917 1795 1926
rect 35 1858 87 1867
rect 35 1824 44 1858
rect 44 1824 78 1858
rect 78 1824 87 1858
rect 35 1815 87 1824
rect 1771 1858 1823 1867
rect 1771 1824 1780 1858
rect 1780 1824 1814 1858
rect 1814 1824 1823 1858
rect 1771 1815 1823 1824
rect 7 1756 59 1765
rect 7 1722 16 1756
rect 16 1722 50 1756
rect 50 1722 59 1756
rect 7 1713 59 1722
rect 1743 1756 1795 1765
rect 1743 1722 1752 1756
rect 1752 1722 1786 1756
rect 1786 1722 1795 1756
rect 1743 1713 1795 1722
rect 35 1654 87 1663
rect 35 1620 44 1654
rect 44 1620 78 1654
rect 78 1620 87 1654
rect 35 1611 87 1620
rect 1771 1654 1823 1663
rect 1771 1620 1780 1654
rect 1780 1620 1814 1654
rect 1814 1620 1823 1654
rect 1771 1611 1823 1620
rect 7 1552 59 1561
rect 7 1518 16 1552
rect 16 1518 50 1552
rect 50 1518 59 1552
rect 7 1509 59 1518
rect 1743 1552 1795 1561
rect 1743 1518 1752 1552
rect 1752 1518 1786 1552
rect 1786 1518 1795 1552
rect 1743 1509 1795 1518
rect 35 1450 87 1459
rect 35 1416 44 1450
rect 44 1416 78 1450
rect 78 1416 87 1450
rect 35 1407 87 1416
rect 1771 1450 1823 1459
rect 1771 1416 1780 1450
rect 1780 1416 1814 1450
rect 1814 1416 1823 1450
rect 1771 1407 1823 1416
rect 7 1348 59 1357
rect 7 1314 16 1348
rect 16 1314 50 1348
rect 50 1314 59 1348
rect 7 1305 59 1314
rect 1743 1348 1795 1357
rect 1743 1314 1752 1348
rect 1752 1314 1786 1348
rect 1786 1314 1795 1348
rect 1743 1305 1795 1314
rect 35 1246 87 1255
rect 35 1212 44 1246
rect 44 1212 78 1246
rect 78 1212 87 1246
rect 35 1203 87 1212
rect 1771 1246 1823 1255
rect 1771 1212 1780 1246
rect 1780 1212 1814 1246
rect 1814 1212 1823 1246
rect 1771 1203 1823 1212
rect 7 1144 59 1153
rect 7 1110 16 1144
rect 16 1110 50 1144
rect 50 1110 59 1144
rect 7 1101 59 1110
rect 1743 1144 1795 1153
rect 1743 1110 1752 1144
rect 1752 1110 1786 1144
rect 1786 1110 1795 1144
rect 1743 1101 1795 1110
rect 35 1042 87 1051
rect 35 1008 44 1042
rect 44 1008 78 1042
rect 78 1008 87 1042
rect 35 999 87 1008
rect 1771 1042 1823 1051
rect 1771 1008 1780 1042
rect 1780 1008 1814 1042
rect 1814 1008 1823 1042
rect 1771 999 1823 1008
rect 7 940 59 949
rect 7 906 16 940
rect 16 906 50 940
rect 50 906 59 940
rect 7 897 59 906
rect 1743 940 1795 949
rect 1743 906 1752 940
rect 1752 906 1786 940
rect 1786 906 1795 940
rect 1743 897 1795 906
<< metal2 >>
rect 33 2303 89 2312
rect 33 2238 89 2247
rect 1769 2303 1825 2312
rect 1769 2238 1825 2247
rect 7 2173 59 2179
rect 1 2126 7 2169
rect 1743 2173 1795 2179
rect 59 2161 65 2169
rect 1737 2161 1743 2169
rect 59 2133 1743 2161
rect 59 2126 65 2133
rect 1737 2126 1743 2133
rect 7 2115 59 2121
rect 1795 2126 1801 2169
rect 1743 2115 1795 2121
rect 24 2017 33 2073
rect 89 2017 98 2073
rect 1760 2017 1769 2073
rect 1825 2017 1834 2073
rect 7 1969 59 1975
rect 1 1922 7 1965
rect 1743 1969 1795 1975
rect 59 1957 65 1965
rect 1737 1957 1743 1965
rect 59 1929 1743 1957
rect 59 1922 65 1929
rect 1737 1922 1743 1929
rect 7 1911 59 1917
rect 1795 1922 1801 1965
rect 1743 1911 1795 1917
rect 24 1813 33 1869
rect 89 1813 98 1869
rect 1760 1813 1769 1869
rect 1825 1813 1834 1869
rect 7 1765 59 1771
rect 1 1718 7 1761
rect 1743 1765 1795 1771
rect 59 1753 65 1761
rect 1737 1753 1743 1761
rect 59 1725 1743 1753
rect 59 1718 65 1725
rect 1737 1718 1743 1725
rect 7 1707 59 1713
rect 1795 1718 1801 1761
rect 1743 1707 1795 1713
rect 24 1609 33 1665
rect 89 1609 98 1665
rect 1760 1609 1769 1665
rect 1825 1609 1834 1665
rect 7 1561 59 1567
rect 1 1514 7 1557
rect 1743 1561 1795 1567
rect 59 1549 65 1557
rect 1737 1549 1743 1557
rect 59 1521 1743 1549
rect 59 1514 65 1521
rect 1737 1514 1743 1521
rect 7 1503 59 1509
rect 1795 1514 1801 1557
rect 1743 1503 1795 1509
rect 24 1405 33 1461
rect 89 1405 98 1461
rect 1760 1405 1769 1461
rect 1825 1405 1834 1461
rect 7 1357 59 1363
rect 1 1310 7 1353
rect 1743 1357 1795 1363
rect 59 1345 65 1353
rect 1737 1345 1743 1353
rect 59 1317 1743 1345
rect 59 1310 65 1317
rect 1737 1310 1743 1317
rect 7 1299 59 1305
rect 1795 1310 1801 1353
rect 1743 1299 1795 1305
rect 24 1201 33 1257
rect 89 1201 98 1257
rect 1760 1201 1769 1257
rect 1825 1201 1834 1257
rect 7 1153 59 1159
rect 1 1106 7 1149
rect 1743 1153 1795 1159
rect 59 1141 65 1149
rect 1737 1141 1743 1149
rect 59 1113 1743 1141
rect 59 1106 65 1113
rect 1737 1106 1743 1113
rect 7 1095 59 1101
rect 1795 1106 1801 1149
rect 1743 1095 1795 1101
rect 24 997 33 1053
rect 89 997 98 1053
rect 1760 997 1769 1053
rect 1825 997 1834 1053
rect 7 949 59 955
rect 1 902 7 945
rect 1743 949 1795 955
rect 59 937 65 945
rect 1737 937 1743 945
rect 59 909 1743 937
rect 59 902 65 909
rect 1737 902 1743 909
rect 7 891 59 897
rect 1795 902 1801 945
rect 1743 891 1795 897
rect 61 368 89 396
rect 12 -32 40 32
<< via2 >>
rect 33 2300 89 2303
rect 33 2248 35 2300
rect 35 2248 87 2300
rect 87 2248 89 2300
rect 33 2247 89 2248
rect 1769 2300 1825 2303
rect 1769 2248 1771 2300
rect 1771 2248 1823 2300
rect 1823 2248 1825 2300
rect 1769 2247 1825 2248
rect 33 2071 89 2073
rect 33 2019 35 2071
rect 35 2019 87 2071
rect 87 2019 89 2071
rect 33 2017 89 2019
rect 1769 2071 1825 2073
rect 1769 2019 1771 2071
rect 1771 2019 1823 2071
rect 1823 2019 1825 2071
rect 1769 2017 1825 2019
rect 33 1867 89 1869
rect 33 1815 35 1867
rect 35 1815 87 1867
rect 87 1815 89 1867
rect 33 1813 89 1815
rect 1769 1867 1825 1869
rect 1769 1815 1771 1867
rect 1771 1815 1823 1867
rect 1823 1815 1825 1867
rect 1769 1813 1825 1815
rect 33 1663 89 1665
rect 33 1611 35 1663
rect 35 1611 87 1663
rect 87 1611 89 1663
rect 33 1609 89 1611
rect 1769 1663 1825 1665
rect 1769 1611 1771 1663
rect 1771 1611 1823 1663
rect 1823 1611 1825 1663
rect 1769 1609 1825 1611
rect 33 1459 89 1461
rect 33 1407 35 1459
rect 35 1407 87 1459
rect 87 1407 89 1459
rect 33 1405 89 1407
rect 1769 1459 1825 1461
rect 1769 1407 1771 1459
rect 1771 1407 1823 1459
rect 1823 1407 1825 1459
rect 1769 1405 1825 1407
rect 33 1255 89 1257
rect 33 1203 35 1255
rect 35 1203 87 1255
rect 87 1203 89 1255
rect 33 1201 89 1203
rect 1769 1255 1825 1257
rect 1769 1203 1771 1255
rect 1771 1203 1823 1255
rect 1823 1203 1825 1255
rect 1769 1201 1825 1203
rect 33 1051 89 1053
rect 33 999 35 1051
rect 35 999 87 1051
rect 87 999 89 1051
rect 33 997 89 999
rect 1769 1051 1825 1053
rect 1769 999 1771 1051
rect 1771 999 1823 1051
rect 1823 999 1825 1051
rect 1769 997 1825 999
<< metal3 >>
rect 28 2303 94 2308
rect 28 2247 33 2303
rect 89 2247 94 2303
rect 28 2242 94 2247
rect 1764 2303 1830 2308
rect 1764 2247 1769 2303
rect 1825 2247 1830 2303
rect 1764 2242 1830 2247
rect 31 2078 91 2242
rect 1767 2078 1827 2242
rect 28 2073 94 2078
rect 28 2017 33 2073
rect 89 2017 94 2073
rect 28 2012 94 2017
rect 1764 2073 1830 2078
rect 1764 2017 1769 2073
rect 1825 2017 1830 2073
rect 1764 2012 1830 2017
rect 31 1874 91 2012
rect 1767 1874 1827 2012
rect 28 1869 94 1874
rect 28 1813 33 1869
rect 89 1813 94 1869
rect 28 1808 94 1813
rect 1764 1869 1830 1874
rect 1764 1813 1769 1869
rect 1825 1813 1830 1869
rect 1764 1808 1830 1813
rect 31 1670 91 1808
rect 1767 1670 1827 1808
rect 28 1665 94 1670
rect 28 1609 33 1665
rect 89 1609 94 1665
rect 28 1604 94 1609
rect 1764 1665 1830 1670
rect 1764 1609 1769 1665
rect 1825 1609 1830 1665
rect 1764 1604 1830 1609
rect 31 1466 91 1604
rect 1767 1466 1827 1604
rect 28 1461 94 1466
rect 28 1405 33 1461
rect 89 1405 94 1461
rect 28 1400 94 1405
rect 1764 1461 1830 1466
rect 1764 1405 1769 1461
rect 1825 1405 1830 1461
rect 1764 1400 1830 1405
rect 31 1262 91 1400
rect 1767 1262 1827 1400
rect 28 1257 94 1262
rect 28 1201 33 1257
rect 89 1201 94 1257
rect 28 1196 94 1201
rect 1764 1257 1830 1262
rect 1764 1201 1769 1257
rect 1825 1201 1830 1257
rect 1764 1196 1830 1201
rect 31 1058 91 1196
rect 1767 1058 1827 1196
rect 28 1053 94 1058
rect 28 997 33 1053
rect 89 997 94 1053
rect 28 992 94 997
rect 1764 1053 1830 1058
rect 1764 997 1769 1053
rect 1825 997 1830 1053
rect 1764 992 1830 997
rect 31 978 91 992
rect 1767 978 1827 992
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_0
timestamp 1581582907
transform 1 0 1532 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1
timestamp 1581582907
transform 1 0 1328 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_2
timestamp 1581582907
transform 1 0 1124 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_3
timestamp 1581582907
transform 1 0 920 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_4
timestamp 1581582907
transform 1 0 716 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_5
timestamp 1581582907
transform 1 0 512 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_6
timestamp 1581582907
transform 1 0 308 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_7
timestamp 1581582907
transform 1 0 104 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_8
timestamp 1581582907
transform 1 0 1532 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_9
timestamp 1581582907
transform 1 0 1124 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_10
timestamp 1581582907
transform 1 0 716 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_11
timestamp 1581582907
transform 1 0 308 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_12
timestamp 1581582907
transform 1 0 1328 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_13
timestamp 1581582907
transform 1 0 920 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_14
timestamp 1581582907
transform 1 0 512 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_15
timestamp 1581582907
transform 1 0 104 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_16
timestamp 1581582907
transform 1 0 1532 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_17
timestamp 1581582907
transform 1 0 1328 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_18
timestamp 1581582907
transform 1 0 716 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_19
timestamp 1581582907
transform 1 0 512 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_20
timestamp 1581582907
transform 1 0 1124 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_21
timestamp 1581582907
transform 1 0 920 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_22
timestamp 1581582907
transform 1 0 308 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_23
timestamp 1581582907
transform 1 0 104 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_24
timestamp 1581582907
transform 1 0 1532 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_25
timestamp 1581582907
transform 1 0 1328 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_26
timestamp 1581582907
transform 1 0 1124 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_27
timestamp 1581582907
transform 1 0 920 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_28
timestamp 1581582907
transform 1 0 716 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_29
timestamp 1581582907
transform 1 0 512 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_30
timestamp 1581582907
transform 1 0 308 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_31
timestamp 1581582907
transform 1 0 104 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_0
timestamp 1581582907
transform 1 0 1328 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1
timestamp 1581582907
transform 1 0 920 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_2
timestamp 1581582907
transform 1 0 512 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_3
timestamp 1581582907
transform 1 0 104 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_4
timestamp 1581582907
transform 1 0 1532 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_5
timestamp 1581582907
transform 1 0 1124 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_6
timestamp 1581582907
transform 1 0 716 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_7
timestamp 1581582907
transform 1 0 308 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_8
timestamp 1581582907
transform 1 0 1124 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_9
timestamp 1581582907
transform 1 0 920 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_10
timestamp 1581582907
transform 1 0 308 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_11
timestamp 1581582907
transform 1 0 104 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_12
timestamp 1581582907
transform 1 0 1532 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_13
timestamp 1581582907
transform 1 0 1328 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_14
timestamp 1581582907
transform 1 0 716 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_15
timestamp 1581582907
transform 1 0 512 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_16
timestamp 1581582907
transform 1 0 716 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_17
timestamp 1581582907
transform 1 0 512 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_18
timestamp 1581582907
transform 1 0 308 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_19
timestamp 1581582907
transform 1 0 104 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_20
timestamp 1581582907
transform 1 0 1532 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_21
timestamp 1581582907
transform 1 0 1328 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_22
timestamp 1581582907
transform 1 0 1124 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_23
timestamp 1581582907
transform 1 0 920 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_0
timestamp 1581582910
transform 1 0 1736 0 1 1893
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_1
timestamp 1581582910
transform 1 0 0 0 1 1893
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_2
timestamp 1581582910
transform 1 0 1736 0 1 1689
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_3
timestamp 1581582910
transform 1 0 0 0 1 1689
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_4
timestamp 1581582910
transform 1 0 1736 0 1 1485
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_5
timestamp 1581582910
transform 1 0 0 0 1 1485
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_6
timestamp 1581582910
transform 1 0 1736 0 1 1281
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_7
timestamp 1581582910
transform 1 0 0 0 1 1281
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_8
timestamp 1581582910
transform 1 0 1736 0 1 1077
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_9
timestamp 1581582910
transform 1 0 0 0 1 1077
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_10
timestamp 1581582910
transform 1 0 1736 0 1 873
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_11
timestamp 1581582910
transform 1 0 0 0 1 873
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_2  sky130_rom_krom_rom_poly_tap_2_0
timestamp 1581582910
transform 1 0 1736 0 1 2097
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_2  sky130_rom_krom_rom_poly_tap_2_1
timestamp 1581582910
transform 1 0 0 0 1 2097
box 0 17 66 83
use sky130_rom_krom_rom_precharge_array_0  sky130_rom_krom_rom_precharge_array_0_0
timestamp 1581582910
transform 1 0 0 0 1 128
box 0 -212 1948 408
<< labels >>
rlabel metal2 s 61 368 89 396 4 precharge
port 3 nsew
rlabel metal2 s 19 909 47 937 4 wl_0_0
port 5 nsew
rlabel metal2 s 19 1113 47 1141 4 wl_0_1
port 7 nsew
rlabel metal2 s 19 1317 47 1345 4 wl_0_2
port 9 nsew
rlabel metal2 s 19 1521 47 1549 4 wl_0_3
port 11 nsew
rlabel metal2 s 19 1725 47 1753 4 wl_0_4
port 13 nsew
rlabel metal2 s 19 1929 47 1957 4 wl_0_5
port 15 nsew
rlabel metal1 s 232 -14 260 14 4 bl_0_0
port 17 nsew
rlabel metal1 s 436 -14 464 14 4 bl_0_1
port 19 nsew
rlabel metal1 s 640 -14 668 14 4 bl_0_2
port 21 nsew
rlabel metal1 s 844 -14 872 14 4 bl_0_3
port 23 nsew
rlabel metal1 s 1048 -14 1076 14 4 bl_0_4
port 25 nsew
rlabel metal1 s 1252 -14 1280 14 4 bl_0_5
port 27 nsew
rlabel metal1 s 1456 -14 1484 14 4 bl_0_6
port 29 nsew
rlabel metal1 s 1660 -14 1688 14 4 bl_0_7
port 31 nsew
rlabel metal1 s 2037 368 2065 396 4 precharge_r
port 33 nsew
rlabel metal3 s 1767 978 1827 1038 4 gnd
port 35 nsew
rlabel metal3 s 31 2244 91 2304 4 gnd
port 35 nsew
rlabel metal3 s 31 978 91 1038 4 gnd
port 35 nsew
rlabel metal3 s 1767 2244 1827 2304 4 gnd
port 35 nsew
rlabel metal2 s 12 -32 40 32 4 vdd
port 37 nsew
<< properties >>
string FIXED_BBOX 0 0 2065 870
<< end >>
