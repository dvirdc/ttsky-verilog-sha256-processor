magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1296 -1277 1772 3436
<< nwell >>
rect -36 1017 512 2176
<< pwell >>
rect 28 159 338 225
rect 28 25 442 159
<< scnmos >>
rect 114 51 144 199
rect 222 51 252 199
<< scpmos >>
rect 114 1816 144 2068
rect 222 1816 252 2068
<< ndiff >>
rect 54 142 114 199
rect 54 108 62 142
rect 96 108 114 142
rect 54 51 114 108
rect 144 142 222 199
rect 144 108 166 142
rect 200 108 222 142
rect 144 51 222 108
rect 252 142 312 199
rect 252 108 270 142
rect 304 108 312 142
rect 252 51 312 108
<< pdiff >>
rect 54 1959 114 2068
rect 54 1925 62 1959
rect 96 1925 114 1959
rect 54 1816 114 1925
rect 144 1959 222 2068
rect 144 1925 166 1959
rect 200 1925 222 1959
rect 144 1816 222 1925
rect 252 1959 312 2068
rect 252 1925 270 1959
rect 304 1925 312 1959
rect 252 1816 312 1925
<< ndiffc >>
rect 62 108 96 142
rect 166 108 200 142
rect 270 108 304 142
<< pdiffc >>
rect 62 1925 96 1959
rect 166 1925 200 1959
rect 270 1925 304 1959
<< psubdiff >>
rect 366 109 416 133
rect 366 75 374 109
rect 408 75 416 109
rect 366 51 416 75
<< nsubdiff >>
rect 366 2031 416 2055
rect 366 1997 374 2031
rect 408 1997 416 2031
rect 366 1973 416 1997
<< psubdiffcont >>
rect 374 75 408 109
<< nsubdiffcont >>
rect 374 1997 408 2031
<< poly >>
rect 114 2068 144 2094
rect 222 2068 252 2094
rect 114 1790 144 1816
rect 222 1790 252 1816
rect 114 1760 252 1790
rect 114 1066 144 1760
rect 48 1050 144 1066
rect 48 1016 64 1050
rect 98 1016 144 1050
rect 48 1000 144 1016
rect 114 255 144 1000
rect 114 225 252 255
rect 114 199 144 225
rect 222 199 252 225
rect 114 25 144 51
rect 222 25 252 51
<< polycont >>
rect 64 1016 98 1050
<< locali >>
rect 0 2102 476 2136
rect 62 1959 96 2102
rect 62 1909 96 1925
rect 166 1959 200 1975
rect 64 1050 98 1066
rect 64 1000 98 1016
rect 166 1050 200 1925
rect 270 1959 304 2102
rect 374 2031 408 2102
rect 374 1981 408 1997
rect 270 1909 304 1925
rect 166 1016 217 1050
rect 62 142 96 158
rect 62 17 96 108
rect 166 142 200 1016
rect 166 92 200 108
rect 270 142 304 158
rect 270 17 304 108
rect 374 109 408 125
rect 374 17 408 75
rect 0 -17 476 17
<< labels >>
rlabel locali s 81 1033 81 1033 4 A
port 1 nsew
rlabel locali s 200 1033 200 1033 4 Z
port 2 nsew
rlabel locali s 238 0 238 0 4 gnd
port 3 nsew
rlabel locali s 238 2119 238 2119 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 476 1858
<< end >>
