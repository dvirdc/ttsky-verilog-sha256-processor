magic
tech sky130A
magscale 1 2
timestamp 1581320207
<< checkpaint >>
rect -1296 -1277 1988 3946
<< nwell >>
rect -36 1262 728 2686
<< pwell >>
rect 28 159 554 677
rect 28 25 658 159
<< scnmos >>
rect 114 51 144 651
rect 222 51 252 651
rect 330 51 360 651
rect 438 51 468 651
<< scpmos >>
rect 114 1578 144 2578
rect 222 1578 252 2578
rect 330 1578 360 2578
rect 438 1578 468 2578
<< ndiff >>
rect 54 368 114 651
rect 54 334 62 368
rect 96 334 114 368
rect 54 51 114 334
rect 144 368 222 651
rect 144 334 166 368
rect 200 334 222 368
rect 144 51 222 334
rect 252 368 330 651
rect 252 334 274 368
rect 308 334 330 368
rect 252 51 330 334
rect 360 368 438 651
rect 360 334 382 368
rect 416 334 438 368
rect 360 51 438 334
rect 468 368 528 651
rect 468 334 486 368
rect 520 334 528 368
rect 468 51 528 334
<< pdiff >>
rect 54 2095 114 2578
rect 54 2061 62 2095
rect 96 2061 114 2095
rect 54 1578 114 2061
rect 144 2095 222 2578
rect 144 2061 166 2095
rect 200 2061 222 2095
rect 144 1578 222 2061
rect 252 2095 330 2578
rect 252 2061 274 2095
rect 308 2061 330 2095
rect 252 1578 330 2061
rect 360 2095 438 2578
rect 360 2061 382 2095
rect 416 2061 438 2095
rect 360 1578 438 2061
rect 468 2095 528 2578
rect 468 2061 486 2095
rect 520 2061 528 2095
rect 468 1578 528 2061
<< ndiffc >>
rect 62 334 96 368
rect 166 334 200 368
rect 274 334 308 368
rect 382 334 416 368
rect 486 334 520 368
<< pdiffc >>
rect 62 2061 96 2095
rect 166 2061 200 2095
rect 274 2061 308 2095
rect 382 2061 416 2095
rect 486 2061 520 2095
<< psubdiff >>
rect 582 109 632 133
rect 582 75 590 109
rect 624 75 632 109
rect 582 51 632 75
<< nsubdiff >>
rect 582 2541 632 2565
rect 582 2507 590 2541
rect 624 2507 632 2541
rect 582 2483 632 2507
<< psubdiffcont >>
rect 590 75 624 109
<< nsubdiffcont >>
rect 590 2507 624 2541
<< poly >>
rect 114 2578 144 2604
rect 222 2578 252 2604
rect 330 2578 360 2604
rect 438 2578 468 2604
rect 114 1552 144 1578
rect 222 1552 252 1578
rect 330 1552 360 1578
rect 438 1552 468 1578
rect 114 1522 468 1552
rect 114 1248 144 1522
rect 48 1232 144 1248
rect 48 1198 64 1232
rect 98 1198 144 1232
rect 48 1182 144 1198
rect 114 707 144 1182
rect 114 677 468 707
rect 114 651 144 677
rect 222 651 252 677
rect 330 651 360 677
rect 438 651 468 677
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
rect 438 25 468 51
<< polycont >>
rect 64 1198 98 1232
<< locali >>
rect 0 2612 692 2646
rect 62 2095 96 2612
rect 62 2045 96 2061
rect 166 2095 200 2111
rect 166 2011 200 2061
rect 274 2095 308 2612
rect 274 2045 308 2061
rect 382 2095 416 2111
rect 382 2011 416 2061
rect 486 2095 520 2612
rect 590 2541 624 2612
rect 590 2491 624 2507
rect 486 2045 520 2061
rect 166 1977 416 2011
rect 64 1232 98 1248
rect 64 1182 98 1198
rect 274 1232 308 1977
rect 274 1198 325 1232
rect 274 452 308 1198
rect 166 418 416 452
rect 62 368 96 384
rect 62 17 96 334
rect 166 368 200 418
rect 166 318 200 334
rect 274 368 308 384
rect 274 17 308 334
rect 382 368 416 418
rect 382 318 416 334
rect 486 368 520 384
rect 486 17 520 334
rect 590 109 624 125
rect 590 17 624 75
rect 0 -17 692 17
<< labels >>
rlabel locali s 81 1215 81 1215 4 A
port 1 nsew
rlabel locali s 308 1215 308 1215 4 Z
port 2 nsew
rlabel locali s 346 0 346 0 4 gnd
port 3 nsew
rlabel locali s 346 2629 346 2629 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 692 1994
<< end >>
