magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1296 -1309 4226 5546
<< locali >>
rect 1427 4220 1443 4254
rect 1477 4220 1493 4254
rect 64 3233 98 3249
rect 2409 3211 2443 3245
rect 64 3183 98 3199
rect 1243 2101 1259 2135
rect 1293 2101 1309 2135
rect 2882 1873 2916 1889
rect 2882 1823 2916 1839
rect 64 988 98 1054
rect 2041 1026 2075 1042
rect 2041 976 2075 992
rect 2764 535 2798 551
rect 2764 485 2798 501
rect 2664 237 2698 303
rect 1243 -17 1259 17
rect 1293 -17 1309 17
<< viali >>
rect 1443 4220 1477 4254
rect 64 3199 98 3233
rect 1259 2101 1293 2135
rect 2882 1839 2916 1873
rect 2041 992 2075 1026
rect 2764 501 2798 535
rect 1259 -17 1293 17
<< metal1 >>
rect 1434 4263 1486 4269
rect 1434 4205 1486 4211
rect 52 3233 110 3239
rect 52 3199 64 3233
rect 98 3199 110 3233
rect 52 3193 110 3199
rect 67 3118 95 3193
rect 67 3090 2913 3118
rect 1250 2144 1302 2150
rect 1250 2086 1302 2092
rect 2885 1879 2913 3090
rect 2870 1873 2928 1879
rect 2870 1839 2882 1873
rect 2916 1839 2928 1873
rect 2870 1833 2928 1839
rect 2029 1026 2087 1032
rect 2029 992 2041 1026
rect 2075 992 2087 1026
rect 2029 986 2087 992
rect 2044 532 2072 986
rect 2752 535 2810 541
rect 2752 532 2764 535
rect 2044 504 2764 532
rect 2752 501 2764 504
rect 2798 501 2810 535
rect 2752 495 2810 501
rect 1250 26 1302 32
rect 1250 -32 1302 -26
<< via1 >>
rect 1434 4254 1486 4263
rect 1434 4220 1443 4254
rect 1443 4220 1477 4254
rect 1477 4220 1486 4254
rect 1434 4211 1486 4220
rect 1250 2135 1302 2144
rect 1250 2101 1259 2135
rect 1259 2101 1293 2135
rect 1293 2101 1302 2135
rect 1250 2092 1302 2101
rect 1250 17 1302 26
rect 1250 -17 1259 17
rect 1259 -17 1293 17
rect 1293 -17 1302 17
rect 1250 -26 1302 -17
<< metal2 >>
rect 1423 4209 1432 4265
rect 1488 4209 1497 4265
rect 1239 2090 1248 2146
rect 1304 2090 1313 2146
rect 1239 -28 1248 28
rect 1304 -28 1313 28
<< via2 >>
rect 1432 4263 1488 4265
rect 1432 4211 1434 4263
rect 1434 4211 1486 4263
rect 1486 4211 1488 4263
rect 1432 4209 1488 4211
rect 1248 2144 1304 2146
rect 1248 2092 1250 2144
rect 1250 2092 1302 2144
rect 1302 2092 1304 2144
rect 1248 2090 1304 2092
rect 1248 26 1304 28
rect 1248 -26 1250 26
rect 1250 -26 1302 26
rect 1302 -26 1304 26
rect 1248 -28 1304 -26
<< metal3 >>
rect 1411 4265 1509 4286
rect 1411 4209 1432 4265
rect 1488 4209 1509 4265
rect 1411 4188 1509 4209
rect 1227 2146 1325 2167
rect 1227 2090 1248 2146
rect 1304 2090 1325 2146
rect 1227 2069 1325 2090
rect 1227 28 1325 49
rect 1227 -28 1248 28
rect 1304 -28 1325 28
rect 1227 -49 1325 -28
use sky130_rom_krom_rom_clock_driver  sky130_rom_krom_rom_clock_driver_0
timestamp 1581321264
transform 1 0 0 0 1 0
box -36 -17 2588 2176
use sky130_rom_krom_rom_control_nand  sky130_rom_krom_rom_control_nand_0
timestamp 1581321264
transform 1 0 2552 0 1 0
box -36 -17 414 2176
use sky130_rom_krom_rom_precharge_driver  sky130_rom_krom_rom_precharge_driver_0
timestamp 1581321264
transform 1 0 0 0 -1 4237
box -36 -17 2956 2176
<< labels >>
rlabel locali s 81 1021 81 1021 4 clk_in
port 2 nsew
rlabel locali s 2058 1009 2058 1009 4 clk_out
port 3 nsew
rlabel locali s 2426 3228 2426 3228 4 prechrg
port 4 nsew
rlabel locali s 2681 270 2681 270 4 CS
port 5 nsew
rlabel metal3 s 1227 -49 1325 49 4 gnd
port 7 nsew
rlabel metal3 s 1411 4188 1509 4286 4 gnd
port 7 nsew
rlabel metal3 s 1227 2069 1325 2167 4 vdd
port 9 nsew
<< properties >>
string FIXED_BBOX 1239 -33 1313 0
<< end >>
