magic
tech sky130A
magscale 1 2
timestamp 1581320207
<< checkpaint >>
rect -1260 -878 14367 4321
<< poly >>
rect 87 641 117 2272
rect 291 845 321 2272
rect 495 1049 525 2272
rect 699 1253 729 2272
rect 903 1457 933 2272
rect 1107 1661 1137 2272
rect 1311 1865 1341 2272
rect 1515 2069 1545 2272
rect 1606 2071 1672 2087
rect 1606 2069 1622 2071
rect 1515 2039 1622 2069
rect 1606 2037 1622 2039
rect 1656 2037 1672 2071
rect 1606 2021 1672 2037
rect 1402 1867 1468 1883
rect 1402 1865 1418 1867
rect 1311 1835 1418 1865
rect 1402 1833 1418 1835
rect 1452 1833 1468 1867
rect 1402 1817 1468 1833
rect 1198 1663 1264 1679
rect 1198 1661 1214 1663
rect 1107 1631 1214 1661
rect 1198 1629 1214 1631
rect 1248 1629 1264 1663
rect 1198 1613 1264 1629
rect 994 1459 1060 1475
rect 994 1457 1010 1459
rect 903 1427 1010 1457
rect 994 1425 1010 1427
rect 1044 1425 1060 1459
rect 994 1409 1060 1425
rect 790 1255 856 1271
rect 790 1253 806 1255
rect 699 1223 806 1253
rect 790 1221 806 1223
rect 840 1221 856 1255
rect 790 1205 856 1221
rect 586 1051 652 1067
rect 586 1049 602 1051
rect 495 1019 602 1049
rect 586 1017 602 1019
rect 636 1017 652 1051
rect 586 1001 652 1017
rect 382 847 448 863
rect 382 845 398 847
rect 291 815 398 845
rect 382 813 398 815
rect 432 813 448 847
rect 382 797 448 813
rect 178 643 244 659
rect 178 641 194 643
rect 87 611 194 641
rect 178 609 194 611
rect 228 609 244 643
rect 1719 641 1749 2272
rect 1923 845 1953 2272
rect 2127 1049 2157 2272
rect 2331 1253 2361 2272
rect 2535 1457 2565 2272
rect 2739 1661 2769 2272
rect 2943 1865 2973 2272
rect 3147 2069 3177 2272
rect 3238 2071 3304 2087
rect 3238 2069 3254 2071
rect 3147 2039 3254 2069
rect 3238 2037 3254 2039
rect 3288 2037 3304 2071
rect 3238 2021 3304 2037
rect 3034 1867 3100 1883
rect 3034 1865 3050 1867
rect 2943 1835 3050 1865
rect 3034 1833 3050 1835
rect 3084 1833 3100 1867
rect 3034 1817 3100 1833
rect 2830 1663 2896 1679
rect 2830 1661 2846 1663
rect 2739 1631 2846 1661
rect 2830 1629 2846 1631
rect 2880 1629 2896 1663
rect 2830 1613 2896 1629
rect 2626 1459 2692 1475
rect 2626 1457 2642 1459
rect 2535 1427 2642 1457
rect 2626 1425 2642 1427
rect 2676 1425 2692 1459
rect 2626 1409 2692 1425
rect 2422 1255 2488 1271
rect 2422 1253 2438 1255
rect 2331 1223 2438 1253
rect 2422 1221 2438 1223
rect 2472 1221 2488 1255
rect 2422 1205 2488 1221
rect 2218 1051 2284 1067
rect 2218 1049 2234 1051
rect 2127 1019 2234 1049
rect 2218 1017 2234 1019
rect 2268 1017 2284 1051
rect 2218 1001 2284 1017
rect 2014 847 2080 863
rect 2014 845 2030 847
rect 1923 815 2030 845
rect 2014 813 2030 815
rect 2064 813 2080 847
rect 2014 797 2080 813
rect 1810 643 1876 659
rect 1810 641 1826 643
rect 1719 611 1826 641
rect 178 593 244 609
rect 1810 609 1826 611
rect 1860 609 1876 643
rect 3351 641 3381 2272
rect 3555 845 3585 2272
rect 3759 1049 3789 2272
rect 3963 1253 3993 2272
rect 4167 1457 4197 2272
rect 4371 1661 4401 2272
rect 4575 1865 4605 2272
rect 4779 2069 4809 2272
rect 4870 2071 4936 2087
rect 4870 2069 4886 2071
rect 4779 2039 4886 2069
rect 4870 2037 4886 2039
rect 4920 2037 4936 2071
rect 4870 2021 4936 2037
rect 4666 1867 4732 1883
rect 4666 1865 4682 1867
rect 4575 1835 4682 1865
rect 4666 1833 4682 1835
rect 4716 1833 4732 1867
rect 4666 1817 4732 1833
rect 4462 1663 4528 1679
rect 4462 1661 4478 1663
rect 4371 1631 4478 1661
rect 4462 1629 4478 1631
rect 4512 1629 4528 1663
rect 4462 1613 4528 1629
rect 4258 1459 4324 1475
rect 4258 1457 4274 1459
rect 4167 1427 4274 1457
rect 4258 1425 4274 1427
rect 4308 1425 4324 1459
rect 4258 1409 4324 1425
rect 4054 1255 4120 1271
rect 4054 1253 4070 1255
rect 3963 1223 4070 1253
rect 4054 1221 4070 1223
rect 4104 1221 4120 1255
rect 4054 1205 4120 1221
rect 3850 1051 3916 1067
rect 3850 1049 3866 1051
rect 3759 1019 3866 1049
rect 3850 1017 3866 1019
rect 3900 1017 3916 1051
rect 3850 1001 3916 1017
rect 3646 847 3712 863
rect 3646 845 3662 847
rect 3555 815 3662 845
rect 3646 813 3662 815
rect 3696 813 3712 847
rect 3646 797 3712 813
rect 3442 643 3508 659
rect 3442 641 3458 643
rect 3351 611 3458 641
rect 1810 593 1876 609
rect 3442 609 3458 611
rect 3492 609 3508 643
rect 4983 641 5013 2272
rect 5187 845 5217 2272
rect 5391 1049 5421 2272
rect 5595 1253 5625 2272
rect 5799 1457 5829 2272
rect 6003 1661 6033 2272
rect 6207 1865 6237 2272
rect 6411 2069 6441 2272
rect 6502 2071 6568 2087
rect 6502 2069 6518 2071
rect 6411 2039 6518 2069
rect 6502 2037 6518 2039
rect 6552 2037 6568 2071
rect 6502 2021 6568 2037
rect 6298 1867 6364 1883
rect 6298 1865 6314 1867
rect 6207 1835 6314 1865
rect 6298 1833 6314 1835
rect 6348 1833 6364 1867
rect 6298 1817 6364 1833
rect 6094 1663 6160 1679
rect 6094 1661 6110 1663
rect 6003 1631 6110 1661
rect 6094 1629 6110 1631
rect 6144 1629 6160 1663
rect 6094 1613 6160 1629
rect 5890 1459 5956 1475
rect 5890 1457 5906 1459
rect 5799 1427 5906 1457
rect 5890 1425 5906 1427
rect 5940 1425 5956 1459
rect 5890 1409 5956 1425
rect 5686 1255 5752 1271
rect 5686 1253 5702 1255
rect 5595 1223 5702 1253
rect 5686 1221 5702 1223
rect 5736 1221 5752 1255
rect 5686 1205 5752 1221
rect 5482 1051 5548 1067
rect 5482 1049 5498 1051
rect 5391 1019 5498 1049
rect 5482 1017 5498 1019
rect 5532 1017 5548 1051
rect 5482 1001 5548 1017
rect 5278 847 5344 863
rect 5278 845 5294 847
rect 5187 815 5294 845
rect 5278 813 5294 815
rect 5328 813 5344 847
rect 5278 797 5344 813
rect 5074 643 5140 659
rect 5074 641 5090 643
rect 4983 611 5090 641
rect 3442 593 3508 609
rect 5074 609 5090 611
rect 5124 609 5140 643
rect 6615 641 6645 2272
rect 6819 845 6849 2272
rect 7023 1049 7053 2272
rect 7227 1253 7257 2272
rect 7431 1457 7461 2272
rect 7635 1661 7665 2272
rect 7839 1865 7869 2272
rect 8043 2069 8073 2272
rect 8134 2071 8200 2087
rect 8134 2069 8150 2071
rect 8043 2039 8150 2069
rect 8134 2037 8150 2039
rect 8184 2037 8200 2071
rect 8134 2021 8200 2037
rect 7930 1867 7996 1883
rect 7930 1865 7946 1867
rect 7839 1835 7946 1865
rect 7930 1833 7946 1835
rect 7980 1833 7996 1867
rect 7930 1817 7996 1833
rect 7726 1663 7792 1679
rect 7726 1661 7742 1663
rect 7635 1631 7742 1661
rect 7726 1629 7742 1631
rect 7776 1629 7792 1663
rect 7726 1613 7792 1629
rect 7522 1459 7588 1475
rect 7522 1457 7538 1459
rect 7431 1427 7538 1457
rect 7522 1425 7538 1427
rect 7572 1425 7588 1459
rect 7522 1409 7588 1425
rect 7318 1255 7384 1271
rect 7318 1253 7334 1255
rect 7227 1223 7334 1253
rect 7318 1221 7334 1223
rect 7368 1221 7384 1255
rect 7318 1205 7384 1221
rect 7114 1051 7180 1067
rect 7114 1049 7130 1051
rect 7023 1019 7130 1049
rect 7114 1017 7130 1019
rect 7164 1017 7180 1051
rect 7114 1001 7180 1017
rect 6910 847 6976 863
rect 6910 845 6926 847
rect 6819 815 6926 845
rect 6910 813 6926 815
rect 6960 813 6976 847
rect 6910 797 6976 813
rect 6706 643 6772 659
rect 6706 641 6722 643
rect 6615 611 6722 641
rect 5074 593 5140 609
rect 6706 609 6722 611
rect 6756 609 6772 643
rect 8247 641 8277 2272
rect 8451 845 8481 2272
rect 8655 1049 8685 2272
rect 8859 1253 8889 2272
rect 9063 1457 9093 2272
rect 9267 1661 9297 2272
rect 9471 1865 9501 2272
rect 9675 2069 9705 2272
rect 9766 2071 9832 2087
rect 9766 2069 9782 2071
rect 9675 2039 9782 2069
rect 9766 2037 9782 2039
rect 9816 2037 9832 2071
rect 9766 2021 9832 2037
rect 9562 1867 9628 1883
rect 9562 1865 9578 1867
rect 9471 1835 9578 1865
rect 9562 1833 9578 1835
rect 9612 1833 9628 1867
rect 9562 1817 9628 1833
rect 9358 1663 9424 1679
rect 9358 1661 9374 1663
rect 9267 1631 9374 1661
rect 9358 1629 9374 1631
rect 9408 1629 9424 1663
rect 9358 1613 9424 1629
rect 9154 1459 9220 1475
rect 9154 1457 9170 1459
rect 9063 1427 9170 1457
rect 9154 1425 9170 1427
rect 9204 1425 9220 1459
rect 9154 1409 9220 1425
rect 8950 1255 9016 1271
rect 8950 1253 8966 1255
rect 8859 1223 8966 1253
rect 8950 1221 8966 1223
rect 9000 1221 9016 1255
rect 8950 1205 9016 1221
rect 8746 1051 8812 1067
rect 8746 1049 8762 1051
rect 8655 1019 8762 1049
rect 8746 1017 8762 1019
rect 8796 1017 8812 1051
rect 8746 1001 8812 1017
rect 8542 847 8608 863
rect 8542 845 8558 847
rect 8451 815 8558 845
rect 8542 813 8558 815
rect 8592 813 8608 847
rect 8542 797 8608 813
rect 8338 643 8404 659
rect 8338 641 8354 643
rect 8247 611 8354 641
rect 6706 593 6772 609
rect 8338 609 8354 611
rect 8388 609 8404 643
rect 9879 641 9909 2272
rect 10083 845 10113 2272
rect 10287 1049 10317 2272
rect 10491 1253 10521 2272
rect 10695 1457 10725 2272
rect 10899 1661 10929 2272
rect 11103 1865 11133 2272
rect 11307 2069 11337 2272
rect 11398 2071 11464 2087
rect 11398 2069 11414 2071
rect 11307 2039 11414 2069
rect 11398 2037 11414 2039
rect 11448 2037 11464 2071
rect 11398 2021 11464 2037
rect 11194 1867 11260 1883
rect 11194 1865 11210 1867
rect 11103 1835 11210 1865
rect 11194 1833 11210 1835
rect 11244 1833 11260 1867
rect 11194 1817 11260 1833
rect 10990 1663 11056 1679
rect 10990 1661 11006 1663
rect 10899 1631 11006 1661
rect 10990 1629 11006 1631
rect 11040 1629 11056 1663
rect 10990 1613 11056 1629
rect 10786 1459 10852 1475
rect 10786 1457 10802 1459
rect 10695 1427 10802 1457
rect 10786 1425 10802 1427
rect 10836 1425 10852 1459
rect 10786 1409 10852 1425
rect 10582 1255 10648 1271
rect 10582 1253 10598 1255
rect 10491 1223 10598 1253
rect 10582 1221 10598 1223
rect 10632 1221 10648 1255
rect 10582 1205 10648 1221
rect 10378 1051 10444 1067
rect 10378 1049 10394 1051
rect 10287 1019 10394 1049
rect 10378 1017 10394 1019
rect 10428 1017 10444 1051
rect 10378 1001 10444 1017
rect 10174 847 10240 863
rect 10174 845 10190 847
rect 10083 815 10190 845
rect 10174 813 10190 815
rect 10224 813 10240 847
rect 10174 797 10240 813
rect 9970 643 10036 659
rect 9970 641 9986 643
rect 9879 611 9986 641
rect 8338 593 8404 609
rect 9970 609 9986 611
rect 10020 609 10036 643
rect 11511 641 11541 2272
rect 11715 845 11745 2272
rect 11919 1049 11949 2272
rect 12123 1253 12153 2272
rect 12327 1457 12357 2272
rect 12531 1661 12561 2272
rect 12735 1865 12765 2272
rect 12939 2069 12969 2272
rect 13030 2071 13096 2087
rect 13030 2069 13046 2071
rect 12939 2039 13046 2069
rect 13030 2037 13046 2039
rect 13080 2037 13096 2071
rect 13030 2021 13096 2037
rect 12826 1867 12892 1883
rect 12826 1865 12842 1867
rect 12735 1835 12842 1865
rect 12826 1833 12842 1835
rect 12876 1833 12892 1867
rect 12826 1817 12892 1833
rect 12622 1663 12688 1679
rect 12622 1661 12638 1663
rect 12531 1631 12638 1661
rect 12622 1629 12638 1631
rect 12672 1629 12688 1663
rect 12622 1613 12688 1629
rect 12418 1459 12484 1475
rect 12418 1457 12434 1459
rect 12327 1427 12434 1457
rect 12418 1425 12434 1427
rect 12468 1425 12484 1459
rect 12418 1409 12484 1425
rect 12214 1255 12280 1271
rect 12214 1253 12230 1255
rect 12123 1223 12230 1253
rect 12214 1221 12230 1223
rect 12264 1221 12280 1255
rect 12214 1205 12280 1221
rect 12010 1051 12076 1067
rect 12010 1049 12026 1051
rect 11919 1019 12026 1049
rect 12010 1017 12026 1019
rect 12060 1017 12076 1051
rect 12010 1001 12076 1017
rect 11806 847 11872 863
rect 11806 845 11822 847
rect 11715 815 11822 845
rect 11806 813 11822 815
rect 11856 813 11872 847
rect 11806 797 11872 813
rect 11602 643 11668 659
rect 11602 641 11618 643
rect 11511 611 11618 641
rect 9970 593 10036 609
rect 11602 609 11618 611
rect 11652 609 11668 643
rect 11602 593 11668 609
<< polycont >>
rect 1622 2037 1656 2071
rect 1418 1833 1452 1867
rect 1214 1629 1248 1663
rect 1010 1425 1044 1459
rect 806 1221 840 1255
rect 602 1017 636 1051
rect 398 813 432 847
rect 194 609 228 643
rect 3254 2037 3288 2071
rect 3050 1833 3084 1867
rect 2846 1629 2880 1663
rect 2642 1425 2676 1459
rect 2438 1221 2472 1255
rect 2234 1017 2268 1051
rect 2030 813 2064 847
rect 1826 609 1860 643
rect 4886 2037 4920 2071
rect 4682 1833 4716 1867
rect 4478 1629 4512 1663
rect 4274 1425 4308 1459
rect 4070 1221 4104 1255
rect 3866 1017 3900 1051
rect 3662 813 3696 847
rect 3458 609 3492 643
rect 6518 2037 6552 2071
rect 6314 1833 6348 1867
rect 6110 1629 6144 1663
rect 5906 1425 5940 1459
rect 5702 1221 5736 1255
rect 5498 1017 5532 1051
rect 5294 813 5328 847
rect 5090 609 5124 643
rect 8150 2037 8184 2071
rect 7946 1833 7980 1867
rect 7742 1629 7776 1663
rect 7538 1425 7572 1459
rect 7334 1221 7368 1255
rect 7130 1017 7164 1051
rect 6926 813 6960 847
rect 6722 609 6756 643
rect 9782 2037 9816 2071
rect 9578 1833 9612 1867
rect 9374 1629 9408 1663
rect 9170 1425 9204 1459
rect 8966 1221 9000 1255
rect 8762 1017 8796 1051
rect 8558 813 8592 847
rect 8354 609 8388 643
rect 11414 2037 11448 2071
rect 11210 1833 11244 1867
rect 11006 1629 11040 1663
rect 10802 1425 10836 1459
rect 10598 1221 10632 1255
rect 10394 1017 10428 1051
rect 10190 813 10224 847
rect 9986 609 10020 643
rect 13046 2037 13080 2071
rect 12842 1833 12876 1867
rect 12638 1629 12672 1663
rect 12434 1425 12468 1459
rect 12230 1221 12264 1255
rect 12026 1017 12060 1051
rect 11822 813 11856 847
rect 11618 609 11652 643
<< locali >>
rect 1606 2037 1622 2071
rect 1656 2037 1672 2071
rect 3238 2037 3254 2071
rect 3288 2037 3304 2071
rect 4870 2037 4886 2071
rect 4920 2037 4936 2071
rect 6502 2037 6518 2071
rect 6552 2037 6568 2071
rect 8134 2037 8150 2071
rect 8184 2037 8200 2071
rect 9766 2037 9782 2071
rect 9816 2037 9832 2071
rect 11398 2037 11414 2071
rect 11448 2037 11464 2071
rect 13030 2037 13046 2071
rect 13080 2037 13096 2071
rect 1402 1833 1418 1867
rect 1452 1833 1468 1867
rect 3034 1833 3050 1867
rect 3084 1833 3100 1867
rect 4666 1833 4682 1867
rect 4716 1833 4732 1867
rect 6298 1833 6314 1867
rect 6348 1833 6364 1867
rect 7930 1833 7946 1867
rect 7980 1833 7996 1867
rect 9562 1833 9578 1867
rect 9612 1833 9628 1867
rect 11194 1833 11210 1867
rect 11244 1833 11260 1867
rect 12826 1833 12842 1867
rect 12876 1833 12892 1867
rect 1198 1629 1214 1663
rect 1248 1629 1264 1663
rect 2830 1629 2846 1663
rect 2880 1629 2896 1663
rect 4462 1629 4478 1663
rect 4512 1629 4528 1663
rect 6094 1629 6110 1663
rect 6144 1629 6160 1663
rect 7726 1629 7742 1663
rect 7776 1629 7792 1663
rect 9358 1629 9374 1663
rect 9408 1629 9424 1663
rect 10990 1629 11006 1663
rect 11040 1629 11056 1663
rect 12622 1629 12638 1663
rect 12672 1629 12688 1663
rect 994 1425 1010 1459
rect 1044 1425 1060 1459
rect 2626 1425 2642 1459
rect 2676 1425 2692 1459
rect 4258 1425 4274 1459
rect 4308 1425 4324 1459
rect 5890 1425 5906 1459
rect 5940 1425 5956 1459
rect 7522 1425 7538 1459
rect 7572 1425 7588 1459
rect 9154 1425 9170 1459
rect 9204 1425 9220 1459
rect 10786 1425 10802 1459
rect 10836 1425 10852 1459
rect 12418 1425 12434 1459
rect 12468 1425 12484 1459
rect 790 1221 806 1255
rect 840 1221 856 1255
rect 2422 1221 2438 1255
rect 2472 1221 2488 1255
rect 4054 1221 4070 1255
rect 4104 1221 4120 1255
rect 5686 1221 5702 1255
rect 5736 1221 5752 1255
rect 7318 1221 7334 1255
rect 7368 1221 7384 1255
rect 8950 1221 8966 1255
rect 9000 1221 9016 1255
rect 10582 1221 10598 1255
rect 10632 1221 10648 1255
rect 12214 1221 12230 1255
rect 12264 1221 12280 1255
rect 586 1017 602 1051
rect 636 1017 652 1051
rect 2218 1017 2234 1051
rect 2268 1017 2284 1051
rect 3850 1017 3866 1051
rect 3900 1017 3916 1051
rect 5482 1017 5498 1051
rect 5532 1017 5548 1051
rect 7114 1017 7130 1051
rect 7164 1017 7180 1051
rect 8746 1017 8762 1051
rect 8796 1017 8812 1051
rect 10378 1017 10394 1051
rect 10428 1017 10444 1051
rect 12010 1017 12026 1051
rect 12060 1017 12076 1051
rect 382 813 398 847
rect 432 813 448 847
rect 2014 813 2030 847
rect 2064 813 2080 847
rect 3646 813 3662 847
rect 3696 813 3712 847
rect 5278 813 5294 847
rect 5328 813 5344 847
rect 6910 813 6926 847
rect 6960 813 6976 847
rect 8542 813 8558 847
rect 8592 813 8608 847
rect 10174 813 10190 847
rect 10224 813 10240 847
rect 11806 813 11822 847
rect 11856 813 11872 847
rect 178 609 194 643
rect 228 609 244 643
rect 1810 609 1826 643
rect 1860 609 1876 643
rect 3442 609 3458 643
rect 3492 609 3508 643
rect 5074 609 5090 643
rect 5124 609 5140 643
rect 6706 609 6722 643
rect 6756 609 6772 643
rect 8338 609 8354 643
rect 8388 609 8404 643
rect 9970 609 9986 643
rect 10020 609 10036 643
rect 11602 609 11618 643
rect 11652 609 11668 643
<< viali >>
rect 1622 2037 1656 2071
rect 3254 2037 3288 2071
rect 4886 2037 4920 2071
rect 6518 2037 6552 2071
rect 8150 2037 8184 2071
rect 9782 2037 9816 2071
rect 11414 2037 11448 2071
rect 13046 2037 13080 2071
rect 1418 1833 1452 1867
rect 3050 1833 3084 1867
rect 4682 1833 4716 1867
rect 6314 1833 6348 1867
rect 7946 1833 7980 1867
rect 9578 1833 9612 1867
rect 11210 1833 11244 1867
rect 12842 1833 12876 1867
rect 1214 1629 1248 1663
rect 2846 1629 2880 1663
rect 4478 1629 4512 1663
rect 6110 1629 6144 1663
rect 7742 1629 7776 1663
rect 9374 1629 9408 1663
rect 11006 1629 11040 1663
rect 12638 1629 12672 1663
rect 1010 1425 1044 1459
rect 2642 1425 2676 1459
rect 4274 1425 4308 1459
rect 5906 1425 5940 1459
rect 7538 1425 7572 1459
rect 9170 1425 9204 1459
rect 10802 1425 10836 1459
rect 12434 1425 12468 1459
rect 806 1221 840 1255
rect 2438 1221 2472 1255
rect 4070 1221 4104 1255
rect 5702 1221 5736 1255
rect 7334 1221 7368 1255
rect 8966 1221 9000 1255
rect 10598 1221 10632 1255
rect 12230 1221 12264 1255
rect 602 1017 636 1051
rect 2234 1017 2268 1051
rect 3866 1017 3900 1051
rect 5498 1017 5532 1051
rect 7130 1017 7164 1051
rect 8762 1017 8796 1051
rect 10394 1017 10428 1051
rect 12026 1017 12060 1051
rect 398 813 432 847
rect 2030 813 2064 847
rect 3662 813 3696 847
rect 5294 813 5328 847
rect 6926 813 6960 847
rect 8558 813 8592 847
rect 10190 813 10224 847
rect 11822 813 11856 847
rect 194 609 228 643
rect 1826 609 1860 643
rect 3458 609 3492 643
rect 5090 609 5124 643
rect 6722 609 6756 643
rect 8354 609 8388 643
rect 9986 609 10020 643
rect 11618 609 11652 643
<< metal1 >>
rect 80 2874 108 3026
rect 172 2968 178 3020
rect 230 2968 236 3020
rect 284 2874 312 3026
rect 376 2968 382 3020
rect 434 2968 440 3020
rect 488 2874 516 3026
rect 580 2968 586 3020
rect 638 2968 644 3020
rect 692 2874 720 3026
rect 784 2968 790 3020
rect 842 2968 848 3020
rect 896 2874 924 3026
rect 988 2968 994 3020
rect 1046 2968 1052 3020
rect 1100 2874 1128 3026
rect 1192 2968 1198 3020
rect 1250 2968 1256 3020
rect 1304 2874 1332 3026
rect 1396 2968 1402 3020
rect 1454 2968 1460 3020
rect 1508 2874 1536 3026
rect 1600 2968 1606 3020
rect 1658 2968 1664 3020
rect 1712 2874 1740 3026
rect 1804 2968 1810 3020
rect 1862 2968 1868 3020
rect 1916 2874 1944 3026
rect 2008 2968 2014 3020
rect 2066 2968 2072 3020
rect 2120 2874 2148 3026
rect 2212 2968 2218 3020
rect 2270 2968 2276 3020
rect 2324 2874 2352 3026
rect 2416 2968 2422 3020
rect 2474 2968 2480 3020
rect 2528 2874 2556 3026
rect 2620 2968 2626 3020
rect 2678 2968 2684 3020
rect 2732 2874 2760 3026
rect 2824 2968 2830 3020
rect 2882 2968 2888 3020
rect 2936 2874 2964 3026
rect 3028 2968 3034 3020
rect 3086 2968 3092 3020
rect 3140 2874 3168 3026
rect 3232 2968 3238 3020
rect 3290 2968 3296 3020
rect 3344 2874 3372 3026
rect 3436 2968 3442 3020
rect 3494 2968 3500 3020
rect 3548 2874 3576 3026
rect 3640 2968 3646 3020
rect 3698 2968 3704 3020
rect 3752 2874 3780 3026
rect 3844 2968 3850 3020
rect 3902 2968 3908 3020
rect 3956 2874 3984 3026
rect 4048 2968 4054 3020
rect 4106 2968 4112 3020
rect 4160 2874 4188 3026
rect 4252 2968 4258 3020
rect 4310 2968 4316 3020
rect 4364 2874 4392 3026
rect 4456 2968 4462 3020
rect 4514 2968 4520 3020
rect 4568 2874 4596 3026
rect 4660 2968 4666 3020
rect 4718 2968 4724 3020
rect 4772 2874 4800 3026
rect 4864 2968 4870 3020
rect 4922 2968 4928 3020
rect 4976 2874 5004 3026
rect 5068 2968 5074 3020
rect 5126 2968 5132 3020
rect 5180 2874 5208 3026
rect 5272 2968 5278 3020
rect 5330 2968 5336 3020
rect 5384 2874 5412 3026
rect 5476 2968 5482 3020
rect 5534 2968 5540 3020
rect 5588 2874 5616 3026
rect 5680 2968 5686 3020
rect 5738 2968 5744 3020
rect 5792 2874 5820 3026
rect 5884 2968 5890 3020
rect 5942 2968 5948 3020
rect 5996 2874 6024 3026
rect 6088 2968 6094 3020
rect 6146 2968 6152 3020
rect 6200 2874 6228 3026
rect 6292 2968 6298 3020
rect 6350 2968 6356 3020
rect 6404 2874 6432 3026
rect 6496 2968 6502 3020
rect 6554 2968 6560 3020
rect 6608 2874 6636 3026
rect 6700 2968 6706 3020
rect 6758 2968 6764 3020
rect 6812 2874 6840 3026
rect 6904 2968 6910 3020
rect 6962 2968 6968 3020
rect 7016 2874 7044 3026
rect 7108 2968 7114 3020
rect 7166 2968 7172 3020
rect 7220 2874 7248 3026
rect 7312 2968 7318 3020
rect 7370 2968 7376 3020
rect 7424 2874 7452 3026
rect 7516 2968 7522 3020
rect 7574 2968 7580 3020
rect 7628 2874 7656 3026
rect 7720 2968 7726 3020
rect 7778 2968 7784 3020
rect 7832 2874 7860 3026
rect 7924 2968 7930 3020
rect 7982 2968 7988 3020
rect 8036 2874 8064 3026
rect 8128 2968 8134 3020
rect 8186 2968 8192 3020
rect 8240 2874 8268 3026
rect 8332 2968 8338 3020
rect 8390 2968 8396 3020
rect 8444 2874 8472 3026
rect 8536 2968 8542 3020
rect 8594 2968 8600 3020
rect 8648 2874 8676 3026
rect 8740 2968 8746 3020
rect 8798 2968 8804 3020
rect 8852 2874 8880 3026
rect 8944 2968 8950 3020
rect 9002 2968 9008 3020
rect 9056 2874 9084 3026
rect 9148 2968 9154 3020
rect 9206 2968 9212 3020
rect 9260 2874 9288 3026
rect 9352 2968 9358 3020
rect 9410 2968 9416 3020
rect 9464 2874 9492 3026
rect 9556 2968 9562 3020
rect 9614 2968 9620 3020
rect 9668 2874 9696 3026
rect 9760 2968 9766 3020
rect 9818 2968 9824 3020
rect 9872 2874 9900 3026
rect 9964 2968 9970 3020
rect 10022 2968 10028 3020
rect 10076 2874 10104 3026
rect 10168 2968 10174 3020
rect 10226 2968 10232 3020
rect 10280 2874 10308 3026
rect 10372 2968 10378 3020
rect 10430 2968 10436 3020
rect 10484 2874 10512 3026
rect 10576 2968 10582 3020
rect 10634 2968 10640 3020
rect 10688 2874 10716 3026
rect 10780 2968 10786 3020
rect 10838 2968 10844 3020
rect 10892 2874 10920 3026
rect 10984 2968 10990 3020
rect 11042 2968 11048 3020
rect 11096 2874 11124 3026
rect 11188 2968 11194 3020
rect 11246 2968 11252 3020
rect 11300 2874 11328 3026
rect 11392 2968 11398 3020
rect 11450 2968 11456 3020
rect 11504 2874 11532 3026
rect 11596 2968 11602 3020
rect 11654 2968 11660 3020
rect 11708 2874 11736 3026
rect 11800 2968 11806 3020
rect 11858 2968 11864 3020
rect 11912 2874 11940 3026
rect 12004 2968 12010 3020
rect 12062 2968 12068 3020
rect 12116 2874 12144 3026
rect 12208 2968 12214 3020
rect 12266 2968 12272 3020
rect 12320 2874 12348 3026
rect 12412 2968 12418 3020
rect 12470 2968 12476 3020
rect 12524 2874 12552 3026
rect 12616 2968 12622 3020
rect 12674 2968 12680 3020
rect 12728 2874 12756 3026
rect 12820 2968 12826 3020
rect 12878 2968 12884 3020
rect 12932 2874 12960 3026
rect 13024 2968 13030 3020
rect 13082 2968 13088 3020
rect 80 434 108 2244
rect 179 600 185 652
rect 237 600 243 652
rect 284 434 312 2244
rect 383 804 389 856
rect 441 804 447 856
rect 488 434 516 2244
rect 587 1008 593 1060
rect 645 1008 651 1060
rect 692 434 720 2244
rect 791 1212 797 1264
rect 849 1212 855 1264
rect 896 434 924 2244
rect 995 1416 1001 1468
rect 1053 1416 1059 1468
rect 1100 434 1128 2244
rect 1199 1620 1205 1672
rect 1257 1620 1263 1672
rect 1304 434 1332 2244
rect 1403 1824 1409 1876
rect 1461 1824 1467 1876
rect 1508 434 1536 2244
rect 1607 2028 1613 2080
rect 1665 2028 1671 2080
rect 1712 434 1740 2244
rect 1811 600 1817 652
rect 1869 600 1875 652
rect 1916 434 1944 2244
rect 2015 804 2021 856
rect 2073 804 2079 856
rect 2120 434 2148 2244
rect 2219 1008 2225 1060
rect 2277 1008 2283 1060
rect 2324 434 2352 2244
rect 2423 1212 2429 1264
rect 2481 1212 2487 1264
rect 2528 434 2556 2244
rect 2627 1416 2633 1468
rect 2685 1416 2691 1468
rect 2732 434 2760 2244
rect 2831 1620 2837 1672
rect 2889 1620 2895 1672
rect 2936 434 2964 2244
rect 3035 1824 3041 1876
rect 3093 1824 3099 1876
rect 3140 434 3168 2244
rect 3239 2028 3245 2080
rect 3297 2028 3303 2080
rect 3344 434 3372 2244
rect 3443 600 3449 652
rect 3501 600 3507 652
rect 3548 434 3576 2244
rect 3647 804 3653 856
rect 3705 804 3711 856
rect 3752 434 3780 2244
rect 3851 1008 3857 1060
rect 3909 1008 3915 1060
rect 3956 434 3984 2244
rect 4055 1212 4061 1264
rect 4113 1212 4119 1264
rect 4160 434 4188 2244
rect 4259 1416 4265 1468
rect 4317 1416 4323 1468
rect 4364 434 4392 2244
rect 4463 1620 4469 1672
rect 4521 1620 4527 1672
rect 4568 434 4596 2244
rect 4667 1824 4673 1876
rect 4725 1824 4731 1876
rect 4772 434 4800 2244
rect 4871 2028 4877 2080
rect 4929 2028 4935 2080
rect 4976 434 5004 2244
rect 5075 600 5081 652
rect 5133 600 5139 652
rect 5180 434 5208 2244
rect 5279 804 5285 856
rect 5337 804 5343 856
rect 5384 434 5412 2244
rect 5483 1008 5489 1060
rect 5541 1008 5547 1060
rect 5588 434 5616 2244
rect 5687 1212 5693 1264
rect 5745 1212 5751 1264
rect 5792 434 5820 2244
rect 5891 1416 5897 1468
rect 5949 1416 5955 1468
rect 5996 434 6024 2244
rect 6095 1620 6101 1672
rect 6153 1620 6159 1672
rect 6200 434 6228 2244
rect 6299 1824 6305 1876
rect 6357 1824 6363 1876
rect 6404 434 6432 2244
rect 6503 2028 6509 2080
rect 6561 2028 6567 2080
rect 6608 434 6636 2244
rect 6707 600 6713 652
rect 6765 600 6771 652
rect 6812 434 6840 2244
rect 6911 804 6917 856
rect 6969 804 6975 856
rect 7016 434 7044 2244
rect 7115 1008 7121 1060
rect 7173 1008 7179 1060
rect 7220 434 7248 2244
rect 7319 1212 7325 1264
rect 7377 1212 7383 1264
rect 7424 434 7452 2244
rect 7523 1416 7529 1468
rect 7581 1416 7587 1468
rect 7628 434 7656 2244
rect 7727 1620 7733 1672
rect 7785 1620 7791 1672
rect 7832 434 7860 2244
rect 7931 1824 7937 1876
rect 7989 1824 7995 1876
rect 8036 434 8064 2244
rect 8135 2028 8141 2080
rect 8193 2028 8199 2080
rect 8240 434 8268 2244
rect 8339 600 8345 652
rect 8397 600 8403 652
rect 8444 434 8472 2244
rect 8543 804 8549 856
rect 8601 804 8607 856
rect 8648 434 8676 2244
rect 8747 1008 8753 1060
rect 8805 1008 8811 1060
rect 8852 434 8880 2244
rect 8951 1212 8957 1264
rect 9009 1212 9015 1264
rect 9056 434 9084 2244
rect 9155 1416 9161 1468
rect 9213 1416 9219 1468
rect 9260 434 9288 2244
rect 9359 1620 9365 1672
rect 9417 1620 9423 1672
rect 9464 434 9492 2244
rect 9563 1824 9569 1876
rect 9621 1824 9627 1876
rect 9668 434 9696 2244
rect 9767 2028 9773 2080
rect 9825 2028 9831 2080
rect 9872 434 9900 2244
rect 9971 600 9977 652
rect 10029 600 10035 652
rect 10076 434 10104 2244
rect 10175 804 10181 856
rect 10233 804 10239 856
rect 10280 434 10308 2244
rect 10379 1008 10385 1060
rect 10437 1008 10443 1060
rect 10484 434 10512 2244
rect 10583 1212 10589 1264
rect 10641 1212 10647 1264
rect 10688 434 10716 2244
rect 10787 1416 10793 1468
rect 10845 1416 10851 1468
rect 10892 434 10920 2244
rect 10991 1620 10997 1672
rect 11049 1620 11055 1672
rect 11096 434 11124 2244
rect 11195 1824 11201 1876
rect 11253 1824 11259 1876
rect 11300 434 11328 2244
rect 11399 2028 11405 2080
rect 11457 2028 11463 2080
rect 11504 434 11532 2244
rect 11603 600 11609 652
rect 11661 600 11667 652
rect 11708 434 11736 2244
rect 11807 804 11813 856
rect 11865 804 11871 856
rect 11912 434 11940 2244
rect 12011 1008 12017 1060
rect 12069 1008 12075 1060
rect 12116 434 12144 2244
rect 12215 1212 12221 1264
rect 12273 1212 12279 1264
rect 12320 434 12348 2244
rect 12419 1416 12425 1468
rect 12477 1416 12483 1468
rect 12524 434 12552 2244
rect 12623 1620 12629 1672
rect 12681 1620 12687 1672
rect 12728 434 12756 2244
rect 12827 1824 12833 1876
rect 12885 1824 12891 1876
rect 12932 434 12960 2244
rect 13031 2028 13037 2080
rect 13089 2028 13095 2080
rect 62 382 68 434
rect 120 382 126 434
rect 266 382 272 434
rect 324 382 330 434
rect 470 382 476 434
rect 528 382 534 434
rect 674 382 680 434
rect 732 382 738 434
rect 878 382 884 434
rect 936 382 942 434
rect 1082 382 1088 434
rect 1140 382 1146 434
rect 1286 382 1292 434
rect 1344 382 1350 434
rect 1490 382 1496 434
rect 1548 382 1554 434
rect 1694 382 1700 434
rect 1752 382 1758 434
rect 1898 382 1904 434
rect 1956 382 1962 434
rect 2102 382 2108 434
rect 2160 382 2166 434
rect 2306 382 2312 434
rect 2364 382 2370 434
rect 2510 382 2516 434
rect 2568 382 2574 434
rect 2714 382 2720 434
rect 2772 382 2778 434
rect 2918 382 2924 434
rect 2976 382 2982 434
rect 3122 382 3128 434
rect 3180 382 3186 434
rect 3326 382 3332 434
rect 3384 382 3390 434
rect 3530 382 3536 434
rect 3588 382 3594 434
rect 3734 382 3740 434
rect 3792 382 3798 434
rect 3938 382 3944 434
rect 3996 382 4002 434
rect 4142 382 4148 434
rect 4200 382 4206 434
rect 4346 382 4352 434
rect 4404 382 4410 434
rect 4550 382 4556 434
rect 4608 382 4614 434
rect 4754 382 4760 434
rect 4812 382 4818 434
rect 4958 382 4964 434
rect 5016 382 5022 434
rect 5162 382 5168 434
rect 5220 382 5226 434
rect 5366 382 5372 434
rect 5424 382 5430 434
rect 5570 382 5576 434
rect 5628 382 5634 434
rect 5774 382 5780 434
rect 5832 382 5838 434
rect 5978 382 5984 434
rect 6036 382 6042 434
rect 6182 382 6188 434
rect 6240 382 6246 434
rect 6386 382 6392 434
rect 6444 382 6450 434
rect 6590 382 6596 434
rect 6648 382 6654 434
rect 6794 382 6800 434
rect 6852 382 6858 434
rect 6998 382 7004 434
rect 7056 382 7062 434
rect 7202 382 7208 434
rect 7260 382 7266 434
rect 7406 382 7412 434
rect 7464 382 7470 434
rect 7610 382 7616 434
rect 7668 382 7674 434
rect 7814 382 7820 434
rect 7872 382 7878 434
rect 8018 382 8024 434
rect 8076 382 8082 434
rect 8222 382 8228 434
rect 8280 382 8286 434
rect 8426 382 8432 434
rect 8484 382 8490 434
rect 8630 382 8636 434
rect 8688 382 8694 434
rect 8834 382 8840 434
rect 8892 382 8898 434
rect 9038 382 9044 434
rect 9096 382 9102 434
rect 9242 382 9248 434
rect 9300 382 9306 434
rect 9446 382 9452 434
rect 9504 382 9510 434
rect 9650 382 9656 434
rect 9708 382 9714 434
rect 9854 382 9860 434
rect 9912 382 9918 434
rect 10058 382 10064 434
rect 10116 382 10122 434
rect 10262 382 10268 434
rect 10320 382 10326 434
rect 10466 382 10472 434
rect 10524 382 10530 434
rect 10670 382 10676 434
rect 10728 382 10734 434
rect 10874 382 10880 434
rect 10932 382 10938 434
rect 11078 382 11084 434
rect 11136 382 11142 434
rect 11282 382 11288 434
rect 11340 382 11346 434
rect 11486 382 11492 434
rect 11544 382 11550 434
rect 11690 382 11696 434
rect 11748 382 11754 434
rect 11894 382 11900 434
rect 11952 382 11958 434
rect 12098 382 12104 434
rect 12156 382 12162 434
rect 12302 382 12308 434
rect 12360 382 12366 434
rect 12506 382 12512 434
rect 12564 382 12570 434
rect 12710 382 12716 434
rect 12768 382 12774 434
rect 12914 382 12920 434
rect 12972 382 12978 434
<< via1 >>
rect 178 2968 230 3020
rect 382 2968 434 3020
rect 586 2968 638 3020
rect 790 2968 842 3020
rect 994 2968 1046 3020
rect 1198 2968 1250 3020
rect 1402 2968 1454 3020
rect 1606 2968 1658 3020
rect 1810 2968 1862 3020
rect 2014 2968 2066 3020
rect 2218 2968 2270 3020
rect 2422 2968 2474 3020
rect 2626 2968 2678 3020
rect 2830 2968 2882 3020
rect 3034 2968 3086 3020
rect 3238 2968 3290 3020
rect 3442 2968 3494 3020
rect 3646 2968 3698 3020
rect 3850 2968 3902 3020
rect 4054 2968 4106 3020
rect 4258 2968 4310 3020
rect 4462 2968 4514 3020
rect 4666 2968 4718 3020
rect 4870 2968 4922 3020
rect 5074 2968 5126 3020
rect 5278 2968 5330 3020
rect 5482 2968 5534 3020
rect 5686 2968 5738 3020
rect 5890 2968 5942 3020
rect 6094 2968 6146 3020
rect 6298 2968 6350 3020
rect 6502 2968 6554 3020
rect 6706 2968 6758 3020
rect 6910 2968 6962 3020
rect 7114 2968 7166 3020
rect 7318 2968 7370 3020
rect 7522 2968 7574 3020
rect 7726 2968 7778 3020
rect 7930 2968 7982 3020
rect 8134 2968 8186 3020
rect 8338 2968 8390 3020
rect 8542 2968 8594 3020
rect 8746 2968 8798 3020
rect 8950 2968 9002 3020
rect 9154 2968 9206 3020
rect 9358 2968 9410 3020
rect 9562 2968 9614 3020
rect 9766 2968 9818 3020
rect 9970 2968 10022 3020
rect 10174 2968 10226 3020
rect 10378 2968 10430 3020
rect 10582 2968 10634 3020
rect 10786 2968 10838 3020
rect 10990 2968 11042 3020
rect 11194 2968 11246 3020
rect 11398 2968 11450 3020
rect 11602 2968 11654 3020
rect 11806 2968 11858 3020
rect 12010 2968 12062 3020
rect 12214 2968 12266 3020
rect 12418 2968 12470 3020
rect 12622 2968 12674 3020
rect 12826 2968 12878 3020
rect 13030 2968 13082 3020
rect 185 643 237 652
rect 185 609 194 643
rect 194 609 228 643
rect 228 609 237 643
rect 185 600 237 609
rect 389 847 441 856
rect 389 813 398 847
rect 398 813 432 847
rect 432 813 441 847
rect 389 804 441 813
rect 593 1051 645 1060
rect 593 1017 602 1051
rect 602 1017 636 1051
rect 636 1017 645 1051
rect 593 1008 645 1017
rect 797 1255 849 1264
rect 797 1221 806 1255
rect 806 1221 840 1255
rect 840 1221 849 1255
rect 797 1212 849 1221
rect 1001 1459 1053 1468
rect 1001 1425 1010 1459
rect 1010 1425 1044 1459
rect 1044 1425 1053 1459
rect 1001 1416 1053 1425
rect 1205 1663 1257 1672
rect 1205 1629 1214 1663
rect 1214 1629 1248 1663
rect 1248 1629 1257 1663
rect 1205 1620 1257 1629
rect 1409 1867 1461 1876
rect 1409 1833 1418 1867
rect 1418 1833 1452 1867
rect 1452 1833 1461 1867
rect 1409 1824 1461 1833
rect 1613 2071 1665 2080
rect 1613 2037 1622 2071
rect 1622 2037 1656 2071
rect 1656 2037 1665 2071
rect 1613 2028 1665 2037
rect 1817 643 1869 652
rect 1817 609 1826 643
rect 1826 609 1860 643
rect 1860 609 1869 643
rect 1817 600 1869 609
rect 2021 847 2073 856
rect 2021 813 2030 847
rect 2030 813 2064 847
rect 2064 813 2073 847
rect 2021 804 2073 813
rect 2225 1051 2277 1060
rect 2225 1017 2234 1051
rect 2234 1017 2268 1051
rect 2268 1017 2277 1051
rect 2225 1008 2277 1017
rect 2429 1255 2481 1264
rect 2429 1221 2438 1255
rect 2438 1221 2472 1255
rect 2472 1221 2481 1255
rect 2429 1212 2481 1221
rect 2633 1459 2685 1468
rect 2633 1425 2642 1459
rect 2642 1425 2676 1459
rect 2676 1425 2685 1459
rect 2633 1416 2685 1425
rect 2837 1663 2889 1672
rect 2837 1629 2846 1663
rect 2846 1629 2880 1663
rect 2880 1629 2889 1663
rect 2837 1620 2889 1629
rect 3041 1867 3093 1876
rect 3041 1833 3050 1867
rect 3050 1833 3084 1867
rect 3084 1833 3093 1867
rect 3041 1824 3093 1833
rect 3245 2071 3297 2080
rect 3245 2037 3254 2071
rect 3254 2037 3288 2071
rect 3288 2037 3297 2071
rect 3245 2028 3297 2037
rect 3449 643 3501 652
rect 3449 609 3458 643
rect 3458 609 3492 643
rect 3492 609 3501 643
rect 3449 600 3501 609
rect 3653 847 3705 856
rect 3653 813 3662 847
rect 3662 813 3696 847
rect 3696 813 3705 847
rect 3653 804 3705 813
rect 3857 1051 3909 1060
rect 3857 1017 3866 1051
rect 3866 1017 3900 1051
rect 3900 1017 3909 1051
rect 3857 1008 3909 1017
rect 4061 1255 4113 1264
rect 4061 1221 4070 1255
rect 4070 1221 4104 1255
rect 4104 1221 4113 1255
rect 4061 1212 4113 1221
rect 4265 1459 4317 1468
rect 4265 1425 4274 1459
rect 4274 1425 4308 1459
rect 4308 1425 4317 1459
rect 4265 1416 4317 1425
rect 4469 1663 4521 1672
rect 4469 1629 4478 1663
rect 4478 1629 4512 1663
rect 4512 1629 4521 1663
rect 4469 1620 4521 1629
rect 4673 1867 4725 1876
rect 4673 1833 4682 1867
rect 4682 1833 4716 1867
rect 4716 1833 4725 1867
rect 4673 1824 4725 1833
rect 4877 2071 4929 2080
rect 4877 2037 4886 2071
rect 4886 2037 4920 2071
rect 4920 2037 4929 2071
rect 4877 2028 4929 2037
rect 5081 643 5133 652
rect 5081 609 5090 643
rect 5090 609 5124 643
rect 5124 609 5133 643
rect 5081 600 5133 609
rect 5285 847 5337 856
rect 5285 813 5294 847
rect 5294 813 5328 847
rect 5328 813 5337 847
rect 5285 804 5337 813
rect 5489 1051 5541 1060
rect 5489 1017 5498 1051
rect 5498 1017 5532 1051
rect 5532 1017 5541 1051
rect 5489 1008 5541 1017
rect 5693 1255 5745 1264
rect 5693 1221 5702 1255
rect 5702 1221 5736 1255
rect 5736 1221 5745 1255
rect 5693 1212 5745 1221
rect 5897 1459 5949 1468
rect 5897 1425 5906 1459
rect 5906 1425 5940 1459
rect 5940 1425 5949 1459
rect 5897 1416 5949 1425
rect 6101 1663 6153 1672
rect 6101 1629 6110 1663
rect 6110 1629 6144 1663
rect 6144 1629 6153 1663
rect 6101 1620 6153 1629
rect 6305 1867 6357 1876
rect 6305 1833 6314 1867
rect 6314 1833 6348 1867
rect 6348 1833 6357 1867
rect 6305 1824 6357 1833
rect 6509 2071 6561 2080
rect 6509 2037 6518 2071
rect 6518 2037 6552 2071
rect 6552 2037 6561 2071
rect 6509 2028 6561 2037
rect 6713 643 6765 652
rect 6713 609 6722 643
rect 6722 609 6756 643
rect 6756 609 6765 643
rect 6713 600 6765 609
rect 6917 847 6969 856
rect 6917 813 6926 847
rect 6926 813 6960 847
rect 6960 813 6969 847
rect 6917 804 6969 813
rect 7121 1051 7173 1060
rect 7121 1017 7130 1051
rect 7130 1017 7164 1051
rect 7164 1017 7173 1051
rect 7121 1008 7173 1017
rect 7325 1255 7377 1264
rect 7325 1221 7334 1255
rect 7334 1221 7368 1255
rect 7368 1221 7377 1255
rect 7325 1212 7377 1221
rect 7529 1459 7581 1468
rect 7529 1425 7538 1459
rect 7538 1425 7572 1459
rect 7572 1425 7581 1459
rect 7529 1416 7581 1425
rect 7733 1663 7785 1672
rect 7733 1629 7742 1663
rect 7742 1629 7776 1663
rect 7776 1629 7785 1663
rect 7733 1620 7785 1629
rect 7937 1867 7989 1876
rect 7937 1833 7946 1867
rect 7946 1833 7980 1867
rect 7980 1833 7989 1867
rect 7937 1824 7989 1833
rect 8141 2071 8193 2080
rect 8141 2037 8150 2071
rect 8150 2037 8184 2071
rect 8184 2037 8193 2071
rect 8141 2028 8193 2037
rect 8345 643 8397 652
rect 8345 609 8354 643
rect 8354 609 8388 643
rect 8388 609 8397 643
rect 8345 600 8397 609
rect 8549 847 8601 856
rect 8549 813 8558 847
rect 8558 813 8592 847
rect 8592 813 8601 847
rect 8549 804 8601 813
rect 8753 1051 8805 1060
rect 8753 1017 8762 1051
rect 8762 1017 8796 1051
rect 8796 1017 8805 1051
rect 8753 1008 8805 1017
rect 8957 1255 9009 1264
rect 8957 1221 8966 1255
rect 8966 1221 9000 1255
rect 9000 1221 9009 1255
rect 8957 1212 9009 1221
rect 9161 1459 9213 1468
rect 9161 1425 9170 1459
rect 9170 1425 9204 1459
rect 9204 1425 9213 1459
rect 9161 1416 9213 1425
rect 9365 1663 9417 1672
rect 9365 1629 9374 1663
rect 9374 1629 9408 1663
rect 9408 1629 9417 1663
rect 9365 1620 9417 1629
rect 9569 1867 9621 1876
rect 9569 1833 9578 1867
rect 9578 1833 9612 1867
rect 9612 1833 9621 1867
rect 9569 1824 9621 1833
rect 9773 2071 9825 2080
rect 9773 2037 9782 2071
rect 9782 2037 9816 2071
rect 9816 2037 9825 2071
rect 9773 2028 9825 2037
rect 9977 643 10029 652
rect 9977 609 9986 643
rect 9986 609 10020 643
rect 10020 609 10029 643
rect 9977 600 10029 609
rect 10181 847 10233 856
rect 10181 813 10190 847
rect 10190 813 10224 847
rect 10224 813 10233 847
rect 10181 804 10233 813
rect 10385 1051 10437 1060
rect 10385 1017 10394 1051
rect 10394 1017 10428 1051
rect 10428 1017 10437 1051
rect 10385 1008 10437 1017
rect 10589 1255 10641 1264
rect 10589 1221 10598 1255
rect 10598 1221 10632 1255
rect 10632 1221 10641 1255
rect 10589 1212 10641 1221
rect 10793 1459 10845 1468
rect 10793 1425 10802 1459
rect 10802 1425 10836 1459
rect 10836 1425 10845 1459
rect 10793 1416 10845 1425
rect 10997 1663 11049 1672
rect 10997 1629 11006 1663
rect 11006 1629 11040 1663
rect 11040 1629 11049 1663
rect 10997 1620 11049 1629
rect 11201 1867 11253 1876
rect 11201 1833 11210 1867
rect 11210 1833 11244 1867
rect 11244 1833 11253 1867
rect 11201 1824 11253 1833
rect 11405 2071 11457 2080
rect 11405 2037 11414 2071
rect 11414 2037 11448 2071
rect 11448 2037 11457 2071
rect 11405 2028 11457 2037
rect 11609 643 11661 652
rect 11609 609 11618 643
rect 11618 609 11652 643
rect 11652 609 11661 643
rect 11609 600 11661 609
rect 11813 847 11865 856
rect 11813 813 11822 847
rect 11822 813 11856 847
rect 11856 813 11865 847
rect 11813 804 11865 813
rect 12017 1051 12069 1060
rect 12017 1017 12026 1051
rect 12026 1017 12060 1051
rect 12060 1017 12069 1051
rect 12017 1008 12069 1017
rect 12221 1255 12273 1264
rect 12221 1221 12230 1255
rect 12230 1221 12264 1255
rect 12264 1221 12273 1255
rect 12221 1212 12273 1221
rect 12425 1459 12477 1468
rect 12425 1425 12434 1459
rect 12434 1425 12468 1459
rect 12468 1425 12477 1459
rect 12425 1416 12477 1425
rect 12629 1663 12681 1672
rect 12629 1629 12638 1663
rect 12638 1629 12672 1663
rect 12672 1629 12681 1663
rect 12629 1620 12681 1629
rect 12833 1867 12885 1876
rect 12833 1833 12842 1867
rect 12842 1833 12876 1867
rect 12876 1833 12885 1867
rect 12833 1824 12885 1833
rect 13037 2071 13089 2080
rect 13037 2037 13046 2071
rect 13046 2037 13080 2071
rect 13080 2037 13089 2071
rect 13037 2028 13089 2037
rect 68 382 120 434
rect 272 382 324 434
rect 476 382 528 434
rect 680 382 732 434
rect 884 382 936 434
rect 1088 382 1140 434
rect 1292 382 1344 434
rect 1496 382 1548 434
rect 1700 382 1752 434
rect 1904 382 1956 434
rect 2108 382 2160 434
rect 2312 382 2364 434
rect 2516 382 2568 434
rect 2720 382 2772 434
rect 2924 382 2976 434
rect 3128 382 3180 434
rect 3332 382 3384 434
rect 3536 382 3588 434
rect 3740 382 3792 434
rect 3944 382 3996 434
rect 4148 382 4200 434
rect 4352 382 4404 434
rect 4556 382 4608 434
rect 4760 382 4812 434
rect 4964 382 5016 434
rect 5168 382 5220 434
rect 5372 382 5424 434
rect 5576 382 5628 434
rect 5780 382 5832 434
rect 5984 382 6036 434
rect 6188 382 6240 434
rect 6392 382 6444 434
rect 6596 382 6648 434
rect 6800 382 6852 434
rect 7004 382 7056 434
rect 7208 382 7260 434
rect 7412 382 7464 434
rect 7616 382 7668 434
rect 7820 382 7872 434
rect 8024 382 8076 434
rect 8228 382 8280 434
rect 8432 382 8484 434
rect 8636 382 8688 434
rect 8840 382 8892 434
rect 9044 382 9096 434
rect 9248 382 9300 434
rect 9452 382 9504 434
rect 9656 382 9708 434
rect 9860 382 9912 434
rect 10064 382 10116 434
rect 10268 382 10320 434
rect 10472 382 10524 434
rect 10676 382 10728 434
rect 10880 382 10932 434
rect 11084 382 11136 434
rect 11288 382 11340 434
rect 11492 382 11544 434
rect 11696 382 11748 434
rect 11900 382 11952 434
rect 12104 382 12156 434
rect 12308 382 12360 434
rect 12512 382 12564 434
rect 12716 382 12768 434
rect 12920 382 12972 434
<< metal2 >>
rect 26 3020 13096 3026
rect 26 2968 178 3020
rect 230 2968 382 3020
rect 434 2968 586 3020
rect 638 2968 790 3020
rect 842 2968 994 3020
rect 1046 2968 1198 3020
rect 1250 2968 1402 3020
rect 1454 2968 1606 3020
rect 1658 2968 1810 3020
rect 1862 2968 2014 3020
rect 2066 2968 2218 3020
rect 2270 2968 2422 3020
rect 2474 2968 2626 3020
rect 2678 2968 2830 3020
rect 2882 2968 3034 3020
rect 3086 2968 3238 3020
rect 3290 2968 3442 3020
rect 3494 2968 3646 3020
rect 3698 2968 3850 3020
rect 3902 2968 4054 3020
rect 4106 2968 4258 3020
rect 4310 2968 4462 3020
rect 4514 2968 4666 3020
rect 4718 2968 4870 3020
rect 4922 2968 5074 3020
rect 5126 2968 5278 3020
rect 5330 2968 5482 3020
rect 5534 2968 5686 3020
rect 5738 2968 5890 3020
rect 5942 2968 6094 3020
rect 6146 2968 6298 3020
rect 6350 2968 6502 3020
rect 6554 2968 6706 3020
rect 6758 2968 6910 3020
rect 6962 2968 7114 3020
rect 7166 2968 7318 3020
rect 7370 2968 7522 3020
rect 7574 2968 7726 3020
rect 7778 2968 7930 3020
rect 7982 2968 8134 3020
rect 8186 2968 8338 3020
rect 8390 2968 8542 3020
rect 8594 2968 8746 3020
rect 8798 2968 8950 3020
rect 9002 2968 9154 3020
rect 9206 2968 9358 3020
rect 9410 2968 9562 3020
rect 9614 2968 9766 3020
rect 9818 2968 9970 3020
rect 10022 2968 10174 3020
rect 10226 2968 10378 3020
rect 10430 2968 10582 3020
rect 10634 2968 10786 3020
rect 10838 2968 10990 3020
rect 11042 2968 11194 3020
rect 11246 2968 11398 3020
rect 11450 2968 11602 3020
rect 11654 2968 11806 3020
rect 11858 2968 12010 3020
rect 12062 2968 12214 3020
rect 12266 2968 12418 3020
rect 12470 2968 12622 3020
rect 12674 2968 12826 3020
rect 12878 2968 13030 3020
rect 13082 2968 13096 3020
rect 26 2962 13096 2968
rect 1607 2068 1613 2080
rect 0 2040 1613 2068
rect 1607 2028 1613 2040
rect 1665 2068 1671 2080
rect 3239 2068 3245 2080
rect 1665 2040 3245 2068
rect 1665 2028 1671 2040
rect 3239 2028 3245 2040
rect 3297 2068 3303 2080
rect 4871 2068 4877 2080
rect 3297 2040 4877 2068
rect 3297 2028 3303 2040
rect 4871 2028 4877 2040
rect 4929 2068 4935 2080
rect 6503 2068 6509 2080
rect 4929 2040 6509 2068
rect 4929 2028 4935 2040
rect 6503 2028 6509 2040
rect 6561 2068 6567 2080
rect 8135 2068 8141 2080
rect 6561 2040 8141 2068
rect 6561 2028 6567 2040
rect 8135 2028 8141 2040
rect 8193 2068 8199 2080
rect 9767 2068 9773 2080
rect 8193 2040 9773 2068
rect 8193 2028 8199 2040
rect 9767 2028 9773 2040
rect 9825 2068 9831 2080
rect 11399 2068 11405 2080
rect 9825 2040 11405 2068
rect 9825 2028 9831 2040
rect 11399 2028 11405 2040
rect 11457 2068 11463 2080
rect 13031 2068 13037 2080
rect 11457 2040 13037 2068
rect 11457 2028 11463 2040
rect 13031 2028 13037 2040
rect 13089 2028 13095 2080
rect 1403 1864 1409 1876
rect 0 1836 1409 1864
rect 1403 1824 1409 1836
rect 1461 1864 1467 1876
rect 3035 1864 3041 1876
rect 1461 1836 3041 1864
rect 1461 1824 1467 1836
rect 3035 1824 3041 1836
rect 3093 1864 3099 1876
rect 4667 1864 4673 1876
rect 3093 1836 4673 1864
rect 3093 1824 3099 1836
rect 4667 1824 4673 1836
rect 4725 1864 4731 1876
rect 6299 1864 6305 1876
rect 4725 1836 6305 1864
rect 4725 1824 4731 1836
rect 6299 1824 6305 1836
rect 6357 1864 6363 1876
rect 7931 1864 7937 1876
rect 6357 1836 7937 1864
rect 6357 1824 6363 1836
rect 7931 1824 7937 1836
rect 7989 1864 7995 1876
rect 9563 1864 9569 1876
rect 7989 1836 9569 1864
rect 7989 1824 7995 1836
rect 9563 1824 9569 1836
rect 9621 1864 9627 1876
rect 11195 1864 11201 1876
rect 9621 1836 11201 1864
rect 9621 1824 9627 1836
rect 11195 1824 11201 1836
rect 11253 1864 11259 1876
rect 12827 1864 12833 1876
rect 11253 1836 12833 1864
rect 11253 1824 11259 1836
rect 12827 1824 12833 1836
rect 12885 1864 12891 1876
rect 12885 1836 13056 1864
rect 12885 1824 12891 1836
rect 1199 1660 1205 1672
rect 0 1632 1205 1660
rect 1199 1620 1205 1632
rect 1257 1660 1263 1672
rect 2831 1660 2837 1672
rect 1257 1632 2837 1660
rect 1257 1620 1263 1632
rect 2831 1620 2837 1632
rect 2889 1660 2895 1672
rect 4463 1660 4469 1672
rect 2889 1632 4469 1660
rect 2889 1620 2895 1632
rect 4463 1620 4469 1632
rect 4521 1660 4527 1672
rect 6095 1660 6101 1672
rect 4521 1632 6101 1660
rect 4521 1620 4527 1632
rect 6095 1620 6101 1632
rect 6153 1660 6159 1672
rect 7727 1660 7733 1672
rect 6153 1632 7733 1660
rect 6153 1620 6159 1632
rect 7727 1620 7733 1632
rect 7785 1660 7791 1672
rect 9359 1660 9365 1672
rect 7785 1632 9365 1660
rect 7785 1620 7791 1632
rect 9359 1620 9365 1632
rect 9417 1660 9423 1672
rect 10991 1660 10997 1672
rect 9417 1632 10997 1660
rect 9417 1620 9423 1632
rect 10991 1620 10997 1632
rect 11049 1660 11055 1672
rect 12623 1660 12629 1672
rect 11049 1632 12629 1660
rect 11049 1620 11055 1632
rect 12623 1620 12629 1632
rect 12681 1660 12687 1672
rect 12681 1632 13056 1660
rect 12681 1620 12687 1632
rect 995 1456 1001 1468
rect 0 1428 1001 1456
rect 995 1416 1001 1428
rect 1053 1456 1059 1468
rect 2627 1456 2633 1468
rect 1053 1428 2633 1456
rect 1053 1416 1059 1428
rect 2627 1416 2633 1428
rect 2685 1456 2691 1468
rect 4259 1456 4265 1468
rect 2685 1428 4265 1456
rect 2685 1416 2691 1428
rect 4259 1416 4265 1428
rect 4317 1456 4323 1468
rect 5891 1456 5897 1468
rect 4317 1428 5897 1456
rect 4317 1416 4323 1428
rect 5891 1416 5897 1428
rect 5949 1456 5955 1468
rect 7523 1456 7529 1468
rect 5949 1428 7529 1456
rect 5949 1416 5955 1428
rect 7523 1416 7529 1428
rect 7581 1456 7587 1468
rect 9155 1456 9161 1468
rect 7581 1428 9161 1456
rect 7581 1416 7587 1428
rect 9155 1416 9161 1428
rect 9213 1456 9219 1468
rect 10787 1456 10793 1468
rect 9213 1428 10793 1456
rect 9213 1416 9219 1428
rect 10787 1416 10793 1428
rect 10845 1456 10851 1468
rect 12419 1456 12425 1468
rect 10845 1428 12425 1456
rect 10845 1416 10851 1428
rect 12419 1416 12425 1428
rect 12477 1456 12483 1468
rect 12477 1428 13056 1456
rect 12477 1416 12483 1428
rect 791 1252 797 1264
rect 0 1224 797 1252
rect 791 1212 797 1224
rect 849 1252 855 1264
rect 2423 1252 2429 1264
rect 849 1224 2429 1252
rect 849 1212 855 1224
rect 2423 1212 2429 1224
rect 2481 1252 2487 1264
rect 4055 1252 4061 1264
rect 2481 1224 4061 1252
rect 2481 1212 2487 1224
rect 4055 1212 4061 1224
rect 4113 1252 4119 1264
rect 5687 1252 5693 1264
rect 4113 1224 5693 1252
rect 4113 1212 4119 1224
rect 5687 1212 5693 1224
rect 5745 1252 5751 1264
rect 7319 1252 7325 1264
rect 5745 1224 7325 1252
rect 5745 1212 5751 1224
rect 7319 1212 7325 1224
rect 7377 1252 7383 1264
rect 8951 1252 8957 1264
rect 7377 1224 8957 1252
rect 7377 1212 7383 1224
rect 8951 1212 8957 1224
rect 9009 1252 9015 1264
rect 10583 1252 10589 1264
rect 9009 1224 10589 1252
rect 9009 1212 9015 1224
rect 10583 1212 10589 1224
rect 10641 1252 10647 1264
rect 12215 1252 12221 1264
rect 10641 1224 12221 1252
rect 10641 1212 10647 1224
rect 12215 1212 12221 1224
rect 12273 1252 12279 1264
rect 12273 1224 13056 1252
rect 12273 1212 12279 1224
rect 587 1048 593 1060
rect 0 1020 593 1048
rect 587 1008 593 1020
rect 645 1048 651 1060
rect 2219 1048 2225 1060
rect 645 1020 2225 1048
rect 645 1008 651 1020
rect 2219 1008 2225 1020
rect 2277 1048 2283 1060
rect 3851 1048 3857 1060
rect 2277 1020 3857 1048
rect 2277 1008 2283 1020
rect 3851 1008 3857 1020
rect 3909 1048 3915 1060
rect 5483 1048 5489 1060
rect 3909 1020 5489 1048
rect 3909 1008 3915 1020
rect 5483 1008 5489 1020
rect 5541 1048 5547 1060
rect 7115 1048 7121 1060
rect 5541 1020 7121 1048
rect 5541 1008 5547 1020
rect 7115 1008 7121 1020
rect 7173 1048 7179 1060
rect 8747 1048 8753 1060
rect 7173 1020 8753 1048
rect 7173 1008 7179 1020
rect 8747 1008 8753 1020
rect 8805 1048 8811 1060
rect 10379 1048 10385 1060
rect 8805 1020 10385 1048
rect 8805 1008 8811 1020
rect 10379 1008 10385 1020
rect 10437 1048 10443 1060
rect 12011 1048 12017 1060
rect 10437 1020 12017 1048
rect 10437 1008 10443 1020
rect 12011 1008 12017 1020
rect 12069 1048 12075 1060
rect 12069 1020 13056 1048
rect 12069 1008 12075 1020
rect 383 844 389 856
rect 0 816 389 844
rect 383 804 389 816
rect 441 844 447 856
rect 2015 844 2021 856
rect 441 816 2021 844
rect 441 804 447 816
rect 2015 804 2021 816
rect 2073 844 2079 856
rect 3647 844 3653 856
rect 2073 816 3653 844
rect 2073 804 2079 816
rect 3647 804 3653 816
rect 3705 844 3711 856
rect 5279 844 5285 856
rect 3705 816 5285 844
rect 3705 804 3711 816
rect 5279 804 5285 816
rect 5337 844 5343 856
rect 6911 844 6917 856
rect 5337 816 6917 844
rect 5337 804 5343 816
rect 6911 804 6917 816
rect 6969 844 6975 856
rect 8543 844 8549 856
rect 6969 816 8549 844
rect 6969 804 6975 816
rect 8543 804 8549 816
rect 8601 844 8607 856
rect 10175 844 10181 856
rect 8601 816 10181 844
rect 8601 804 8607 816
rect 10175 804 10181 816
rect 10233 844 10239 856
rect 11807 844 11813 856
rect 10233 816 11813 844
rect 10233 804 10239 816
rect 11807 804 11813 816
rect 11865 844 11871 856
rect 11865 816 13056 844
rect 11865 804 11871 816
rect 179 640 185 652
rect 0 612 185 640
rect 179 600 185 612
rect 237 640 243 652
rect 1811 640 1817 652
rect 237 612 1817 640
rect 237 600 243 612
rect 1811 600 1817 612
rect 1869 640 1875 652
rect 3443 640 3449 652
rect 1869 612 3449 640
rect 1869 600 1875 612
rect 3443 600 3449 612
rect 3501 640 3507 652
rect 5075 640 5081 652
rect 3501 612 5081 640
rect 3501 600 3507 612
rect 5075 600 5081 612
rect 5133 640 5139 652
rect 6707 640 6713 652
rect 5133 612 6713 640
rect 5133 600 5139 612
rect 6707 600 6713 612
rect 6765 640 6771 652
rect 8339 640 8345 652
rect 6765 612 8345 640
rect 6765 600 6771 612
rect 8339 600 8345 612
rect 8397 640 8403 652
rect 9971 640 9977 652
rect 8397 612 9977 640
rect 8397 600 8403 612
rect 9971 600 9977 612
rect 10029 640 10035 652
rect 11603 640 11609 652
rect 10029 612 11609 640
rect 10029 600 10035 612
rect 11603 600 11609 612
rect 11661 640 11667 652
rect 11661 612 13056 640
rect 11661 600 11667 612
rect 62 382 68 434
rect 120 422 126 434
rect 266 422 272 434
rect 120 394 272 422
rect 120 382 126 394
rect 266 382 272 394
rect 324 422 330 434
rect 470 422 476 434
rect 324 394 476 422
rect 324 382 330 394
rect 470 382 476 394
rect 528 422 534 434
rect 674 422 680 434
rect 528 394 680 422
rect 528 382 534 394
rect 674 382 680 394
rect 732 422 738 434
rect 878 422 884 434
rect 732 394 884 422
rect 732 382 738 394
rect 878 382 884 394
rect 936 422 942 434
rect 1082 422 1088 434
rect 936 394 1088 422
rect 936 382 942 394
rect 1082 382 1088 394
rect 1140 422 1146 434
rect 1286 422 1292 434
rect 1140 394 1292 422
rect 1140 382 1146 394
rect 1286 382 1292 394
rect 1344 422 1350 434
rect 1490 422 1496 434
rect 1344 394 1496 422
rect 1344 382 1350 394
rect 1490 382 1496 394
rect 1548 382 1554 434
rect 1694 382 1700 434
rect 1752 422 1758 434
rect 1898 422 1904 434
rect 1752 394 1904 422
rect 1752 382 1758 394
rect 1898 382 1904 394
rect 1956 422 1962 434
rect 2102 422 2108 434
rect 1956 394 2108 422
rect 1956 382 1962 394
rect 2102 382 2108 394
rect 2160 422 2166 434
rect 2306 422 2312 434
rect 2160 394 2312 422
rect 2160 382 2166 394
rect 2306 382 2312 394
rect 2364 422 2370 434
rect 2510 422 2516 434
rect 2364 394 2516 422
rect 2364 382 2370 394
rect 2510 382 2516 394
rect 2568 422 2574 434
rect 2714 422 2720 434
rect 2568 394 2720 422
rect 2568 382 2574 394
rect 2714 382 2720 394
rect 2772 422 2778 434
rect 2918 422 2924 434
rect 2772 394 2924 422
rect 2772 382 2778 394
rect 2918 382 2924 394
rect 2976 422 2982 434
rect 3122 422 3128 434
rect 2976 394 3128 422
rect 2976 382 2982 394
rect 3122 382 3128 394
rect 3180 382 3186 434
rect 3326 382 3332 434
rect 3384 422 3390 434
rect 3530 422 3536 434
rect 3384 394 3536 422
rect 3384 382 3390 394
rect 3530 382 3536 394
rect 3588 422 3594 434
rect 3734 422 3740 434
rect 3588 394 3740 422
rect 3588 382 3594 394
rect 3734 382 3740 394
rect 3792 422 3798 434
rect 3938 422 3944 434
rect 3792 394 3944 422
rect 3792 382 3798 394
rect 3938 382 3944 394
rect 3996 422 4002 434
rect 4142 422 4148 434
rect 3996 394 4148 422
rect 3996 382 4002 394
rect 4142 382 4148 394
rect 4200 422 4206 434
rect 4346 422 4352 434
rect 4200 394 4352 422
rect 4200 382 4206 394
rect 4346 382 4352 394
rect 4404 422 4410 434
rect 4550 422 4556 434
rect 4404 394 4556 422
rect 4404 382 4410 394
rect 4550 382 4556 394
rect 4608 422 4614 434
rect 4754 422 4760 434
rect 4608 394 4760 422
rect 4608 382 4614 394
rect 4754 382 4760 394
rect 4812 382 4818 434
rect 4958 382 4964 434
rect 5016 422 5022 434
rect 5162 422 5168 434
rect 5016 394 5168 422
rect 5016 382 5022 394
rect 5162 382 5168 394
rect 5220 422 5226 434
rect 5366 422 5372 434
rect 5220 394 5372 422
rect 5220 382 5226 394
rect 5366 382 5372 394
rect 5424 422 5430 434
rect 5570 422 5576 434
rect 5424 394 5576 422
rect 5424 382 5430 394
rect 5570 382 5576 394
rect 5628 422 5634 434
rect 5774 422 5780 434
rect 5628 394 5780 422
rect 5628 382 5634 394
rect 5774 382 5780 394
rect 5832 422 5838 434
rect 5978 422 5984 434
rect 5832 394 5984 422
rect 5832 382 5838 394
rect 5978 382 5984 394
rect 6036 422 6042 434
rect 6182 422 6188 434
rect 6036 394 6188 422
rect 6036 382 6042 394
rect 6182 382 6188 394
rect 6240 422 6246 434
rect 6386 422 6392 434
rect 6240 394 6392 422
rect 6240 382 6246 394
rect 6386 382 6392 394
rect 6444 382 6450 434
rect 6590 382 6596 434
rect 6648 422 6654 434
rect 6794 422 6800 434
rect 6648 394 6800 422
rect 6648 382 6654 394
rect 6794 382 6800 394
rect 6852 422 6858 434
rect 6998 422 7004 434
rect 6852 394 7004 422
rect 6852 382 6858 394
rect 6998 382 7004 394
rect 7056 422 7062 434
rect 7202 422 7208 434
rect 7056 394 7208 422
rect 7056 382 7062 394
rect 7202 382 7208 394
rect 7260 422 7266 434
rect 7406 422 7412 434
rect 7260 394 7412 422
rect 7260 382 7266 394
rect 7406 382 7412 394
rect 7464 422 7470 434
rect 7610 422 7616 434
rect 7464 394 7616 422
rect 7464 382 7470 394
rect 7610 382 7616 394
rect 7668 422 7674 434
rect 7814 422 7820 434
rect 7668 394 7820 422
rect 7668 382 7674 394
rect 7814 382 7820 394
rect 7872 422 7878 434
rect 8018 422 8024 434
rect 7872 394 8024 422
rect 7872 382 7878 394
rect 8018 382 8024 394
rect 8076 382 8082 434
rect 8222 382 8228 434
rect 8280 422 8286 434
rect 8426 422 8432 434
rect 8280 394 8432 422
rect 8280 382 8286 394
rect 8426 382 8432 394
rect 8484 422 8490 434
rect 8630 422 8636 434
rect 8484 394 8636 422
rect 8484 382 8490 394
rect 8630 382 8636 394
rect 8688 422 8694 434
rect 8834 422 8840 434
rect 8688 394 8840 422
rect 8688 382 8694 394
rect 8834 382 8840 394
rect 8892 422 8898 434
rect 9038 422 9044 434
rect 8892 394 9044 422
rect 8892 382 8898 394
rect 9038 382 9044 394
rect 9096 422 9102 434
rect 9242 422 9248 434
rect 9096 394 9248 422
rect 9096 382 9102 394
rect 9242 382 9248 394
rect 9300 422 9306 434
rect 9446 422 9452 434
rect 9300 394 9452 422
rect 9300 382 9306 394
rect 9446 382 9452 394
rect 9504 422 9510 434
rect 9650 422 9656 434
rect 9504 394 9656 422
rect 9504 382 9510 394
rect 9650 382 9656 394
rect 9708 382 9714 434
rect 9854 382 9860 434
rect 9912 422 9918 434
rect 10058 422 10064 434
rect 9912 394 10064 422
rect 9912 382 9918 394
rect 10058 382 10064 394
rect 10116 422 10122 434
rect 10262 422 10268 434
rect 10116 394 10268 422
rect 10116 382 10122 394
rect 10262 382 10268 394
rect 10320 422 10326 434
rect 10466 422 10472 434
rect 10320 394 10472 422
rect 10320 382 10326 394
rect 10466 382 10472 394
rect 10524 422 10530 434
rect 10670 422 10676 434
rect 10524 394 10676 422
rect 10524 382 10530 394
rect 10670 382 10676 394
rect 10728 422 10734 434
rect 10874 422 10880 434
rect 10728 394 10880 422
rect 10728 382 10734 394
rect 10874 382 10880 394
rect 10932 422 10938 434
rect 11078 422 11084 434
rect 10932 394 11084 422
rect 10932 382 10938 394
rect 11078 382 11084 394
rect 11136 422 11142 434
rect 11282 422 11288 434
rect 11136 394 11288 422
rect 11136 382 11142 394
rect 11282 382 11288 394
rect 11340 382 11346 434
rect 11486 382 11492 434
rect 11544 422 11550 434
rect 11690 422 11696 434
rect 11544 394 11696 422
rect 11544 382 11550 394
rect 11690 382 11696 394
rect 11748 422 11754 434
rect 11894 422 11900 434
rect 11748 394 11900 422
rect 11748 382 11754 394
rect 11894 382 11900 394
rect 11952 422 11958 434
rect 12098 422 12104 434
rect 11952 394 12104 422
rect 11952 382 11958 394
rect 12098 382 12104 394
rect 12156 422 12162 434
rect 12302 422 12308 434
rect 12156 394 12308 422
rect 12156 382 12162 394
rect 12302 382 12308 394
rect 12360 422 12366 434
rect 12506 422 12512 434
rect 12360 394 12512 422
rect 12360 382 12366 394
rect 12506 382 12512 394
rect 12564 422 12570 434
rect 12710 422 12716 434
rect 12564 394 12716 422
rect 12564 382 12570 394
rect 12710 382 12716 394
rect 12768 422 12774 434
rect 12914 422 12920 434
rect 12768 394 12920 422
rect 12768 382 12774 394
rect 12914 382 12920 394
rect 12972 382 12978 434
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_0
timestamp 1581320207
transform 1 0 12852 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_1
timestamp 1581320207
transform 1 0 12648 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_2
timestamp 1581320207
transform 1 0 12444 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_3
timestamp 1581320207
transform 1 0 12240 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_4
timestamp 1581320207
transform 1 0 12036 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_5
timestamp 1581320207
transform 1 0 11832 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_6
timestamp 1581320207
transform 1 0 11628 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_7
timestamp 1581320207
transform 1 0 11424 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_8
timestamp 1581320207
transform 1 0 11220 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_9
timestamp 1581320207
transform 1 0 11016 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_10
timestamp 1581320207
transform 1 0 10812 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_11
timestamp 1581320207
transform 1 0 10608 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_12
timestamp 1581320207
transform 1 0 10404 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_13
timestamp 1581320207
transform 1 0 10200 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_14
timestamp 1581320207
transform 1 0 9996 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_15
timestamp 1581320207
transform 1 0 9792 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_16
timestamp 1581320207
transform 1 0 9588 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_17
timestamp 1581320207
transform 1 0 9384 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_18
timestamp 1581320207
transform 1 0 9180 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_19
timestamp 1581320207
transform 1 0 8976 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_20
timestamp 1581320207
transform 1 0 8772 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_21
timestamp 1581320207
transform 1 0 8568 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_22
timestamp 1581320207
transform 1 0 8364 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_23
timestamp 1581320207
transform 1 0 8160 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_24
timestamp 1581320207
transform 1 0 7956 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_25
timestamp 1581320207
transform 1 0 7752 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_26
timestamp 1581320207
transform 1 0 7548 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_27
timestamp 1581320207
transform 1 0 7344 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_28
timestamp 1581320207
transform 1 0 7140 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_29
timestamp 1581320207
transform 1 0 6936 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_30
timestamp 1581320207
transform 1 0 6732 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_31
timestamp 1581320207
transform 1 0 6528 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_32
timestamp 1581320207
transform 1 0 6324 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_33
timestamp 1581320207
transform 1 0 6120 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_34
timestamp 1581320207
transform 1 0 5916 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_35
timestamp 1581320207
transform 1 0 5712 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_36
timestamp 1581320207
transform 1 0 5508 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_37
timestamp 1581320207
transform 1 0 5304 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_38
timestamp 1581320207
transform 1 0 5100 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_39
timestamp 1581320207
transform 1 0 4896 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_40
timestamp 1581320207
transform 1 0 4692 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_41
timestamp 1581320207
transform 1 0 4488 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_42
timestamp 1581320207
transform 1 0 4284 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_43
timestamp 1581320207
transform 1 0 4080 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_44
timestamp 1581320207
transform 1 0 3876 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_45
timestamp 1581320207
transform 1 0 3672 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_46
timestamp 1581320207
transform 1 0 3468 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_47
timestamp 1581320207
transform 1 0 3264 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_48
timestamp 1581320207
transform 1 0 3060 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_49
timestamp 1581320207
transform 1 0 2856 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_50
timestamp 1581320207
transform 1 0 2652 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_51
timestamp 1581320207
transform 1 0 2448 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_52
timestamp 1581320207
transform 1 0 2244 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_53
timestamp 1581320207
transform 1 0 2040 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_54
timestamp 1581320207
transform 1 0 1836 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_55
timestamp 1581320207
transform 1 0 1632 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_56
timestamp 1581320207
transform 1 0 1428 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_57
timestamp 1581320207
transform 1 0 1224 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_58
timestamp 1581320207
transform 1 0 1020 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_59
timestamp 1581320207
transform 1 0 816 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_60
timestamp 1581320207
transform 1 0 612 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_61
timestamp 1581320207
transform 1 0 408 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_62
timestamp 1581320207
transform 1 0 204 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_63
timestamp 1581320207
transform 1 0 0 0 1 2244
box 1 0 255 817
<< labels >>
rlabel metal2 s 0 612 13056 640 4 sel_0
port 3 nsew
rlabel metal2 s 0 816 13056 844 4 sel_1
port 5 nsew
rlabel metal2 s 0 1020 13056 1048 4 sel_2
port 7 nsew
rlabel metal2 s 0 1224 13056 1252 4 sel_3
port 9 nsew
rlabel metal2 s 0 1428 13056 1456 4 sel_4
port 11 nsew
rlabel metal2 s 0 1632 13056 1660 4 sel_5
port 13 nsew
rlabel metal2 s 0 1836 13056 1864 4 sel_6
port 15 nsew
rlabel metal2 s 0 2040 13056 2068 4 sel_7
port 17 nsew
rlabel metal1 s 80 408 108 2244 4 bl_out_0
port 19 nsew
rlabel metal1 s 1712 408 1740 2244 4 bl_out_1
port 21 nsew
rlabel metal1 s 3344 408 3372 2244 4 bl_out_2
port 23 nsew
rlabel metal1 s 4976 408 5004 2244 4 bl_out_3
port 25 nsew
rlabel metal1 s 6608 408 6636 2244 4 bl_out_4
port 27 nsew
rlabel metal1 s 8240 408 8268 2244 4 bl_out_5
port 29 nsew
rlabel metal1 s 9872 408 9900 2244 4 bl_out_6
port 31 nsew
rlabel metal1 s 11504 408 11532 2244 4 bl_out_7
port 33 nsew
rlabel metal2 s 26 2962 13096 3026 4 gnd
port 35 nsew
rlabel metal1 s 80 2874 108 3026 4 bl_0
port 37 nsew
rlabel metal1 s 284 2874 312 3026 4 bl_1
port 39 nsew
rlabel metal1 s 488 2874 516 3026 4 bl_2
port 41 nsew
rlabel metal1 s 692 2874 720 3026 4 bl_3
port 43 nsew
rlabel metal1 s 896 2874 924 3026 4 bl_4
port 45 nsew
rlabel metal1 s 1100 2874 1128 3026 4 bl_5
port 47 nsew
rlabel metal1 s 1304 2874 1332 3026 4 bl_6
port 49 nsew
rlabel metal1 s 1508 2874 1536 3026 4 bl_7
port 51 nsew
rlabel metal1 s 1712 2874 1740 3026 4 bl_8
port 53 nsew
rlabel metal1 s 1916 2874 1944 3026 4 bl_9
port 55 nsew
rlabel metal1 s 2120 2874 2148 3026 4 bl_10
port 57 nsew
rlabel metal1 s 2324 2874 2352 3026 4 bl_11
port 59 nsew
rlabel metal1 s 2528 2874 2556 3026 4 bl_12
port 61 nsew
rlabel metal1 s 2732 2874 2760 3026 4 bl_13
port 63 nsew
rlabel metal1 s 2936 2874 2964 3026 4 bl_14
port 65 nsew
rlabel metal1 s 3140 2874 3168 3026 4 bl_15
port 67 nsew
rlabel metal1 s 3344 2874 3372 3026 4 bl_16
port 69 nsew
rlabel metal1 s 3548 2874 3576 3026 4 bl_17
port 71 nsew
rlabel metal1 s 3752 2874 3780 3026 4 bl_18
port 73 nsew
rlabel metal1 s 3956 2874 3984 3026 4 bl_19
port 75 nsew
rlabel metal1 s 4160 2874 4188 3026 4 bl_20
port 77 nsew
rlabel metal1 s 4364 2874 4392 3026 4 bl_21
port 79 nsew
rlabel metal1 s 4568 2874 4596 3026 4 bl_22
port 81 nsew
rlabel metal1 s 4772 2874 4800 3026 4 bl_23
port 83 nsew
rlabel metal1 s 4976 2874 5004 3026 4 bl_24
port 85 nsew
rlabel metal1 s 5180 2874 5208 3026 4 bl_25
port 87 nsew
rlabel metal1 s 5384 2874 5412 3026 4 bl_26
port 89 nsew
rlabel metal1 s 5588 2874 5616 3026 4 bl_27
port 91 nsew
rlabel metal1 s 5792 2874 5820 3026 4 bl_28
port 93 nsew
rlabel metal1 s 5996 2874 6024 3026 4 bl_29
port 95 nsew
rlabel metal1 s 6200 2874 6228 3026 4 bl_30
port 97 nsew
rlabel metal1 s 6404 2874 6432 3026 4 bl_31
port 99 nsew
rlabel metal1 s 6608 2874 6636 3026 4 bl_32
port 101 nsew
rlabel metal1 s 6812 2874 6840 3026 4 bl_33
port 103 nsew
rlabel metal1 s 7016 2874 7044 3026 4 bl_34
port 105 nsew
rlabel metal1 s 7220 2874 7248 3026 4 bl_35
port 107 nsew
rlabel metal1 s 7424 2874 7452 3026 4 bl_36
port 109 nsew
rlabel metal1 s 7628 2874 7656 3026 4 bl_37
port 111 nsew
rlabel metal1 s 7832 2874 7860 3026 4 bl_38
port 113 nsew
rlabel metal1 s 8036 2874 8064 3026 4 bl_39
port 115 nsew
rlabel metal1 s 8240 2874 8268 3026 4 bl_40
port 117 nsew
rlabel metal1 s 8444 2874 8472 3026 4 bl_41
port 119 nsew
rlabel metal1 s 8648 2874 8676 3026 4 bl_42
port 121 nsew
rlabel metal1 s 8852 2874 8880 3026 4 bl_43
port 123 nsew
rlabel metal1 s 9056 2874 9084 3026 4 bl_44
port 125 nsew
rlabel metal1 s 9260 2874 9288 3026 4 bl_45
port 127 nsew
rlabel metal1 s 9464 2874 9492 3026 4 bl_46
port 129 nsew
rlabel metal1 s 9668 2874 9696 3026 4 bl_47
port 131 nsew
rlabel metal1 s 9872 2874 9900 3026 4 bl_48
port 133 nsew
rlabel metal1 s 10076 2874 10104 3026 4 bl_49
port 135 nsew
rlabel metal1 s 10280 2874 10308 3026 4 bl_50
port 137 nsew
rlabel metal1 s 10484 2874 10512 3026 4 bl_51
port 139 nsew
rlabel metal1 s 10688 2874 10716 3026 4 bl_52
port 141 nsew
rlabel metal1 s 10892 2874 10920 3026 4 bl_53
port 143 nsew
rlabel metal1 s 11096 2874 11124 3026 4 bl_54
port 145 nsew
rlabel metal1 s 11300 2874 11328 3026 4 bl_55
port 147 nsew
rlabel metal1 s 11504 2874 11532 3026 4 bl_56
port 149 nsew
rlabel metal1 s 11708 2874 11736 3026 4 bl_57
port 151 nsew
rlabel metal1 s 11912 2874 11940 3026 4 bl_58
port 153 nsew
rlabel metal1 s 12116 2874 12144 3026 4 bl_59
port 155 nsew
rlabel metal1 s 12320 2874 12348 3026 4 bl_60
port 157 nsew
rlabel metal1 s 12524 2874 12552 3026 4 bl_61
port 159 nsew
rlabel metal1 s 12728 2874 12756 3026 4 bl_62
port 161 nsew
rlabel metal1 s 12932 2874 12960 3026 4 bl_63
port 163 nsew
<< properties >>
string FIXED_BBOX 0 0 13056 2001
<< end >>
