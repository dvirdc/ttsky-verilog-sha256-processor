magic
tech sky130A
magscale 1 2
timestamp 1581321280
<< checkpaint >>
rect -2756 -2756 19622 20168
<< locali >>
rect 6679 17038 6713 17054
rect 6679 16988 6713 17004
rect 6679 16834 6713 16850
rect 6679 16784 6713 16800
rect 6679 16526 6713 16542
rect 6679 16476 6713 16492
rect 6679 16322 6713 16338
rect 6679 16272 6713 16288
rect 6679 16118 6713 16134
rect 6679 16068 6713 16084
rect 6679 15914 6713 15930
rect 6679 15864 6713 15880
rect 6679 15710 6713 15726
rect 6679 15660 6713 15676
rect 6679 15506 6713 15522
rect 6679 15456 6713 15472
rect 6679 15302 6713 15318
rect 6679 15252 6713 15268
rect 6679 15098 6713 15114
rect 6679 15048 6713 15064
rect 6679 14790 6713 14806
rect 6679 14740 6713 14756
rect 6679 14586 6713 14602
rect 6679 14536 6713 14552
rect 6679 14382 6713 14398
rect 6679 14332 6713 14348
rect 6679 14178 6713 14194
rect 6679 14128 6713 14144
rect 6679 13974 6713 13990
rect 6679 13924 6713 13940
rect 6679 13770 6713 13786
rect 6679 13720 6713 13736
rect 6679 13566 6713 13582
rect 6679 13516 6713 13532
rect 6679 13362 6713 13378
rect 6679 13312 6713 13328
rect 6679 13054 6713 13070
rect 6679 13004 6713 13020
rect 6679 12850 6713 12866
rect 6679 12800 6713 12816
rect 6679 12646 6713 12662
rect 6679 12596 6713 12612
rect 6679 12442 6713 12458
rect 6679 12392 6713 12408
rect 6679 12238 6713 12254
rect 6679 12188 6713 12204
rect 6679 12034 6713 12050
rect 6679 11984 6713 12000
rect 6679 11830 6713 11846
rect 6679 11780 6713 11796
rect 6679 11626 6713 11642
rect 6679 11576 6713 11592
rect 6679 11318 6713 11334
rect 6679 11268 6713 11284
rect 6679 11114 6713 11130
rect 6679 11064 6713 11080
rect 6679 10910 6713 10926
rect 6679 10860 6713 10876
rect 6679 10706 6713 10722
rect 6679 10656 6713 10672
rect 6679 10502 6713 10518
rect 6679 10452 6713 10468
rect 6679 10298 6713 10314
rect 6679 10248 6713 10264
rect 6679 10094 6713 10110
rect 6679 10044 6713 10060
rect 6679 9890 6713 9906
rect 6679 9840 6713 9856
rect 6679 9582 6713 9598
rect 6679 9532 6713 9548
rect 6679 9378 6713 9394
rect 6679 9328 6713 9344
rect 6679 9174 6713 9190
rect 6679 9124 6713 9140
rect 6679 8970 6713 8986
rect 6679 8920 6713 8936
rect 6679 8766 6713 8782
rect 6679 8716 6713 8732
rect 6679 8562 6713 8578
rect 6679 8512 6713 8528
rect 6679 8358 6713 8374
rect 6679 8308 6713 8324
rect 6679 8154 6713 8170
rect 6679 8104 6713 8120
rect 6934 7029 6950 7063
rect 6984 7029 7000 7063
rect 7138 7029 7154 7063
rect 7188 7029 7204 7063
rect 7342 7029 7358 7063
rect 7392 7029 7408 7063
rect 7546 7029 7562 7063
rect 7596 7029 7612 7063
rect 7750 7029 7766 7063
rect 7800 7029 7816 7063
rect 7954 7029 7970 7063
rect 8004 7029 8020 7063
rect 8158 7029 8174 7063
rect 8208 7029 8224 7063
rect 8362 7029 8378 7063
rect 8412 7029 8428 7063
rect 8566 7029 8582 7063
rect 8616 7029 8632 7063
rect 8770 7029 8786 7063
rect 8820 7029 8836 7063
rect 8974 7029 8990 7063
rect 9024 7029 9040 7063
rect 9178 7029 9194 7063
rect 9228 7029 9244 7063
rect 9382 7029 9398 7063
rect 9432 7029 9448 7063
rect 9586 7029 9602 7063
rect 9636 7029 9652 7063
rect 9790 7029 9806 7063
rect 9840 7029 9856 7063
rect 9994 7029 10010 7063
rect 10044 7029 10060 7063
rect 10198 7029 10214 7063
rect 10248 7029 10264 7063
rect 10402 7029 10418 7063
rect 10452 7029 10468 7063
rect 10606 7029 10622 7063
rect 10656 7029 10672 7063
rect 10810 7029 10826 7063
rect 10860 7029 10876 7063
rect 11014 7029 11030 7063
rect 11064 7029 11080 7063
rect 11218 7029 11234 7063
rect 11268 7029 11284 7063
rect 11422 7029 11438 7063
rect 11472 7029 11488 7063
rect 11626 7029 11642 7063
rect 11676 7029 11692 7063
rect 11830 7029 11846 7063
rect 11880 7029 11896 7063
rect 12034 7029 12050 7063
rect 12084 7029 12100 7063
rect 12238 7029 12254 7063
rect 12288 7029 12304 7063
rect 12442 7029 12458 7063
rect 12492 7029 12508 7063
rect 12646 7029 12662 7063
rect 12696 7029 12712 7063
rect 12850 7029 12866 7063
rect 12900 7029 12916 7063
rect 13054 7029 13070 7063
rect 13104 7029 13120 7063
rect 13258 7029 13274 7063
rect 13308 7029 13324 7063
rect 13462 7029 13478 7063
rect 13512 7029 13528 7063
rect 13666 7029 13682 7063
rect 13716 7029 13732 7063
rect 13870 7029 13886 7063
rect 13920 7029 13936 7063
rect 14074 7029 14090 7063
rect 14124 7029 14140 7063
rect 14278 7029 14294 7063
rect 14328 7029 14344 7063
rect 14482 7029 14498 7063
rect 14532 7029 14548 7063
rect 14686 7029 14702 7063
rect 14736 7029 14752 7063
rect 14890 7029 14906 7063
rect 14940 7029 14956 7063
rect 15094 7029 15110 7063
rect 15144 7029 15160 7063
rect 15298 7029 15314 7063
rect 15348 7029 15364 7063
rect 15502 7029 15518 7063
rect 15552 7029 15568 7063
rect 15706 7029 15722 7063
rect 15756 7029 15772 7063
rect 15910 7029 15926 7063
rect 15960 7029 15976 7063
rect 16114 7029 16130 7063
rect 16164 7029 16180 7063
rect 16318 7029 16334 7063
rect 16368 7029 16384 7063
rect 16522 7029 16538 7063
rect 16572 7029 16588 7063
rect 6934 5434 6950 5468
rect 6984 5434 7000 5468
rect 7138 5434 7154 5468
rect 7188 5434 7204 5468
rect 7342 5434 7358 5468
rect 7392 5434 7408 5468
rect 7546 5434 7562 5468
rect 7596 5434 7612 5468
rect 7750 5434 7766 5468
rect 7800 5434 7816 5468
rect 7954 5434 7970 5468
rect 8004 5434 8020 5468
rect 8158 5434 8174 5468
rect 8208 5434 8224 5468
rect 8362 5434 8378 5468
rect 8412 5434 8428 5468
rect 8566 5434 8582 5468
rect 8616 5434 8632 5468
rect 8770 5434 8786 5468
rect 8820 5434 8836 5468
rect 8974 5434 8990 5468
rect 9024 5434 9040 5468
rect 9178 5434 9194 5468
rect 9228 5434 9244 5468
rect 9382 5434 9398 5468
rect 9432 5434 9448 5468
rect 9586 5434 9602 5468
rect 9636 5434 9652 5468
rect 9790 5434 9806 5468
rect 9840 5434 9856 5468
rect 9994 5434 10010 5468
rect 10044 5434 10060 5468
rect 10198 5434 10214 5468
rect 10248 5434 10264 5468
rect 10402 5434 10418 5468
rect 10452 5434 10468 5468
rect 10606 5434 10622 5468
rect 10656 5434 10672 5468
rect 10810 5434 10826 5468
rect 10860 5434 10876 5468
rect 11014 5434 11030 5468
rect 11064 5434 11080 5468
rect 11218 5434 11234 5468
rect 11268 5434 11284 5468
rect 11422 5434 11438 5468
rect 11472 5434 11488 5468
rect 11626 5434 11642 5468
rect 11676 5434 11692 5468
rect 11830 5434 11846 5468
rect 11880 5434 11896 5468
rect 12034 5434 12050 5468
rect 12084 5434 12100 5468
rect 12238 5434 12254 5468
rect 12288 5434 12304 5468
rect 12442 5434 12458 5468
rect 12492 5434 12508 5468
rect 12646 5434 12662 5468
rect 12696 5434 12712 5468
rect 12850 5434 12866 5468
rect 12900 5434 12916 5468
rect 13054 5434 13070 5468
rect 13104 5434 13120 5468
rect 13258 5434 13274 5468
rect 13308 5434 13324 5468
rect 13462 5434 13478 5468
rect 13512 5434 13528 5468
rect 13666 5434 13682 5468
rect 13716 5434 13732 5468
rect 13870 5434 13886 5468
rect 13920 5434 13936 5468
rect 14074 5434 14090 5468
rect 14124 5434 14140 5468
rect 14278 5434 14294 5468
rect 14328 5434 14344 5468
rect 14482 5434 14498 5468
rect 14532 5434 14548 5468
rect 14686 5434 14702 5468
rect 14736 5434 14752 5468
rect 14890 5434 14906 5468
rect 14940 5434 14956 5468
rect 15094 5434 15110 5468
rect 15144 5434 15160 5468
rect 15298 5434 15314 5468
rect 15348 5434 15364 5468
rect 15502 5434 15518 5468
rect 15552 5434 15568 5468
rect 15706 5434 15722 5468
rect 15756 5434 15772 5468
rect 15910 5434 15926 5468
rect 15960 5434 15976 5468
rect 16114 5434 16130 5468
rect 16164 5434 16180 5468
rect 16318 5434 16334 5468
rect 16368 5434 16384 5468
rect 16522 5434 16538 5468
rect 16572 5434 16588 5468
rect 337 4793 371 4809
rect 337 4743 371 4759
rect 745 4793 779 4809
rect 745 4743 779 4759
rect 1153 4793 1187 4809
rect 1153 4743 1187 4759
rect 1561 4793 1595 4809
rect 1561 4743 1595 4759
rect 1969 4793 2003 4809
rect 1969 4743 2003 4759
rect 2377 4793 2411 4809
rect 2377 4743 2411 4759
rect 6679 4113 6713 4129
rect 6679 4063 6713 4079
rect 6679 3909 6713 3925
rect 6679 3859 6713 3875
rect 6679 3705 6713 3721
rect 6679 3655 6713 3671
rect 2865 3628 2899 3644
rect 2865 3578 2899 3594
rect 10148 1739 10182 1755
rect 10148 1689 10182 1705
rect 10456 1739 10490 1755
rect 10456 1689 10490 1705
rect 10764 1739 10798 1755
rect 10764 1689 10798 1705
rect 11072 1739 11106 1755
rect 11072 1689 11106 1705
rect 11380 1739 11414 1755
rect 11380 1689 11414 1705
rect 11688 1739 11722 1755
rect 11688 1689 11722 1705
rect 11996 1739 12030 1755
rect 11996 1689 12030 1705
rect 12304 1739 12338 1755
rect 12304 1689 12338 1705
rect 12612 1739 12646 1755
rect 12612 1689 12646 1705
rect 12920 1739 12954 1755
rect 12920 1689 12954 1705
rect 13228 1739 13262 1755
rect 13228 1689 13262 1705
rect 13536 1739 13570 1755
rect 13536 1689 13570 1705
rect 13844 1739 13878 1755
rect 13844 1689 13878 1705
rect 14152 1739 14186 1755
rect 14152 1689 14186 1705
rect 14460 1739 14494 1755
rect 14460 1689 14494 1705
rect 14768 1739 14802 1755
rect 14768 1689 14802 1705
rect 520 1421 554 1437
rect 520 1371 554 1387
rect 2497 1409 2531 1425
rect 2497 1359 2531 1375
rect 3120 670 3154 686
rect 3120 620 3154 636
rect 3963 344 3997 360
rect 3963 294 3997 310
rect 4371 344 4405 360
rect 4371 294 4405 310
rect 10132 0 10148 34
rect 10182 0 10198 34
rect 10440 0 10456 34
rect 10490 0 10506 34
rect 10748 0 10764 34
rect 10798 0 10814 34
rect 11056 0 11072 34
rect 11106 0 11122 34
rect 11364 0 11380 34
rect 11414 0 11430 34
rect 11672 0 11688 34
rect 11722 0 11738 34
rect 11980 0 11996 34
rect 12030 0 12046 34
rect 12288 0 12304 34
rect 12338 0 12354 34
rect 12596 0 12612 34
rect 12646 0 12662 34
rect 12904 0 12920 34
rect 12954 0 12970 34
rect 13212 0 13228 34
rect 13262 0 13278 34
rect 13520 0 13536 34
rect 13570 0 13586 34
rect 13828 0 13844 34
rect 13878 0 13894 34
rect 14136 0 14152 34
rect 14186 0 14202 34
rect 14444 0 14460 34
rect 14494 0 14510 34
rect 14752 0 14768 34
rect 14802 0 14818 34
<< viali >>
rect 6679 17004 6713 17038
rect 6679 16800 6713 16834
rect 6679 16492 6713 16526
rect 6679 16288 6713 16322
rect 6679 16084 6713 16118
rect 6679 15880 6713 15914
rect 6679 15676 6713 15710
rect 6679 15472 6713 15506
rect 6679 15268 6713 15302
rect 6679 15064 6713 15098
rect 6679 14756 6713 14790
rect 6679 14552 6713 14586
rect 6679 14348 6713 14382
rect 6679 14144 6713 14178
rect 6679 13940 6713 13974
rect 6679 13736 6713 13770
rect 6679 13532 6713 13566
rect 6679 13328 6713 13362
rect 6679 13020 6713 13054
rect 6679 12816 6713 12850
rect 6679 12612 6713 12646
rect 6679 12408 6713 12442
rect 6679 12204 6713 12238
rect 6679 12000 6713 12034
rect 6679 11796 6713 11830
rect 6679 11592 6713 11626
rect 6679 11284 6713 11318
rect 6679 11080 6713 11114
rect 6679 10876 6713 10910
rect 6679 10672 6713 10706
rect 6679 10468 6713 10502
rect 6679 10264 6713 10298
rect 6679 10060 6713 10094
rect 6679 9856 6713 9890
rect 6679 9548 6713 9582
rect 6679 9344 6713 9378
rect 6679 9140 6713 9174
rect 6679 8936 6713 8970
rect 6679 8732 6713 8766
rect 6679 8528 6713 8562
rect 6679 8324 6713 8358
rect 6679 8120 6713 8154
rect 6950 7029 6984 7063
rect 7154 7029 7188 7063
rect 7358 7029 7392 7063
rect 7562 7029 7596 7063
rect 7766 7029 7800 7063
rect 7970 7029 8004 7063
rect 8174 7029 8208 7063
rect 8378 7029 8412 7063
rect 8582 7029 8616 7063
rect 8786 7029 8820 7063
rect 8990 7029 9024 7063
rect 9194 7029 9228 7063
rect 9398 7029 9432 7063
rect 9602 7029 9636 7063
rect 9806 7029 9840 7063
rect 10010 7029 10044 7063
rect 10214 7029 10248 7063
rect 10418 7029 10452 7063
rect 10622 7029 10656 7063
rect 10826 7029 10860 7063
rect 11030 7029 11064 7063
rect 11234 7029 11268 7063
rect 11438 7029 11472 7063
rect 11642 7029 11676 7063
rect 11846 7029 11880 7063
rect 12050 7029 12084 7063
rect 12254 7029 12288 7063
rect 12458 7029 12492 7063
rect 12662 7029 12696 7063
rect 12866 7029 12900 7063
rect 13070 7029 13104 7063
rect 13274 7029 13308 7063
rect 13478 7029 13512 7063
rect 13682 7029 13716 7063
rect 13886 7029 13920 7063
rect 14090 7029 14124 7063
rect 14294 7029 14328 7063
rect 14498 7029 14532 7063
rect 14702 7029 14736 7063
rect 14906 7029 14940 7063
rect 15110 7029 15144 7063
rect 15314 7029 15348 7063
rect 15518 7029 15552 7063
rect 15722 7029 15756 7063
rect 15926 7029 15960 7063
rect 16130 7029 16164 7063
rect 16334 7029 16368 7063
rect 16538 7029 16572 7063
rect 6950 5434 6984 5468
rect 7154 5434 7188 5468
rect 7358 5434 7392 5468
rect 7562 5434 7596 5468
rect 7766 5434 7800 5468
rect 7970 5434 8004 5468
rect 8174 5434 8208 5468
rect 8378 5434 8412 5468
rect 8582 5434 8616 5468
rect 8786 5434 8820 5468
rect 8990 5434 9024 5468
rect 9194 5434 9228 5468
rect 9398 5434 9432 5468
rect 9602 5434 9636 5468
rect 9806 5434 9840 5468
rect 10010 5434 10044 5468
rect 10214 5434 10248 5468
rect 10418 5434 10452 5468
rect 10622 5434 10656 5468
rect 10826 5434 10860 5468
rect 11030 5434 11064 5468
rect 11234 5434 11268 5468
rect 11438 5434 11472 5468
rect 11642 5434 11676 5468
rect 11846 5434 11880 5468
rect 12050 5434 12084 5468
rect 12254 5434 12288 5468
rect 12458 5434 12492 5468
rect 12662 5434 12696 5468
rect 12866 5434 12900 5468
rect 13070 5434 13104 5468
rect 13274 5434 13308 5468
rect 13478 5434 13512 5468
rect 13682 5434 13716 5468
rect 13886 5434 13920 5468
rect 14090 5434 14124 5468
rect 14294 5434 14328 5468
rect 14498 5434 14532 5468
rect 14702 5434 14736 5468
rect 14906 5434 14940 5468
rect 15110 5434 15144 5468
rect 15314 5434 15348 5468
rect 15518 5434 15552 5468
rect 15722 5434 15756 5468
rect 15926 5434 15960 5468
rect 16130 5434 16164 5468
rect 16334 5434 16368 5468
rect 16538 5434 16572 5468
rect 337 4759 371 4793
rect 745 4759 779 4793
rect 1153 4759 1187 4793
rect 1561 4759 1595 4793
rect 1969 4759 2003 4793
rect 2377 4759 2411 4793
rect 6679 4079 6713 4113
rect 6679 3875 6713 3909
rect 6679 3671 6713 3705
rect 2865 3594 2899 3628
rect 10148 1705 10182 1739
rect 10456 1705 10490 1739
rect 10764 1705 10798 1739
rect 11072 1705 11106 1739
rect 11380 1705 11414 1739
rect 11688 1705 11722 1739
rect 11996 1705 12030 1739
rect 12304 1705 12338 1739
rect 12612 1705 12646 1739
rect 12920 1705 12954 1739
rect 13228 1705 13262 1739
rect 13536 1705 13570 1739
rect 13844 1705 13878 1739
rect 14152 1705 14186 1739
rect 14460 1705 14494 1739
rect 14768 1705 14802 1739
rect 520 1387 554 1421
rect 2497 1375 2531 1409
rect 3120 636 3154 670
rect 3963 310 3997 344
rect 4371 310 4405 344
rect 10148 0 10182 34
rect 10456 0 10490 34
rect 10764 0 10798 34
rect 11072 0 11106 34
rect 11380 0 11414 34
rect 11688 0 11722 34
rect 11996 0 12030 34
rect 12304 0 12338 34
rect 12612 0 12646 34
rect 12920 0 12954 34
rect 13228 0 13262 34
rect 13536 0 13570 34
rect 13844 0 13878 34
rect 14152 0 14186 34
rect 14460 0 14494 34
rect 14768 0 14802 34
<< metal1 >>
rect 6921 17326 6927 17378
rect 6979 17326 6985 17378
rect 16537 17326 16543 17378
rect 16595 17326 16601 17378
rect 3691 17115 3697 17167
rect 3749 17115 3755 17167
rect 4087 17115 4093 17167
rect 4145 17115 4151 17167
rect 4697 17115 4703 17167
rect 4755 17115 4761 17167
rect 5945 17115 5951 17167
rect 6003 17115 6009 17167
rect 6667 17038 6725 17044
rect 6667 17004 6679 17038
rect 6713 17035 6725 17038
rect 6826 17035 6832 17047
rect 6713 17007 6832 17035
rect 6713 17004 6725 17007
rect 6667 16998 6725 17004
rect 6826 16995 6832 17007
rect 6884 16995 6890 17047
rect 6667 16834 6725 16840
rect 6667 16800 6679 16834
rect 6713 16831 6725 16834
rect 6826 16831 6832 16843
rect 6713 16803 6832 16831
rect 6713 16800 6725 16803
rect 6667 16794 6725 16800
rect 6826 16791 6832 16803
rect 6884 16791 6890 16843
rect 6667 16526 6725 16532
rect 6667 16492 6679 16526
rect 6713 16523 6725 16526
rect 6826 16523 6832 16535
rect 6713 16495 6832 16523
rect 6713 16492 6725 16495
rect 6667 16486 6725 16492
rect 6826 16483 6832 16495
rect 6884 16483 6890 16535
rect 6667 16322 6725 16328
rect 6667 16288 6679 16322
rect 6713 16319 6725 16322
rect 6826 16319 6832 16331
rect 6713 16291 6832 16319
rect 6713 16288 6725 16291
rect 6667 16282 6725 16288
rect 6826 16279 6832 16291
rect 6884 16279 6890 16331
rect 6667 16118 6725 16124
rect 6667 16084 6679 16118
rect 6713 16115 6725 16118
rect 6826 16115 6832 16127
rect 6713 16087 6832 16115
rect 6713 16084 6725 16087
rect 6667 16078 6725 16084
rect 6826 16075 6832 16087
rect 6884 16075 6890 16127
rect 6667 15914 6725 15920
rect 6667 15880 6679 15914
rect 6713 15911 6725 15914
rect 6826 15911 6832 15923
rect 6713 15883 6832 15911
rect 6713 15880 6725 15883
rect 6667 15874 6725 15880
rect 6826 15871 6832 15883
rect 6884 15871 6890 15923
rect 6667 15710 6725 15716
rect 6667 15676 6679 15710
rect 6713 15707 6725 15710
rect 6826 15707 6832 15719
rect 6713 15679 6832 15707
rect 6713 15676 6725 15679
rect 6667 15670 6725 15676
rect 6826 15667 6832 15679
rect 6884 15667 6890 15719
rect 6667 15506 6725 15512
rect 6667 15472 6679 15506
rect 6713 15503 6725 15506
rect 6826 15503 6832 15515
rect 6713 15475 6832 15503
rect 6713 15472 6725 15475
rect 6667 15466 6725 15472
rect 6826 15463 6832 15475
rect 6884 15463 6890 15515
rect 6667 15302 6725 15308
rect 6667 15268 6679 15302
rect 6713 15299 6725 15302
rect 6826 15299 6832 15311
rect 6713 15271 6832 15299
rect 6713 15268 6725 15271
rect 6667 15262 6725 15268
rect 6826 15259 6832 15271
rect 6884 15259 6890 15311
rect 6667 15098 6725 15104
rect 6667 15064 6679 15098
rect 6713 15095 6725 15098
rect 6826 15095 6832 15107
rect 6713 15067 6832 15095
rect 6713 15064 6725 15067
rect 6667 15058 6725 15064
rect 6826 15055 6832 15067
rect 6884 15055 6890 15107
rect 6667 14790 6725 14796
rect 6667 14756 6679 14790
rect 6713 14787 6725 14790
rect 6826 14787 6832 14799
rect 6713 14759 6832 14787
rect 6713 14756 6725 14759
rect 6667 14750 6725 14756
rect 6826 14747 6832 14759
rect 6884 14747 6890 14799
rect 6667 14586 6725 14592
rect 6667 14552 6679 14586
rect 6713 14583 6725 14586
rect 6826 14583 6832 14595
rect 6713 14555 6832 14583
rect 6713 14552 6725 14555
rect 6667 14546 6725 14552
rect 6826 14543 6832 14555
rect 6884 14543 6890 14595
rect 6667 14382 6725 14388
rect 6667 14348 6679 14382
rect 6713 14379 6725 14382
rect 6826 14379 6832 14391
rect 6713 14351 6832 14379
rect 6713 14348 6725 14351
rect 6667 14342 6725 14348
rect 6826 14339 6832 14351
rect 6884 14339 6890 14391
rect 6667 14178 6725 14184
rect 6667 14144 6679 14178
rect 6713 14175 6725 14178
rect 6826 14175 6832 14187
rect 6713 14147 6832 14175
rect 6713 14144 6725 14147
rect 6667 14138 6725 14144
rect 6826 14135 6832 14147
rect 6884 14135 6890 14187
rect 6667 13974 6725 13980
rect 6667 13940 6679 13974
rect 6713 13971 6725 13974
rect 6826 13971 6832 13983
rect 6713 13943 6832 13971
rect 6713 13940 6725 13943
rect 6667 13934 6725 13940
rect 6826 13931 6832 13943
rect 6884 13931 6890 13983
rect 6667 13770 6725 13776
rect 6667 13736 6679 13770
rect 6713 13767 6725 13770
rect 6826 13767 6832 13779
rect 6713 13739 6832 13767
rect 6713 13736 6725 13739
rect 6667 13730 6725 13736
rect 6826 13727 6832 13739
rect 6884 13727 6890 13779
rect 6667 13566 6725 13572
rect 6667 13532 6679 13566
rect 6713 13563 6725 13566
rect 6826 13563 6832 13575
rect 6713 13535 6832 13563
rect 6713 13532 6725 13535
rect 6667 13526 6725 13532
rect 6826 13523 6832 13535
rect 6884 13523 6890 13575
rect 6667 13362 6725 13368
rect 6667 13328 6679 13362
rect 6713 13359 6725 13362
rect 6826 13359 6832 13371
rect 6713 13331 6832 13359
rect 6713 13328 6725 13331
rect 6667 13322 6725 13328
rect 6826 13319 6832 13331
rect 6884 13319 6890 13371
rect 6667 13054 6725 13060
rect 6667 13020 6679 13054
rect 6713 13051 6725 13054
rect 6826 13051 6832 13063
rect 6713 13023 6832 13051
rect 6713 13020 6725 13023
rect 6667 13014 6725 13020
rect 6826 13011 6832 13023
rect 6884 13011 6890 13063
rect 6667 12850 6725 12856
rect 6667 12816 6679 12850
rect 6713 12847 6725 12850
rect 6826 12847 6832 12859
rect 6713 12819 6832 12847
rect 6713 12816 6725 12819
rect 6667 12810 6725 12816
rect 6826 12807 6832 12819
rect 6884 12807 6890 12859
rect 6667 12646 6725 12652
rect 6667 12612 6679 12646
rect 6713 12643 6725 12646
rect 6826 12643 6832 12655
rect 6713 12615 6832 12643
rect 6713 12612 6725 12615
rect 6667 12606 6725 12612
rect 6826 12603 6832 12615
rect 6884 12603 6890 12655
rect 6667 12442 6725 12448
rect 6667 12408 6679 12442
rect 6713 12439 6725 12442
rect 6826 12439 6832 12451
rect 6713 12411 6832 12439
rect 6713 12408 6725 12411
rect 6667 12402 6725 12408
rect 6826 12399 6832 12411
rect 6884 12399 6890 12451
rect 6667 12238 6725 12244
rect 6667 12204 6679 12238
rect 6713 12235 6725 12238
rect 6826 12235 6832 12247
rect 6713 12207 6832 12235
rect 6713 12204 6725 12207
rect 6667 12198 6725 12204
rect 6826 12195 6832 12207
rect 6884 12195 6890 12247
rect 6667 12034 6725 12040
rect 6667 12000 6679 12034
rect 6713 12031 6725 12034
rect 6826 12031 6832 12043
rect 6713 12003 6832 12031
rect 6713 12000 6725 12003
rect 6667 11994 6725 12000
rect 6826 11991 6832 12003
rect 6884 11991 6890 12043
rect 6667 11830 6725 11836
rect 6667 11796 6679 11830
rect 6713 11827 6725 11830
rect 6826 11827 6832 11839
rect 6713 11799 6832 11827
rect 6713 11796 6725 11799
rect 6667 11790 6725 11796
rect 6826 11787 6832 11799
rect 6884 11787 6890 11839
rect 6667 11626 6725 11632
rect 6667 11592 6679 11626
rect 6713 11623 6725 11626
rect 6826 11623 6832 11635
rect 6713 11595 6832 11623
rect 6713 11592 6725 11595
rect 6667 11586 6725 11592
rect 6826 11583 6832 11595
rect 6884 11583 6890 11635
rect 6667 11318 6725 11324
rect 6667 11284 6679 11318
rect 6713 11315 6725 11318
rect 6826 11315 6832 11327
rect 6713 11287 6832 11315
rect 6713 11284 6725 11287
rect 6667 11278 6725 11284
rect 6826 11275 6832 11287
rect 6884 11275 6890 11327
rect 6667 11114 6725 11120
rect 6667 11080 6679 11114
rect 6713 11111 6725 11114
rect 6826 11111 6832 11123
rect 6713 11083 6832 11111
rect 6713 11080 6725 11083
rect 6667 11074 6725 11080
rect 6826 11071 6832 11083
rect 6884 11071 6890 11123
rect 6667 10910 6725 10916
rect 6667 10876 6679 10910
rect 6713 10907 6725 10910
rect 6826 10907 6832 10919
rect 6713 10879 6832 10907
rect 6713 10876 6725 10879
rect 6667 10870 6725 10876
rect 6826 10867 6832 10879
rect 6884 10867 6890 10919
rect 6667 10706 6725 10712
rect 6667 10672 6679 10706
rect 6713 10703 6725 10706
rect 6826 10703 6832 10715
rect 6713 10675 6832 10703
rect 6713 10672 6725 10675
rect 6667 10666 6725 10672
rect 6826 10663 6832 10675
rect 6884 10663 6890 10715
rect 6667 10502 6725 10508
rect 6667 10468 6679 10502
rect 6713 10499 6725 10502
rect 6826 10499 6832 10511
rect 6713 10471 6832 10499
rect 6713 10468 6725 10471
rect 6667 10462 6725 10468
rect 6826 10459 6832 10471
rect 6884 10459 6890 10511
rect 6667 10298 6725 10304
rect 6667 10264 6679 10298
rect 6713 10295 6725 10298
rect 6826 10295 6832 10307
rect 6713 10267 6832 10295
rect 6713 10264 6725 10267
rect 6667 10258 6725 10264
rect 6826 10255 6832 10267
rect 6884 10255 6890 10307
rect 6667 10094 6725 10100
rect 6667 10060 6679 10094
rect 6713 10091 6725 10094
rect 6826 10091 6832 10103
rect 6713 10063 6832 10091
rect 6713 10060 6725 10063
rect 6667 10054 6725 10060
rect 6826 10051 6832 10063
rect 6884 10051 6890 10103
rect 6667 9890 6725 9896
rect 6667 9856 6679 9890
rect 6713 9887 6725 9890
rect 6826 9887 6832 9899
rect 6713 9859 6832 9887
rect 6713 9856 6725 9859
rect 6667 9850 6725 9856
rect 6826 9847 6832 9859
rect 6884 9847 6890 9899
rect 6667 9582 6725 9588
rect 6667 9548 6679 9582
rect 6713 9579 6725 9582
rect 6826 9579 6832 9591
rect 6713 9551 6832 9579
rect 6713 9548 6725 9551
rect 6667 9542 6725 9548
rect 6826 9539 6832 9551
rect 6884 9539 6890 9591
rect 6667 9378 6725 9384
rect 6667 9344 6679 9378
rect 6713 9375 6725 9378
rect 6826 9375 6832 9387
rect 6713 9347 6832 9375
rect 6713 9344 6725 9347
rect 6667 9338 6725 9344
rect 6826 9335 6832 9347
rect 6884 9335 6890 9387
rect 6667 9174 6725 9180
rect 6667 9140 6679 9174
rect 6713 9171 6725 9174
rect 6826 9171 6832 9183
rect 6713 9143 6832 9171
rect 6713 9140 6725 9143
rect 6667 9134 6725 9140
rect 6826 9131 6832 9143
rect 6884 9131 6890 9183
rect 6667 8970 6725 8976
rect 6667 8936 6679 8970
rect 6713 8967 6725 8970
rect 6826 8967 6832 8979
rect 6713 8939 6832 8967
rect 6713 8936 6725 8939
rect 6667 8930 6725 8936
rect 6826 8927 6832 8939
rect 6884 8927 6890 8979
rect 6667 8766 6725 8772
rect 6667 8732 6679 8766
rect 6713 8763 6725 8766
rect 6826 8763 6832 8775
rect 6713 8735 6832 8763
rect 6713 8732 6725 8735
rect 6667 8726 6725 8732
rect 6826 8723 6832 8735
rect 6884 8723 6890 8775
rect 6667 8562 6725 8568
rect 6667 8528 6679 8562
rect 6713 8559 6725 8562
rect 6826 8559 6832 8571
rect 6713 8531 6832 8559
rect 6713 8528 6725 8531
rect 6667 8522 6725 8528
rect 6826 8519 6832 8531
rect 6884 8519 6890 8571
rect 6667 8358 6725 8364
rect 6667 8324 6679 8358
rect 6713 8355 6725 8358
rect 6826 8355 6832 8367
rect 6713 8327 6832 8355
rect 6713 8324 6725 8327
rect 6667 8318 6725 8324
rect 6826 8315 6832 8327
rect 6884 8315 6890 8367
rect 6667 8154 6725 8160
rect 6667 8120 6679 8154
rect 6713 8151 6725 8154
rect 6826 8151 6832 8163
rect 6713 8123 6832 8151
rect 6713 8120 6725 8123
rect 6667 8114 6725 8120
rect 6826 8111 6832 8123
rect 6884 8111 6890 8163
rect 3691 7943 3697 7995
rect 3749 7943 3755 7995
rect 4087 7943 4093 7995
rect 4145 7943 4151 7995
rect 4697 7943 4703 7995
rect 4755 7943 4761 7995
rect 5945 7943 5951 7995
rect 6003 7943 6009 7995
rect 109 7520 115 7572
rect 167 7520 173 7572
rect 6868 7506 6874 7518
rect 5095 7478 6874 7506
rect 2557 7095 2563 7147
rect 2615 7095 2621 7147
rect 2627 6887 2633 6899
rect 2575 6859 2633 6887
rect 2627 6847 2633 6859
rect 2685 6847 2691 6899
rect 109 6568 115 6620
rect 167 6568 173 6620
rect 2557 6143 2563 6195
rect 2615 6143 2621 6195
rect 109 5531 115 5583
rect 167 5531 173 5583
rect 2557 4909 2563 4961
rect 2615 4909 2621 4961
rect 322 4750 328 4802
rect 380 4750 386 4802
rect 730 4750 736 4802
rect 788 4750 794 4802
rect 1138 4750 1144 4802
rect 1196 4750 1202 4802
rect 1546 4750 1552 4802
rect 1604 4750 1610 4802
rect 1954 4750 1960 4802
rect 2012 4750 2018 4802
rect 2362 4750 2368 4802
rect 2420 4750 2426 4802
rect 5095 4487 5123 7478
rect 6868 7466 6874 7478
rect 6926 7466 6932 7518
rect 6953 7075 6981 7124
rect 7157 7075 7185 7124
rect 7361 7075 7389 7124
rect 7565 7075 7593 7124
rect 7769 7075 7797 7124
rect 7973 7075 8001 7124
rect 8177 7075 8205 7124
rect 8381 7075 8409 7124
rect 8585 7075 8613 7124
rect 8789 7075 8817 7124
rect 8993 7075 9021 7124
rect 9197 7075 9225 7124
rect 9401 7075 9429 7124
rect 9605 7075 9633 7124
rect 9809 7075 9837 7124
rect 10013 7075 10041 7124
rect 10217 7075 10245 7124
rect 10421 7075 10449 7124
rect 10625 7075 10653 7124
rect 10829 7075 10857 7124
rect 11033 7075 11061 7124
rect 11237 7075 11265 7124
rect 11441 7075 11469 7124
rect 11645 7075 11673 7124
rect 11849 7075 11877 7124
rect 12053 7075 12081 7124
rect 12257 7075 12285 7124
rect 12461 7075 12489 7124
rect 12665 7075 12693 7124
rect 12869 7075 12897 7124
rect 13073 7075 13101 7124
rect 13277 7075 13305 7124
rect 13481 7075 13509 7124
rect 13685 7075 13713 7124
rect 13889 7075 13917 7124
rect 14093 7075 14121 7124
rect 14297 7075 14325 7124
rect 14501 7075 14529 7124
rect 14705 7075 14733 7124
rect 14909 7075 14937 7124
rect 15113 7075 15141 7124
rect 15317 7075 15345 7124
rect 15521 7075 15549 7124
rect 15725 7075 15753 7124
rect 15929 7075 15957 7124
rect 16133 7075 16161 7124
rect 16337 7075 16365 7124
rect 16541 7075 16569 7124
rect 6944 7063 6990 7075
rect 6944 7029 6950 7063
rect 6984 7029 6990 7063
rect 6944 7017 6990 7029
rect 7148 7063 7194 7075
rect 7148 7029 7154 7063
rect 7188 7029 7194 7063
rect 7148 7017 7194 7029
rect 7352 7063 7398 7075
rect 7352 7029 7358 7063
rect 7392 7029 7398 7063
rect 7352 7017 7398 7029
rect 7556 7063 7602 7075
rect 7556 7029 7562 7063
rect 7596 7029 7602 7063
rect 7556 7017 7602 7029
rect 7760 7063 7806 7075
rect 7760 7029 7766 7063
rect 7800 7029 7806 7063
rect 7760 7017 7806 7029
rect 7964 7063 8010 7075
rect 7964 7029 7970 7063
rect 8004 7029 8010 7063
rect 7964 7017 8010 7029
rect 8168 7063 8214 7075
rect 8168 7029 8174 7063
rect 8208 7029 8214 7063
rect 8168 7017 8214 7029
rect 8372 7063 8418 7075
rect 8372 7029 8378 7063
rect 8412 7029 8418 7063
rect 8372 7017 8418 7029
rect 8576 7063 8622 7075
rect 8576 7029 8582 7063
rect 8616 7029 8622 7063
rect 8576 7017 8622 7029
rect 8780 7063 8826 7075
rect 8780 7029 8786 7063
rect 8820 7029 8826 7063
rect 8780 7017 8826 7029
rect 8984 7063 9030 7075
rect 8984 7029 8990 7063
rect 9024 7029 9030 7063
rect 8984 7017 9030 7029
rect 9188 7063 9234 7075
rect 9188 7029 9194 7063
rect 9228 7029 9234 7063
rect 9188 7017 9234 7029
rect 9392 7063 9438 7075
rect 9392 7029 9398 7063
rect 9432 7029 9438 7063
rect 9392 7017 9438 7029
rect 9596 7063 9642 7075
rect 9596 7029 9602 7063
rect 9636 7029 9642 7063
rect 9596 7017 9642 7029
rect 9800 7063 9846 7075
rect 9800 7029 9806 7063
rect 9840 7029 9846 7063
rect 9800 7017 9846 7029
rect 10004 7063 10050 7075
rect 10004 7029 10010 7063
rect 10044 7029 10050 7063
rect 10004 7017 10050 7029
rect 10208 7063 10254 7075
rect 10208 7029 10214 7063
rect 10248 7029 10254 7063
rect 10208 7017 10254 7029
rect 10412 7063 10458 7075
rect 10412 7029 10418 7063
rect 10452 7029 10458 7063
rect 10412 7017 10458 7029
rect 10616 7063 10662 7075
rect 10616 7029 10622 7063
rect 10656 7029 10662 7063
rect 10616 7017 10662 7029
rect 10820 7063 10866 7075
rect 10820 7029 10826 7063
rect 10860 7029 10866 7063
rect 10820 7017 10866 7029
rect 11024 7063 11070 7075
rect 11024 7029 11030 7063
rect 11064 7029 11070 7063
rect 11024 7017 11070 7029
rect 11228 7063 11274 7075
rect 11228 7029 11234 7063
rect 11268 7029 11274 7063
rect 11228 7017 11274 7029
rect 11432 7063 11478 7075
rect 11432 7029 11438 7063
rect 11472 7029 11478 7063
rect 11432 7017 11478 7029
rect 11636 7063 11682 7075
rect 11636 7029 11642 7063
rect 11676 7029 11682 7063
rect 11636 7017 11682 7029
rect 11840 7063 11886 7075
rect 11840 7029 11846 7063
rect 11880 7029 11886 7063
rect 11840 7017 11886 7029
rect 12044 7063 12090 7075
rect 12044 7029 12050 7063
rect 12084 7029 12090 7063
rect 12044 7017 12090 7029
rect 12248 7063 12294 7075
rect 12248 7029 12254 7063
rect 12288 7029 12294 7063
rect 12248 7017 12294 7029
rect 12452 7063 12498 7075
rect 12452 7029 12458 7063
rect 12492 7029 12498 7063
rect 12452 7017 12498 7029
rect 12656 7063 12702 7075
rect 12656 7029 12662 7063
rect 12696 7029 12702 7063
rect 12656 7017 12702 7029
rect 12860 7063 12906 7075
rect 12860 7029 12866 7063
rect 12900 7029 12906 7063
rect 12860 7017 12906 7029
rect 13064 7063 13110 7075
rect 13064 7029 13070 7063
rect 13104 7029 13110 7063
rect 13064 7017 13110 7029
rect 13268 7063 13314 7075
rect 13268 7029 13274 7063
rect 13308 7029 13314 7063
rect 13268 7017 13314 7029
rect 13472 7063 13518 7075
rect 13472 7029 13478 7063
rect 13512 7029 13518 7063
rect 13472 7017 13518 7029
rect 13676 7063 13722 7075
rect 13676 7029 13682 7063
rect 13716 7029 13722 7063
rect 13676 7017 13722 7029
rect 13880 7063 13926 7075
rect 13880 7029 13886 7063
rect 13920 7029 13926 7063
rect 13880 7017 13926 7029
rect 14084 7063 14130 7075
rect 14084 7029 14090 7063
rect 14124 7029 14130 7063
rect 14084 7017 14130 7029
rect 14288 7063 14334 7075
rect 14288 7029 14294 7063
rect 14328 7029 14334 7063
rect 14288 7017 14334 7029
rect 14492 7063 14538 7075
rect 14492 7029 14498 7063
rect 14532 7029 14538 7063
rect 14492 7017 14538 7029
rect 14696 7063 14742 7075
rect 14696 7029 14702 7063
rect 14736 7029 14742 7063
rect 14696 7017 14742 7029
rect 14900 7063 14946 7075
rect 14900 7029 14906 7063
rect 14940 7029 14946 7063
rect 14900 7017 14946 7029
rect 15104 7063 15150 7075
rect 15104 7029 15110 7063
rect 15144 7029 15150 7063
rect 15104 7017 15150 7029
rect 15308 7063 15354 7075
rect 15308 7029 15314 7063
rect 15348 7029 15354 7063
rect 15308 7017 15354 7029
rect 15512 7063 15558 7075
rect 15512 7029 15518 7063
rect 15552 7029 15558 7063
rect 15512 7017 15558 7029
rect 15716 7063 15762 7075
rect 15716 7029 15722 7063
rect 15756 7029 15762 7063
rect 15716 7017 15762 7029
rect 15920 7063 15966 7075
rect 15920 7029 15926 7063
rect 15960 7029 15966 7063
rect 15920 7017 15966 7029
rect 16124 7063 16170 7075
rect 16124 7029 16130 7063
rect 16164 7029 16170 7063
rect 16124 7017 16170 7029
rect 16328 7063 16374 7075
rect 16328 7029 16334 7063
rect 16368 7029 16374 7063
rect 16328 7017 16374 7029
rect 16532 7063 16578 7075
rect 16532 7029 16538 7063
rect 16572 7029 16578 7063
rect 16532 7017 16578 7029
rect 6815 6428 6821 6480
rect 6873 6428 6879 6480
rect 16607 6428 16613 6480
rect 16665 6428 16671 6480
rect 6815 5512 6821 5564
rect 6873 5512 6879 5564
rect 16607 5512 16613 5564
rect 16665 5512 16671 5564
rect 6944 5468 6990 5480
rect 6944 5434 6950 5468
rect 6984 5434 6990 5468
rect 6944 5422 6990 5434
rect 7148 5468 7194 5480
rect 7148 5434 7154 5468
rect 7188 5434 7194 5468
rect 7148 5422 7194 5434
rect 7352 5468 7398 5480
rect 7352 5434 7358 5468
rect 7392 5434 7398 5468
rect 7352 5422 7398 5434
rect 7556 5468 7602 5480
rect 7556 5434 7562 5468
rect 7596 5434 7602 5468
rect 7556 5422 7602 5434
rect 7760 5468 7806 5480
rect 7760 5434 7766 5468
rect 7800 5434 7806 5468
rect 7760 5422 7806 5434
rect 7964 5468 8010 5480
rect 7964 5434 7970 5468
rect 8004 5434 8010 5468
rect 7964 5422 8010 5434
rect 8168 5468 8214 5480
rect 8168 5434 8174 5468
rect 8208 5434 8214 5468
rect 8168 5422 8214 5434
rect 8372 5468 8418 5480
rect 8372 5434 8378 5468
rect 8412 5434 8418 5468
rect 8372 5422 8418 5434
rect 8576 5468 8622 5480
rect 8576 5434 8582 5468
rect 8616 5434 8622 5468
rect 8576 5422 8622 5434
rect 8780 5468 8826 5480
rect 8780 5434 8786 5468
rect 8820 5434 8826 5468
rect 8780 5422 8826 5434
rect 8984 5468 9030 5480
rect 8984 5434 8990 5468
rect 9024 5434 9030 5468
rect 8984 5422 9030 5434
rect 9188 5468 9234 5480
rect 9188 5434 9194 5468
rect 9228 5434 9234 5468
rect 9188 5422 9234 5434
rect 9392 5468 9438 5480
rect 9392 5434 9398 5468
rect 9432 5434 9438 5468
rect 9392 5422 9438 5434
rect 9596 5468 9642 5480
rect 9596 5434 9602 5468
rect 9636 5434 9642 5468
rect 9596 5422 9642 5434
rect 9800 5468 9846 5480
rect 9800 5434 9806 5468
rect 9840 5434 9846 5468
rect 9800 5422 9846 5434
rect 10004 5468 10050 5480
rect 10004 5434 10010 5468
rect 10044 5434 10050 5468
rect 10004 5422 10050 5434
rect 10208 5468 10254 5480
rect 10208 5434 10214 5468
rect 10248 5434 10254 5468
rect 10208 5422 10254 5434
rect 10412 5468 10458 5480
rect 10412 5434 10418 5468
rect 10452 5434 10458 5468
rect 10412 5422 10458 5434
rect 10616 5468 10662 5480
rect 10616 5434 10622 5468
rect 10656 5434 10662 5468
rect 10616 5422 10662 5434
rect 10820 5468 10866 5480
rect 10820 5434 10826 5468
rect 10860 5434 10866 5468
rect 10820 5422 10866 5434
rect 11024 5468 11070 5480
rect 11024 5434 11030 5468
rect 11064 5434 11070 5468
rect 11024 5422 11070 5434
rect 11228 5468 11274 5480
rect 11228 5434 11234 5468
rect 11268 5434 11274 5468
rect 11228 5422 11274 5434
rect 11432 5468 11478 5480
rect 11432 5434 11438 5468
rect 11472 5434 11478 5468
rect 11432 5422 11478 5434
rect 11636 5468 11682 5480
rect 11636 5434 11642 5468
rect 11676 5434 11682 5468
rect 11636 5422 11682 5434
rect 11840 5468 11886 5480
rect 11840 5434 11846 5468
rect 11880 5434 11886 5468
rect 11840 5422 11886 5434
rect 12044 5468 12090 5480
rect 12044 5434 12050 5468
rect 12084 5434 12090 5468
rect 12044 5422 12090 5434
rect 12248 5468 12294 5480
rect 12248 5434 12254 5468
rect 12288 5434 12294 5468
rect 12248 5422 12294 5434
rect 12452 5468 12498 5480
rect 12452 5434 12458 5468
rect 12492 5434 12498 5468
rect 12452 5422 12498 5434
rect 12656 5468 12702 5480
rect 12656 5434 12662 5468
rect 12696 5434 12702 5468
rect 12656 5422 12702 5434
rect 12860 5468 12906 5480
rect 12860 5434 12866 5468
rect 12900 5434 12906 5468
rect 12860 5422 12906 5434
rect 13064 5468 13110 5480
rect 13064 5434 13070 5468
rect 13104 5434 13110 5468
rect 13064 5422 13110 5434
rect 13268 5468 13314 5480
rect 13268 5434 13274 5468
rect 13308 5434 13314 5468
rect 13268 5422 13314 5434
rect 13472 5468 13518 5480
rect 13472 5434 13478 5468
rect 13512 5434 13518 5468
rect 13472 5422 13518 5434
rect 13676 5468 13722 5480
rect 13676 5434 13682 5468
rect 13716 5434 13722 5468
rect 13676 5422 13722 5434
rect 13880 5468 13926 5480
rect 13880 5434 13886 5468
rect 13920 5434 13926 5468
rect 13880 5422 13926 5434
rect 14084 5468 14130 5480
rect 14084 5434 14090 5468
rect 14124 5434 14130 5468
rect 14084 5422 14130 5434
rect 14288 5468 14334 5480
rect 14288 5434 14294 5468
rect 14328 5434 14334 5468
rect 14288 5422 14334 5434
rect 14492 5468 14538 5480
rect 14492 5434 14498 5468
rect 14532 5434 14538 5468
rect 14492 5422 14538 5434
rect 14696 5468 14742 5480
rect 14696 5434 14702 5468
rect 14736 5434 14742 5468
rect 14696 5422 14742 5434
rect 14900 5468 14946 5480
rect 14900 5434 14906 5468
rect 14940 5434 14946 5468
rect 14900 5422 14946 5434
rect 15104 5468 15150 5480
rect 15104 5434 15110 5468
rect 15144 5434 15150 5468
rect 15104 5422 15150 5434
rect 15308 5468 15354 5480
rect 15308 5434 15314 5468
rect 15348 5434 15354 5468
rect 15308 5422 15354 5434
rect 15512 5468 15558 5480
rect 15512 5434 15518 5468
rect 15552 5434 15558 5468
rect 15512 5422 15558 5434
rect 15716 5468 15762 5480
rect 15716 5434 15722 5468
rect 15756 5434 15762 5468
rect 15716 5422 15762 5434
rect 15920 5468 15966 5480
rect 15920 5434 15926 5468
rect 15960 5434 15966 5468
rect 15920 5422 15966 5434
rect 16124 5468 16170 5480
rect 16124 5434 16130 5468
rect 16164 5434 16170 5468
rect 16124 5422 16170 5434
rect 16328 5468 16374 5480
rect 16328 5434 16334 5468
rect 16368 5434 16374 5468
rect 16328 5422 16374 5434
rect 16532 5468 16578 5480
rect 16532 5434 16538 5468
rect 16572 5434 16578 5468
rect 16532 5422 16578 5434
rect 6953 4916 6981 5422
rect 7157 4916 7185 5422
rect 7361 4916 7389 5422
rect 7565 4916 7593 5422
rect 7769 4916 7797 5422
rect 7973 4916 8001 5422
rect 8177 4916 8205 5422
rect 8381 4916 8409 5422
rect 8585 4916 8613 5422
rect 8789 4916 8817 5422
rect 8993 4916 9021 5422
rect 9197 4916 9225 5422
rect 9401 4916 9429 5422
rect 9605 4916 9633 5422
rect 9809 4916 9837 5422
rect 10013 4916 10041 5422
rect 10217 4916 10245 5422
rect 10421 4916 10449 5422
rect 10625 4916 10653 5422
rect 10829 4916 10857 5422
rect 11033 4916 11061 5422
rect 11237 4916 11265 5422
rect 11441 4916 11469 5422
rect 11645 4916 11673 5422
rect 11849 4916 11877 5422
rect 12053 4916 12081 5422
rect 12257 4916 12285 5422
rect 12461 4916 12489 5422
rect 12665 4916 12693 5422
rect 12869 4916 12897 5422
rect 13073 4916 13101 5422
rect 13277 4916 13305 5422
rect 13481 4916 13509 5422
rect 13685 4916 13713 5422
rect 13889 4916 13917 5422
rect 14093 4916 14121 5422
rect 14297 4916 14325 5422
rect 14501 4916 14529 5422
rect 14705 4916 14733 5422
rect 14909 4916 14937 5422
rect 15113 4916 15141 5422
rect 15317 4916 15345 5422
rect 15521 4916 15549 5422
rect 15725 4916 15753 5422
rect 15929 4916 15957 5422
rect 16133 4916 16161 5422
rect 16337 4916 16365 5422
rect 16541 4916 16569 5422
rect 3406 4459 5123 4487
rect 2853 3628 2911 3634
rect 2853 3594 2865 3628
rect 2899 3625 2911 3628
rect 3406 3625 3434 4459
rect 5723 4190 5729 4242
rect 5781 4190 5787 4242
rect 6345 4190 6351 4242
rect 6403 4190 6409 4242
rect 6664 4070 6670 4122
rect 6722 4070 6728 4122
rect 6664 3866 6670 3918
rect 6722 3866 6728 3918
rect 6664 3662 6670 3714
rect 6722 3662 6728 3714
rect 2899 3597 3434 3625
rect 2899 3594 2911 3597
rect 2853 3588 2911 3594
rect 3406 2438 3434 3597
rect 5723 3494 5729 3546
rect 5781 3494 5787 3546
rect 6345 3494 6351 3546
rect 6403 3494 6409 3546
rect 6935 3444 6941 3496
rect 6993 3444 6999 3496
rect 7547 3444 7553 3496
rect 7605 3444 7611 3496
rect 8159 3444 8165 3496
rect 8217 3444 8223 3496
rect 8771 3444 8777 3496
rect 8829 3444 8835 3496
rect 9383 3444 9389 3496
rect 9441 3444 9447 3496
rect 9995 3444 10001 3496
rect 10053 3444 10059 3496
rect 10607 3444 10613 3496
rect 10665 3444 10671 3496
rect 11219 3444 11225 3496
rect 11277 3444 11283 3496
rect 11831 3444 11837 3496
rect 11889 3444 11895 3496
rect 12443 3444 12449 3496
rect 12501 3444 12507 3496
rect 13055 3444 13061 3496
rect 13113 3444 13119 3496
rect 13667 3444 13673 3496
rect 13725 3444 13731 3496
rect 14279 3444 14285 3496
rect 14337 3444 14343 3496
rect 14891 3444 14897 3496
rect 14949 3444 14955 3496
rect 15503 3444 15509 3496
rect 15561 3444 15567 3496
rect 16115 3444 16121 3496
rect 16173 3444 16179 3496
rect 3735 3071 3741 3123
rect 3793 3071 3799 3123
rect 4551 2646 4557 2698
rect 4609 2646 4615 2698
rect 3406 2410 4161 2438
rect 9995 2429 10001 2481
rect 10053 2469 10059 2481
rect 11673 2469 11679 2481
rect 10053 2441 11679 2469
rect 10053 2429 10059 2441
rect 11673 2429 11679 2441
rect 11731 2429 11737 2481
rect 9383 2327 9389 2379
rect 9441 2367 9447 2379
rect 11365 2367 11371 2379
rect 9441 2339 11371 2367
rect 9441 2327 9447 2339
rect 11365 2327 11371 2339
rect 11423 2327 11429 2379
rect 8771 2225 8777 2277
rect 8829 2265 8835 2277
rect 11057 2265 11063 2277
rect 8829 2237 11063 2265
rect 8829 2225 8835 2237
rect 11057 2225 11063 2237
rect 11115 2225 11121 2277
rect 3735 2119 3741 2171
rect 3793 2119 3799 2171
rect 8159 2123 8165 2175
rect 8217 2163 8223 2175
rect 10749 2163 10755 2175
rect 8217 2135 10755 2163
rect 8217 2123 8223 2135
rect 10749 2123 10755 2135
rect 10807 2123 10813 2175
rect 11831 2123 11837 2175
rect 11889 2163 11895 2175
rect 12597 2163 12603 2175
rect 11889 2135 12603 2163
rect 11889 2123 11895 2135
rect 12597 2123 12603 2135
rect 12655 2123 12661 2175
rect 14753 2123 14759 2175
rect 14811 2163 14817 2175
rect 16115 2163 16121 2175
rect 14811 2135 16121 2163
rect 14811 2123 14817 2135
rect 16115 2123 16121 2135
rect 16173 2123 16179 2175
rect 7547 2021 7553 2073
rect 7605 2061 7611 2073
rect 10441 2061 10447 2073
rect 7605 2033 10447 2061
rect 7605 2021 7611 2033
rect 10441 2021 10447 2033
rect 10499 2021 10505 2073
rect 11219 2021 11225 2073
rect 11277 2061 11283 2073
rect 12289 2061 12295 2073
rect 11277 2033 12295 2061
rect 11277 2021 11283 2033
rect 12289 2021 12295 2033
rect 12347 2021 12353 2073
rect 14137 2021 14143 2073
rect 14195 2061 14201 2073
rect 14891 2061 14897 2073
rect 14195 2033 14897 2061
rect 14195 2021 14201 2033
rect 14891 2021 14897 2033
rect 14949 2021 14955 2073
rect 6935 1919 6941 1971
rect 6993 1959 6999 1971
rect 10133 1959 10139 1971
rect 6993 1931 10139 1959
rect 6993 1919 6999 1931
rect 10133 1919 10139 1931
rect 10191 1919 10197 1971
rect 10607 1919 10613 1971
rect 10665 1959 10671 1971
rect 11981 1959 11987 1971
rect 10665 1931 11987 1959
rect 10665 1919 10671 1931
rect 11981 1919 11987 1931
rect 12039 1919 12045 1971
rect 12443 1919 12449 1971
rect 12501 1959 12507 1971
rect 12905 1959 12911 1971
rect 12501 1931 12911 1959
rect 12501 1919 12507 1931
rect 12905 1919 12911 1931
rect 12963 1919 12969 1971
rect 13055 1919 13061 1971
rect 13113 1959 13119 1971
rect 13213 1959 13219 1971
rect 13113 1931 13219 1959
rect 13113 1919 13119 1931
rect 13213 1919 13219 1931
rect 13271 1919 13277 1971
rect 13521 1919 13527 1971
rect 13579 1959 13585 1971
rect 13667 1959 13673 1971
rect 13579 1931 13673 1959
rect 13579 1919 13585 1931
rect 13667 1919 13673 1931
rect 13725 1919 13731 1971
rect 13829 1919 13835 1971
rect 13887 1959 13893 1971
rect 14279 1959 14285 1971
rect 13887 1931 14285 1959
rect 13887 1919 13893 1931
rect 14279 1919 14285 1931
rect 14337 1919 14343 1971
rect 14445 1919 14451 1971
rect 14503 1959 14509 1971
rect 15503 1959 15509 1971
rect 14503 1931 15509 1959
rect 14503 1919 14509 1931
rect 15503 1919 15509 1931
rect 15561 1919 15567 1971
rect 4551 1694 4557 1746
rect 4609 1694 4615 1746
rect 10133 1696 10139 1748
rect 10191 1696 10197 1748
rect 10441 1696 10447 1748
rect 10499 1696 10505 1748
rect 10749 1696 10755 1748
rect 10807 1696 10813 1748
rect 11057 1696 11063 1748
rect 11115 1696 11121 1748
rect 11365 1696 11371 1748
rect 11423 1696 11429 1748
rect 11673 1696 11679 1748
rect 11731 1696 11737 1748
rect 11981 1696 11987 1748
rect 12039 1696 12045 1748
rect 12289 1696 12295 1748
rect 12347 1696 12353 1748
rect 12597 1696 12603 1748
rect 12655 1696 12661 1748
rect 12905 1696 12911 1748
rect 12963 1696 12969 1748
rect 13213 1696 13219 1748
rect 13271 1696 13277 1748
rect 13521 1696 13527 1748
rect 13579 1696 13585 1748
rect 13829 1696 13835 1748
rect 13887 1696 13893 1748
rect 14137 1696 14143 1748
rect 14195 1696 14201 1748
rect 14445 1696 14451 1748
rect 14503 1696 14509 1748
rect 14753 1696 14759 1748
rect 14811 1696 14817 1748
rect 505 1378 511 1430
rect 563 1378 569 1430
rect 9965 1426 9971 1478
rect 10023 1426 10029 1478
rect 14873 1426 14879 1478
rect 14931 1426 14937 1478
rect 2482 1366 2488 1418
rect 2540 1366 2546 1418
rect 3735 1082 3741 1134
rect 3793 1082 3799 1134
rect 3105 627 3111 679
rect 3163 627 3169 679
rect 4551 460 4557 512
rect 4609 460 4615 512
rect 9965 510 9971 562
rect 10023 510 10029 562
rect 14873 510 14879 562
rect 14931 510 14937 562
rect 3948 301 3954 353
rect 4006 301 4012 353
rect 4356 301 4362 353
rect 4414 301 4420 353
rect 10139 43 10191 49
rect 10139 -15 10191 -9
rect 10447 43 10499 49
rect 10447 -15 10499 -9
rect 10755 43 10807 49
rect 10755 -15 10807 -9
rect 11063 43 11115 49
rect 11063 -15 11115 -9
rect 11371 43 11423 49
rect 11371 -15 11423 -9
rect 11679 43 11731 49
rect 11679 -15 11731 -9
rect 11987 43 12039 49
rect 11987 -15 12039 -9
rect 12295 43 12347 49
rect 12295 -15 12347 -9
rect 12603 43 12655 49
rect 12603 -15 12655 -9
rect 12911 43 12963 49
rect 12911 -15 12963 -9
rect 13219 43 13271 49
rect 13219 -15 13271 -9
rect 13527 43 13579 49
rect 13527 -15 13579 -9
rect 13835 43 13887 49
rect 13835 -15 13887 -9
rect 14143 43 14195 49
rect 14143 -15 14195 -9
rect 14451 43 14503 49
rect 14451 -15 14503 -9
rect 14759 43 14811 49
rect 14759 -15 14811 -9
<< via1 >>
rect 6927 17326 6979 17378
rect 16543 17326 16595 17378
rect 3697 17115 3749 17167
rect 4093 17115 4145 17167
rect 4703 17115 4755 17167
rect 5951 17115 6003 17167
rect 6832 16995 6884 17047
rect 6832 16791 6884 16843
rect 6832 16483 6884 16535
rect 6832 16279 6884 16331
rect 6832 16075 6884 16127
rect 6832 15871 6884 15923
rect 6832 15667 6884 15719
rect 6832 15463 6884 15515
rect 6832 15259 6884 15311
rect 6832 15055 6884 15107
rect 6832 14747 6884 14799
rect 6832 14543 6884 14595
rect 6832 14339 6884 14391
rect 6832 14135 6884 14187
rect 6832 13931 6884 13983
rect 6832 13727 6884 13779
rect 6832 13523 6884 13575
rect 6832 13319 6884 13371
rect 6832 13011 6884 13063
rect 6832 12807 6884 12859
rect 6832 12603 6884 12655
rect 6832 12399 6884 12451
rect 6832 12195 6884 12247
rect 6832 11991 6884 12043
rect 6832 11787 6884 11839
rect 6832 11583 6884 11635
rect 6832 11275 6884 11327
rect 6832 11071 6884 11123
rect 6832 10867 6884 10919
rect 6832 10663 6884 10715
rect 6832 10459 6884 10511
rect 6832 10255 6884 10307
rect 6832 10051 6884 10103
rect 6832 9847 6884 9899
rect 6832 9539 6884 9591
rect 6832 9335 6884 9387
rect 6832 9131 6884 9183
rect 6832 8927 6884 8979
rect 6832 8723 6884 8775
rect 6832 8519 6884 8571
rect 6832 8315 6884 8367
rect 6832 8111 6884 8163
rect 3697 7943 3749 7995
rect 4093 7943 4145 7995
rect 4703 7943 4755 7995
rect 5951 7943 6003 7995
rect 115 7520 167 7572
rect 2563 7095 2615 7147
rect 2633 6847 2685 6899
rect 115 6568 167 6620
rect 2563 6143 2615 6195
rect 115 5531 167 5583
rect 2563 4909 2615 4961
rect 328 4793 380 4802
rect 328 4759 337 4793
rect 337 4759 371 4793
rect 371 4759 380 4793
rect 328 4750 380 4759
rect 736 4793 788 4802
rect 736 4759 745 4793
rect 745 4759 779 4793
rect 779 4759 788 4793
rect 736 4750 788 4759
rect 1144 4793 1196 4802
rect 1144 4759 1153 4793
rect 1153 4759 1187 4793
rect 1187 4759 1196 4793
rect 1144 4750 1196 4759
rect 1552 4793 1604 4802
rect 1552 4759 1561 4793
rect 1561 4759 1595 4793
rect 1595 4759 1604 4793
rect 1552 4750 1604 4759
rect 1960 4793 2012 4802
rect 1960 4759 1969 4793
rect 1969 4759 2003 4793
rect 2003 4759 2012 4793
rect 1960 4750 2012 4759
rect 2368 4793 2420 4802
rect 2368 4759 2377 4793
rect 2377 4759 2411 4793
rect 2411 4759 2420 4793
rect 2368 4750 2420 4759
rect 6874 7466 6926 7518
rect 6821 6428 6873 6480
rect 16613 6428 16665 6480
rect 6821 5512 6873 5564
rect 16613 5512 16665 5564
rect 5729 4190 5781 4242
rect 6351 4190 6403 4242
rect 6670 4113 6722 4122
rect 6670 4079 6679 4113
rect 6679 4079 6713 4113
rect 6713 4079 6722 4113
rect 6670 4070 6722 4079
rect 6670 3909 6722 3918
rect 6670 3875 6679 3909
rect 6679 3875 6713 3909
rect 6713 3875 6722 3909
rect 6670 3866 6722 3875
rect 6670 3705 6722 3714
rect 6670 3671 6679 3705
rect 6679 3671 6713 3705
rect 6713 3671 6722 3705
rect 6670 3662 6722 3671
rect 5729 3494 5781 3546
rect 6351 3494 6403 3546
rect 6941 3444 6993 3496
rect 7553 3444 7605 3496
rect 8165 3444 8217 3496
rect 8777 3444 8829 3496
rect 9389 3444 9441 3496
rect 10001 3444 10053 3496
rect 10613 3444 10665 3496
rect 11225 3444 11277 3496
rect 11837 3444 11889 3496
rect 12449 3444 12501 3496
rect 13061 3444 13113 3496
rect 13673 3444 13725 3496
rect 14285 3444 14337 3496
rect 14897 3444 14949 3496
rect 15509 3444 15561 3496
rect 16121 3444 16173 3496
rect 3741 3071 3793 3123
rect 4557 2646 4609 2698
rect 10001 2429 10053 2481
rect 11679 2429 11731 2481
rect 9389 2327 9441 2379
rect 11371 2327 11423 2379
rect 8777 2225 8829 2277
rect 11063 2225 11115 2277
rect 3741 2119 3793 2171
rect 8165 2123 8217 2175
rect 10755 2123 10807 2175
rect 11837 2123 11889 2175
rect 12603 2123 12655 2175
rect 14759 2123 14811 2175
rect 16121 2123 16173 2175
rect 7553 2021 7605 2073
rect 10447 2021 10499 2073
rect 11225 2021 11277 2073
rect 12295 2021 12347 2073
rect 14143 2021 14195 2073
rect 14897 2021 14949 2073
rect 6941 1919 6993 1971
rect 10139 1919 10191 1971
rect 10613 1919 10665 1971
rect 11987 1919 12039 1971
rect 12449 1919 12501 1971
rect 12911 1919 12963 1971
rect 13061 1919 13113 1971
rect 13219 1919 13271 1971
rect 13527 1919 13579 1971
rect 13673 1919 13725 1971
rect 13835 1919 13887 1971
rect 14285 1919 14337 1971
rect 14451 1919 14503 1971
rect 15509 1919 15561 1971
rect 4557 1694 4609 1746
rect 10139 1739 10191 1748
rect 10139 1705 10148 1739
rect 10148 1705 10182 1739
rect 10182 1705 10191 1739
rect 10139 1696 10191 1705
rect 10447 1739 10499 1748
rect 10447 1705 10456 1739
rect 10456 1705 10490 1739
rect 10490 1705 10499 1739
rect 10447 1696 10499 1705
rect 10755 1739 10807 1748
rect 10755 1705 10764 1739
rect 10764 1705 10798 1739
rect 10798 1705 10807 1739
rect 10755 1696 10807 1705
rect 11063 1739 11115 1748
rect 11063 1705 11072 1739
rect 11072 1705 11106 1739
rect 11106 1705 11115 1739
rect 11063 1696 11115 1705
rect 11371 1739 11423 1748
rect 11371 1705 11380 1739
rect 11380 1705 11414 1739
rect 11414 1705 11423 1739
rect 11371 1696 11423 1705
rect 11679 1739 11731 1748
rect 11679 1705 11688 1739
rect 11688 1705 11722 1739
rect 11722 1705 11731 1739
rect 11679 1696 11731 1705
rect 11987 1739 12039 1748
rect 11987 1705 11996 1739
rect 11996 1705 12030 1739
rect 12030 1705 12039 1739
rect 11987 1696 12039 1705
rect 12295 1739 12347 1748
rect 12295 1705 12304 1739
rect 12304 1705 12338 1739
rect 12338 1705 12347 1739
rect 12295 1696 12347 1705
rect 12603 1739 12655 1748
rect 12603 1705 12612 1739
rect 12612 1705 12646 1739
rect 12646 1705 12655 1739
rect 12603 1696 12655 1705
rect 12911 1739 12963 1748
rect 12911 1705 12920 1739
rect 12920 1705 12954 1739
rect 12954 1705 12963 1739
rect 12911 1696 12963 1705
rect 13219 1739 13271 1748
rect 13219 1705 13228 1739
rect 13228 1705 13262 1739
rect 13262 1705 13271 1739
rect 13219 1696 13271 1705
rect 13527 1739 13579 1748
rect 13527 1705 13536 1739
rect 13536 1705 13570 1739
rect 13570 1705 13579 1739
rect 13527 1696 13579 1705
rect 13835 1739 13887 1748
rect 13835 1705 13844 1739
rect 13844 1705 13878 1739
rect 13878 1705 13887 1739
rect 13835 1696 13887 1705
rect 14143 1739 14195 1748
rect 14143 1705 14152 1739
rect 14152 1705 14186 1739
rect 14186 1705 14195 1739
rect 14143 1696 14195 1705
rect 14451 1739 14503 1748
rect 14451 1705 14460 1739
rect 14460 1705 14494 1739
rect 14494 1705 14503 1739
rect 14451 1696 14503 1705
rect 14759 1739 14811 1748
rect 14759 1705 14768 1739
rect 14768 1705 14802 1739
rect 14802 1705 14811 1739
rect 14759 1696 14811 1705
rect 511 1421 563 1430
rect 511 1387 520 1421
rect 520 1387 554 1421
rect 554 1387 563 1421
rect 511 1378 563 1387
rect 9971 1426 10023 1478
rect 14879 1426 14931 1478
rect 2488 1409 2540 1418
rect 2488 1375 2497 1409
rect 2497 1375 2531 1409
rect 2531 1375 2540 1409
rect 2488 1366 2540 1375
rect 3741 1082 3793 1134
rect 3111 670 3163 679
rect 3111 636 3120 670
rect 3120 636 3154 670
rect 3154 636 3163 670
rect 3111 627 3163 636
rect 4557 460 4609 512
rect 9971 510 10023 562
rect 14879 510 14931 562
rect 3954 344 4006 353
rect 3954 310 3963 344
rect 3963 310 3997 344
rect 3997 310 4006 344
rect 3954 301 4006 310
rect 4362 344 4414 353
rect 4362 310 4371 344
rect 4371 310 4405 344
rect 4405 310 4414 344
rect 4362 301 4414 310
rect 10139 34 10191 43
rect 10139 0 10148 34
rect 10148 0 10182 34
rect 10182 0 10191 34
rect 10139 -9 10191 0
rect 10447 34 10499 43
rect 10447 0 10456 34
rect 10456 0 10490 34
rect 10490 0 10499 34
rect 10447 -9 10499 0
rect 10755 34 10807 43
rect 10755 0 10764 34
rect 10764 0 10798 34
rect 10798 0 10807 34
rect 10755 -9 10807 0
rect 11063 34 11115 43
rect 11063 0 11072 34
rect 11072 0 11106 34
rect 11106 0 11115 34
rect 11063 -9 11115 0
rect 11371 34 11423 43
rect 11371 0 11380 34
rect 11380 0 11414 34
rect 11414 0 11423 34
rect 11371 -9 11423 0
rect 11679 34 11731 43
rect 11679 0 11688 34
rect 11688 0 11722 34
rect 11722 0 11731 34
rect 11679 -9 11731 0
rect 11987 34 12039 43
rect 11987 0 11996 34
rect 11996 0 12030 34
rect 12030 0 12039 34
rect 11987 -9 12039 0
rect 12295 34 12347 43
rect 12295 0 12304 34
rect 12304 0 12338 34
rect 12338 0 12347 34
rect 12295 -9 12347 0
rect 12603 34 12655 43
rect 12603 0 12612 34
rect 12612 0 12646 34
rect 12646 0 12655 34
rect 12603 -9 12655 0
rect 12911 34 12963 43
rect 12911 0 12920 34
rect 12920 0 12954 34
rect 12954 0 12963 34
rect 12911 -9 12963 0
rect 13219 34 13271 43
rect 13219 0 13228 34
rect 13228 0 13262 34
rect 13262 0 13271 34
rect 13219 -9 13271 0
rect 13527 34 13579 43
rect 13527 0 13536 34
rect 13536 0 13570 34
rect 13570 0 13579 34
rect 13527 -9 13579 0
rect 13835 34 13887 43
rect 13835 0 13844 34
rect 13844 0 13878 34
rect 13878 0 13887 34
rect 13835 -9 13887 0
rect 14143 34 14195 43
rect 14143 0 14152 34
rect 14152 0 14186 34
rect 14186 0 14195 34
rect 14143 -9 14195 0
rect 14451 34 14503 43
rect 14451 0 14460 34
rect 14460 0 14494 34
rect 14494 0 14503 34
rect 14451 -9 14503 0
rect 14759 34 14811 43
rect 14759 0 14768 34
rect 14768 0 14802 34
rect 14802 0 14811 34
rect 14759 -9 14811 0
<< metal2 >>
rect 6925 17380 6981 17389
rect 6925 17315 6981 17324
rect 16541 17380 16597 17389
rect 16541 17315 16597 17324
rect 3695 17169 3751 17178
rect 3695 17104 3751 17113
rect 4091 17169 4147 17178
rect 4091 17104 4147 17113
rect 4701 17169 4757 17178
rect 4701 17104 4757 17113
rect 5949 17169 6005 17178
rect 5949 17104 6005 17113
rect 6832 17047 6884 17053
rect 6826 17000 6832 17043
rect 6884 17000 6890 17043
rect 6832 16989 6884 16995
rect 6832 16843 6884 16849
rect 6826 16796 6832 16839
rect 6884 16796 6890 16839
rect 6832 16785 6884 16791
rect 11842 16691 11898 16700
rect 11842 16626 11898 16635
rect 6832 16535 6884 16541
rect 6826 16488 6832 16531
rect 6884 16488 6890 16531
rect 6832 16477 6884 16483
rect 6832 16331 6884 16337
rect 6826 16284 6832 16327
rect 6884 16284 6890 16327
rect 6832 16273 6884 16279
rect 6832 16127 6884 16133
rect 6826 16080 6832 16123
rect 6884 16080 6890 16123
rect 6832 16069 6884 16075
rect 6832 15923 6884 15929
rect 6826 15876 6832 15919
rect 6884 15876 6890 15919
rect 6832 15865 6884 15871
rect 6832 15719 6884 15725
rect 6826 15672 6832 15715
rect 6884 15672 6890 15715
rect 6832 15661 6884 15667
rect 6832 15515 6884 15521
rect 6826 15468 6832 15511
rect 6884 15468 6890 15511
rect 6832 15457 6884 15463
rect 6832 15311 6884 15317
rect 6826 15264 6832 15307
rect 6884 15264 6890 15307
rect 6832 15253 6884 15259
rect 6832 15107 6884 15113
rect 6826 15060 6832 15103
rect 6884 15060 6890 15103
rect 6832 15049 6884 15055
rect 11842 14955 11898 14964
rect 11842 14890 11898 14899
rect 6832 14799 6884 14805
rect 6826 14752 6832 14795
rect 6884 14752 6890 14795
rect 6832 14741 6884 14747
rect 6832 14595 6884 14601
rect 6826 14548 6832 14591
rect 6884 14548 6890 14591
rect 6832 14537 6884 14543
rect 6832 14391 6884 14397
rect 6826 14344 6832 14387
rect 6884 14344 6890 14387
rect 6832 14333 6884 14339
rect 6832 14187 6884 14193
rect 6826 14140 6832 14183
rect 6884 14140 6890 14183
rect 6832 14129 6884 14135
rect 6832 13983 6884 13989
rect 6826 13936 6832 13979
rect 6884 13936 6890 13979
rect 6832 13925 6884 13931
rect 6832 13779 6884 13785
rect 6826 13732 6832 13775
rect 6884 13732 6890 13775
rect 6832 13721 6884 13727
rect 6832 13575 6884 13581
rect 6826 13528 6832 13571
rect 6884 13528 6890 13571
rect 6832 13517 6884 13523
rect 6832 13371 6884 13377
rect 6826 13324 6832 13367
rect 6884 13324 6890 13367
rect 6832 13313 6884 13319
rect 11842 13219 11898 13228
rect 11842 13154 11898 13163
rect 6832 13063 6884 13069
rect 6826 13016 6832 13059
rect 6884 13016 6890 13059
rect 6832 13005 6884 13011
rect 6832 12859 6884 12865
rect 6826 12812 6832 12855
rect 6884 12812 6890 12855
rect 6832 12801 6884 12807
rect 6832 12655 6884 12661
rect 6826 12608 6832 12651
rect 6884 12608 6890 12651
rect 6832 12597 6884 12603
rect 6832 12451 6884 12457
rect 6826 12404 6832 12447
rect 6884 12404 6890 12447
rect 6832 12393 6884 12399
rect 6832 12247 6884 12253
rect 6826 12200 6832 12243
rect 6884 12200 6890 12243
rect 6832 12189 6884 12195
rect 6832 12043 6884 12049
rect 6826 11996 6832 12039
rect 6884 11996 6890 12039
rect 6832 11985 6884 11991
rect 6832 11839 6884 11845
rect 6826 11792 6832 11835
rect 6884 11792 6890 11835
rect 6832 11781 6884 11787
rect 6832 11635 6884 11641
rect 6826 11588 6832 11631
rect 6884 11588 6890 11631
rect 6832 11577 6884 11583
rect 11842 11483 11898 11492
rect 11842 11418 11898 11427
rect 6832 11327 6884 11333
rect 6826 11280 6832 11323
rect 6884 11280 6890 11323
rect 6832 11269 6884 11275
rect 6832 11123 6884 11129
rect 6826 11076 6832 11119
rect 6884 11076 6890 11119
rect 6832 11065 6884 11071
rect 6832 10919 6884 10925
rect 6826 10872 6832 10915
rect 6884 10872 6890 10915
rect 6832 10861 6884 10867
rect 6832 10715 6884 10721
rect 6826 10668 6832 10711
rect 6884 10668 6890 10711
rect 6832 10657 6884 10663
rect 6832 10511 6884 10517
rect 6826 10464 6832 10507
rect 6884 10464 6890 10507
rect 6832 10453 6884 10459
rect 6832 10307 6884 10313
rect 6826 10260 6832 10303
rect 6884 10260 6890 10303
rect 6832 10249 6884 10255
rect 6832 10103 6884 10109
rect 6826 10056 6832 10099
rect 6884 10056 6890 10099
rect 6832 10045 6884 10051
rect 6832 9899 6884 9905
rect 6826 9852 6832 9895
rect 6884 9852 6890 9895
rect 6832 9841 6884 9847
rect 11842 9747 11898 9756
rect 11842 9682 11898 9691
rect 6832 9591 6884 9597
rect 6826 9544 6832 9587
rect 6884 9544 6890 9587
rect 6832 9533 6884 9539
rect 6832 9387 6884 9393
rect 6826 9340 6832 9383
rect 6884 9340 6890 9383
rect 6832 9329 6884 9335
rect 6832 9183 6884 9189
rect 6826 9136 6832 9179
rect 6884 9136 6890 9179
rect 6832 9125 6884 9131
rect 6832 8979 6884 8985
rect 6826 8932 6832 8975
rect 6884 8932 6890 8975
rect 6832 8921 6884 8927
rect 6832 8775 6884 8781
rect 6826 8728 6832 8771
rect 6884 8728 6890 8771
rect 6832 8717 6884 8723
rect 6832 8571 6884 8577
rect 6826 8524 6832 8567
rect 6884 8524 6890 8567
rect 6832 8513 6884 8519
rect 6832 8367 6884 8373
rect 6826 8320 6832 8363
rect 6884 8320 6890 8363
rect 6832 8309 6884 8315
rect 6832 8163 6884 8169
rect 6826 8116 6832 8159
rect 6884 8116 6890 8159
rect 6832 8105 6884 8111
rect 11842 8011 11898 8020
rect 3695 7997 3751 8006
rect 2645 7952 3129 7980
rect 113 7574 169 7583
rect 113 7509 169 7518
rect 2561 7149 2617 7158
rect 2561 7084 2617 7093
rect 2645 6905 2673 7952
rect 3469 7945 3525 7954
rect 3695 7932 3751 7941
rect 4091 7997 4147 8006
rect 4091 7932 4147 7941
rect 4701 7997 4757 8006
rect 4701 7932 4757 7941
rect 5949 7997 6005 8006
rect 11842 7946 11898 7955
rect 5949 7932 6005 7941
rect 3469 7880 3525 7889
rect 6874 7518 6926 7524
rect 6874 7460 6926 7466
rect 6823 7138 6879 7147
rect 6823 7073 6879 7082
rect 2633 6899 2685 6905
rect 2685 6859 3480 6887
rect 2633 6841 2685 6847
rect 113 6622 169 6631
rect 113 6557 169 6566
rect 2561 6197 2617 6206
rect 2561 6132 2617 6141
rect 113 5585 169 5594
rect 113 5520 169 5529
rect 2561 4963 2617 4972
rect 2561 4898 2617 4907
rect 326 4804 382 4813
rect 326 4739 382 4748
rect 734 4804 790 4813
rect 734 4739 790 4748
rect 1142 4804 1198 4813
rect 1142 4739 1198 4748
rect 1550 4804 1606 4813
rect 1550 4739 1606 4748
rect 1958 4804 2014 4813
rect 1958 4739 2014 4748
rect 2366 4804 2422 4813
rect 2366 4739 2422 4748
rect 509 1432 565 1441
rect 509 1367 565 1376
rect 2488 1418 2540 1424
rect 3452 1406 3480 6859
rect 6819 6482 6875 6491
rect 6819 6417 6875 6426
rect 16611 6482 16667 6491
rect 16611 6417 16667 6426
rect 6819 5566 6875 5575
rect 6819 5501 6875 5510
rect 16611 5566 16667 5575
rect 16611 5501 16667 5510
rect 11774 5064 11830 5073
rect 11774 4999 11830 5008
rect 5727 4244 5783 4253
rect 5727 4179 5783 4188
rect 6349 4244 6405 4253
rect 6349 4179 6405 4188
rect 6670 4122 6722 4128
rect 6722 4082 16665 4110
rect 6670 4064 6722 4070
rect 6670 3918 6722 3924
rect 6722 3878 16665 3906
rect 6670 3860 6722 3866
rect 6670 3714 6722 3720
rect 6722 3674 16665 3702
rect 6670 3656 6722 3662
rect 5727 3548 5783 3557
rect 5463 3496 5519 3505
rect 5727 3483 5783 3492
rect 6349 3548 6405 3557
rect 6349 3483 6405 3492
rect 6941 3496 6993 3502
rect 5463 3431 5519 3440
rect 6941 3438 6993 3444
rect 7553 3496 7605 3502
rect 7553 3438 7605 3444
rect 8165 3496 8217 3502
rect 8165 3438 8217 3444
rect 8777 3496 8829 3502
rect 8777 3438 8829 3444
rect 9389 3496 9441 3502
rect 9389 3438 9441 3444
rect 10001 3496 10053 3502
rect 10001 3438 10053 3444
rect 10613 3496 10665 3502
rect 10613 3438 10665 3444
rect 11225 3496 11277 3502
rect 11225 3438 11277 3444
rect 11837 3496 11889 3502
rect 11837 3438 11889 3444
rect 12449 3496 12501 3502
rect 12449 3438 12501 3444
rect 13061 3496 13113 3502
rect 13061 3438 13113 3444
rect 13673 3496 13725 3502
rect 13673 3438 13725 3444
rect 14285 3496 14337 3502
rect 14285 3438 14337 3444
rect 14897 3496 14949 3502
rect 14897 3438 14949 3444
rect 15509 3496 15561 3502
rect 15509 3438 15561 3444
rect 16121 3496 16173 3502
rect 16121 3438 16173 3444
rect 3739 3125 3795 3134
rect 3739 3060 3795 3069
rect 4555 2700 4611 2709
rect 4555 2635 4611 2644
rect 3739 2173 3795 2182
rect 3739 2108 3795 2117
rect 6953 1977 6981 3438
rect 7565 2079 7593 3438
rect 8177 2181 8205 3438
rect 8789 2283 8817 3438
rect 9401 2385 9429 3438
rect 10013 2487 10041 3438
rect 10001 2481 10053 2487
rect 10001 2423 10053 2429
rect 9389 2379 9441 2385
rect 9389 2321 9441 2327
rect 8777 2277 8829 2283
rect 8777 2219 8829 2225
rect 8165 2175 8217 2181
rect 8165 2117 8217 2123
rect 7553 2073 7605 2079
rect 7553 2015 7605 2021
rect 10447 2073 10499 2079
rect 10447 2015 10499 2021
rect 6941 1971 6993 1977
rect 6941 1913 6993 1919
rect 10139 1971 10191 1977
rect 10139 1913 10191 1919
rect 4555 1748 4611 1757
rect 10151 1754 10179 1913
rect 10459 1754 10487 2015
rect 10625 1977 10653 3438
rect 11063 2277 11115 2283
rect 11063 2219 11115 2225
rect 10755 2175 10807 2181
rect 10755 2117 10807 2123
rect 10613 1971 10665 1977
rect 10613 1913 10665 1919
rect 10767 1754 10795 2117
rect 11075 1754 11103 2219
rect 11237 2079 11265 3438
rect 11679 2481 11731 2487
rect 11679 2423 11731 2429
rect 11371 2379 11423 2385
rect 11371 2321 11423 2327
rect 11225 2073 11277 2079
rect 11225 2015 11277 2021
rect 11383 1754 11411 2321
rect 11691 1754 11719 2423
rect 11849 2181 11877 3438
rect 11837 2175 11889 2181
rect 11837 2117 11889 2123
rect 12295 2073 12347 2079
rect 12295 2015 12347 2021
rect 11987 1971 12039 1977
rect 11987 1913 12039 1919
rect 11999 1754 12027 1913
rect 12307 1754 12335 2015
rect 12461 1977 12489 3438
rect 12603 2175 12655 2181
rect 12603 2117 12655 2123
rect 12449 1971 12501 1977
rect 12449 1913 12501 1919
rect 12615 1754 12643 2117
rect 13073 1977 13101 3438
rect 13685 1977 13713 3438
rect 14143 2073 14195 2079
rect 14143 2015 14195 2021
rect 12911 1971 12963 1977
rect 12911 1913 12963 1919
rect 13061 1971 13113 1977
rect 13061 1913 13113 1919
rect 13219 1971 13271 1977
rect 13219 1913 13271 1919
rect 13527 1971 13579 1977
rect 13527 1913 13579 1919
rect 13673 1971 13725 1977
rect 13673 1913 13725 1919
rect 13835 1971 13887 1977
rect 13835 1913 13887 1919
rect 12923 1754 12951 1913
rect 13231 1754 13259 1913
rect 13539 1754 13567 1913
rect 13847 1754 13875 1913
rect 14155 1754 14183 2015
rect 14297 1977 14325 3438
rect 14759 2175 14811 2181
rect 14759 2117 14811 2123
rect 14285 1971 14337 1977
rect 14285 1913 14337 1919
rect 14451 1971 14503 1977
rect 14451 1913 14503 1919
rect 14463 1754 14491 1913
rect 14771 1754 14799 2117
rect 14909 2079 14937 3438
rect 14897 2073 14949 2079
rect 14897 2015 14949 2021
rect 15521 1977 15549 3438
rect 16133 2181 16161 3438
rect 16121 2175 16173 2181
rect 16121 2117 16173 2123
rect 15509 1971 15561 1977
rect 15509 1913 15561 1919
rect 4555 1683 4611 1692
rect 10139 1748 10191 1754
rect 10139 1690 10191 1696
rect 10447 1748 10499 1754
rect 10447 1690 10499 1696
rect 10755 1748 10807 1754
rect 10755 1690 10807 1696
rect 11063 1748 11115 1754
rect 11063 1690 11115 1696
rect 11371 1748 11423 1754
rect 11371 1690 11423 1696
rect 11679 1748 11731 1754
rect 11679 1690 11731 1696
rect 11987 1748 12039 1754
rect 11987 1690 12039 1696
rect 12295 1748 12347 1754
rect 12295 1690 12347 1696
rect 12603 1748 12655 1754
rect 12603 1690 12655 1696
rect 12911 1748 12963 1754
rect 12911 1690 12963 1696
rect 13219 1748 13271 1754
rect 13219 1690 13271 1696
rect 13527 1748 13579 1754
rect 13527 1690 13579 1696
rect 13835 1748 13887 1754
rect 13835 1690 13887 1696
rect 14143 1748 14195 1754
rect 14143 1690 14195 1696
rect 14451 1748 14503 1754
rect 14451 1690 14503 1696
rect 14759 1748 14811 1754
rect 14759 1690 14811 1696
rect 9969 1480 10025 1489
rect 9969 1415 10025 1424
rect 14877 1480 14933 1489
rect 14877 1415 14933 1424
rect 2540 1378 3480 1406
rect 2488 1360 2540 1366
rect 3739 1136 3795 1145
rect 3739 1071 3795 1080
rect 3109 681 3165 690
rect 3109 616 3165 625
rect 9969 564 10025 573
rect 4555 514 4611 523
rect 9969 499 10025 508
rect 14877 564 14933 573
rect 14877 499 14933 508
rect 4555 449 4611 458
rect 3952 355 4008 364
rect 3952 290 4008 299
rect 4360 355 4416 364
rect 4360 290 4416 299
rect 10128 -11 10137 45
rect 10193 -11 10202 45
rect 10436 -11 10445 45
rect 10501 -11 10510 45
rect 10744 -11 10753 45
rect 10809 -11 10818 45
rect 11052 -11 11061 45
rect 11117 -11 11126 45
rect 11360 -11 11369 45
rect 11425 -11 11434 45
rect 11668 -11 11677 45
rect 11733 -11 11742 45
rect 11976 -11 11985 45
rect 12041 -11 12050 45
rect 12284 -11 12293 45
rect 12349 -11 12358 45
rect 12592 -11 12601 45
rect 12657 -11 12666 45
rect 12900 -11 12909 45
rect 12965 -11 12974 45
rect 13208 -11 13217 45
rect 13273 -11 13282 45
rect 13516 -11 13525 45
rect 13581 -11 13590 45
rect 13824 -11 13833 45
rect 13889 -11 13898 45
rect 14132 -11 14141 45
rect 14197 -11 14206 45
rect 14440 -11 14449 45
rect 14505 -11 14514 45
rect 14748 -11 14757 45
rect 14813 -11 14822 45
<< via2 >>
rect 6925 17378 6981 17380
rect 6925 17326 6927 17378
rect 6927 17326 6979 17378
rect 6979 17326 6981 17378
rect 6925 17324 6981 17326
rect 16541 17378 16597 17380
rect 16541 17326 16543 17378
rect 16543 17326 16595 17378
rect 16595 17326 16597 17378
rect 16541 17324 16597 17326
rect 3695 17167 3751 17169
rect 3695 17115 3697 17167
rect 3697 17115 3749 17167
rect 3749 17115 3751 17167
rect 3695 17113 3751 17115
rect 4091 17167 4147 17169
rect 4091 17115 4093 17167
rect 4093 17115 4145 17167
rect 4145 17115 4147 17167
rect 4091 17113 4147 17115
rect 4701 17167 4757 17169
rect 4701 17115 4703 17167
rect 4703 17115 4755 17167
rect 4755 17115 4757 17167
rect 4701 17113 4757 17115
rect 5949 17167 6005 17169
rect 5949 17115 5951 17167
rect 5951 17115 6003 17167
rect 6003 17115 6005 17167
rect 5949 17113 6005 17115
rect 11842 16635 11898 16691
rect 11842 14899 11898 14955
rect 11842 13163 11898 13219
rect 11842 11427 11898 11483
rect 11842 9691 11898 9747
rect 3695 7995 3751 7997
rect 113 7572 169 7574
rect 113 7520 115 7572
rect 115 7520 167 7572
rect 167 7520 169 7572
rect 113 7518 169 7520
rect 2561 7147 2617 7149
rect 2561 7095 2563 7147
rect 2563 7095 2615 7147
rect 2615 7095 2617 7147
rect 2561 7093 2617 7095
rect 3469 7889 3525 7945
rect 3695 7943 3697 7995
rect 3697 7943 3749 7995
rect 3749 7943 3751 7995
rect 3695 7941 3751 7943
rect 4091 7995 4147 7997
rect 4091 7943 4093 7995
rect 4093 7943 4145 7995
rect 4145 7943 4147 7995
rect 4091 7941 4147 7943
rect 4701 7995 4757 7997
rect 4701 7943 4703 7995
rect 4703 7943 4755 7995
rect 4755 7943 4757 7995
rect 4701 7941 4757 7943
rect 5949 7995 6005 7997
rect 5949 7943 5951 7995
rect 5951 7943 6003 7995
rect 6003 7943 6005 7995
rect 11842 7955 11898 8011
rect 5949 7941 6005 7943
rect 6823 7082 6879 7138
rect 113 6620 169 6622
rect 113 6568 115 6620
rect 115 6568 167 6620
rect 167 6568 169 6620
rect 113 6566 169 6568
rect 2561 6195 2617 6197
rect 2561 6143 2563 6195
rect 2563 6143 2615 6195
rect 2615 6143 2617 6195
rect 2561 6141 2617 6143
rect 113 5583 169 5585
rect 113 5531 115 5583
rect 115 5531 167 5583
rect 167 5531 169 5583
rect 113 5529 169 5531
rect 2561 4961 2617 4963
rect 2561 4909 2563 4961
rect 2563 4909 2615 4961
rect 2615 4909 2617 4961
rect 2561 4907 2617 4909
rect 326 4802 382 4804
rect 326 4750 328 4802
rect 328 4750 380 4802
rect 380 4750 382 4802
rect 326 4748 382 4750
rect 734 4802 790 4804
rect 734 4750 736 4802
rect 736 4750 788 4802
rect 788 4750 790 4802
rect 734 4748 790 4750
rect 1142 4802 1198 4804
rect 1142 4750 1144 4802
rect 1144 4750 1196 4802
rect 1196 4750 1198 4802
rect 1142 4748 1198 4750
rect 1550 4802 1606 4804
rect 1550 4750 1552 4802
rect 1552 4750 1604 4802
rect 1604 4750 1606 4802
rect 1550 4748 1606 4750
rect 1958 4802 2014 4804
rect 1958 4750 1960 4802
rect 1960 4750 2012 4802
rect 2012 4750 2014 4802
rect 1958 4748 2014 4750
rect 2366 4802 2422 4804
rect 2366 4750 2368 4802
rect 2368 4750 2420 4802
rect 2420 4750 2422 4802
rect 2366 4748 2422 4750
rect 509 1430 565 1432
rect 509 1378 511 1430
rect 511 1378 563 1430
rect 563 1378 565 1430
rect 509 1376 565 1378
rect 6819 6480 6875 6482
rect 6819 6428 6821 6480
rect 6821 6428 6873 6480
rect 6873 6428 6875 6480
rect 6819 6426 6875 6428
rect 16611 6480 16667 6482
rect 16611 6428 16613 6480
rect 16613 6428 16665 6480
rect 16665 6428 16667 6480
rect 16611 6426 16667 6428
rect 6819 5564 6875 5566
rect 6819 5512 6821 5564
rect 6821 5512 6873 5564
rect 6873 5512 6875 5564
rect 6819 5510 6875 5512
rect 16611 5564 16667 5566
rect 16611 5512 16613 5564
rect 16613 5512 16665 5564
rect 16665 5512 16667 5564
rect 16611 5510 16667 5512
rect 11774 5008 11830 5064
rect 5727 4242 5783 4244
rect 5727 4190 5729 4242
rect 5729 4190 5781 4242
rect 5781 4190 5783 4242
rect 5727 4188 5783 4190
rect 6349 4242 6405 4244
rect 6349 4190 6351 4242
rect 6351 4190 6403 4242
rect 6403 4190 6405 4242
rect 6349 4188 6405 4190
rect 5727 3546 5783 3548
rect 5463 3440 5519 3496
rect 5727 3494 5729 3546
rect 5729 3494 5781 3546
rect 5781 3494 5783 3546
rect 5727 3492 5783 3494
rect 6349 3546 6405 3548
rect 6349 3494 6351 3546
rect 6351 3494 6403 3546
rect 6403 3494 6405 3546
rect 6349 3492 6405 3494
rect 3739 3123 3795 3125
rect 3739 3071 3741 3123
rect 3741 3071 3793 3123
rect 3793 3071 3795 3123
rect 3739 3069 3795 3071
rect 4555 2698 4611 2700
rect 4555 2646 4557 2698
rect 4557 2646 4609 2698
rect 4609 2646 4611 2698
rect 4555 2644 4611 2646
rect 3739 2171 3795 2173
rect 3739 2119 3741 2171
rect 3741 2119 3793 2171
rect 3793 2119 3795 2171
rect 3739 2117 3795 2119
rect 4555 1746 4611 1748
rect 4555 1694 4557 1746
rect 4557 1694 4609 1746
rect 4609 1694 4611 1746
rect 4555 1692 4611 1694
rect 9969 1478 10025 1480
rect 9969 1426 9971 1478
rect 9971 1426 10023 1478
rect 10023 1426 10025 1478
rect 9969 1424 10025 1426
rect 14877 1478 14933 1480
rect 14877 1426 14879 1478
rect 14879 1426 14931 1478
rect 14931 1426 14933 1478
rect 14877 1424 14933 1426
rect 3739 1134 3795 1136
rect 3739 1082 3741 1134
rect 3741 1082 3793 1134
rect 3793 1082 3795 1134
rect 3739 1080 3795 1082
rect 3109 679 3165 681
rect 3109 627 3111 679
rect 3111 627 3163 679
rect 3163 627 3165 679
rect 3109 625 3165 627
rect 9969 562 10025 564
rect 4555 512 4611 514
rect 4555 460 4557 512
rect 4557 460 4609 512
rect 4609 460 4611 512
rect 9969 510 9971 562
rect 9971 510 10023 562
rect 10023 510 10025 562
rect 9969 508 10025 510
rect 14877 562 14933 564
rect 14877 510 14879 562
rect 14879 510 14931 562
rect 14931 510 14933 562
rect 14877 508 14933 510
rect 4555 458 4611 460
rect 3952 353 4008 355
rect 3952 301 3954 353
rect 3954 301 4006 353
rect 4006 301 4008 353
rect 3952 299 4008 301
rect 4360 353 4416 355
rect 4360 301 4362 353
rect 4362 301 4414 353
rect 4414 301 4416 353
rect 4360 299 4416 301
rect 10137 43 10193 45
rect 10137 -9 10139 43
rect 10139 -9 10191 43
rect 10191 -9 10193 43
rect 10137 -11 10193 -9
rect 10445 43 10501 45
rect 10445 -9 10447 43
rect 10447 -9 10499 43
rect 10499 -9 10501 43
rect 10445 -11 10501 -9
rect 10753 43 10809 45
rect 10753 -9 10755 43
rect 10755 -9 10807 43
rect 10807 -9 10809 43
rect 10753 -11 10809 -9
rect 11061 43 11117 45
rect 11061 -9 11063 43
rect 11063 -9 11115 43
rect 11115 -9 11117 43
rect 11061 -11 11117 -9
rect 11369 43 11425 45
rect 11369 -9 11371 43
rect 11371 -9 11423 43
rect 11423 -9 11425 43
rect 11369 -11 11425 -9
rect 11677 43 11733 45
rect 11677 -9 11679 43
rect 11679 -9 11731 43
rect 11731 -9 11733 43
rect 11677 -11 11733 -9
rect 11985 43 12041 45
rect 11985 -9 11987 43
rect 11987 -9 12039 43
rect 12039 -9 12041 43
rect 11985 -11 12041 -9
rect 12293 43 12349 45
rect 12293 -9 12295 43
rect 12295 -9 12347 43
rect 12347 -9 12349 43
rect 12293 -11 12349 -9
rect 12601 43 12657 45
rect 12601 -9 12603 43
rect 12603 -9 12655 43
rect 12655 -9 12657 43
rect 12601 -11 12657 -9
rect 12909 43 12965 45
rect 12909 -9 12911 43
rect 12911 -9 12963 43
rect 12963 -9 12965 43
rect 12909 -11 12965 -9
rect 13217 43 13273 45
rect 13217 -9 13219 43
rect 13219 -9 13271 43
rect 13271 -9 13273 43
rect 13217 -11 13273 -9
rect 13525 43 13581 45
rect 13525 -9 13527 43
rect 13527 -9 13579 43
rect 13579 -9 13581 43
rect 13525 -11 13581 -9
rect 13833 43 13889 45
rect 13833 -9 13835 43
rect 13835 -9 13887 43
rect 13887 -9 13889 43
rect 13833 -11 13889 -9
rect 14141 43 14197 45
rect 14141 -9 14143 43
rect 14143 -9 14195 43
rect 14195 -9 14197 43
rect 14141 -11 14197 -9
rect 14449 43 14505 45
rect 14449 -9 14451 43
rect 14451 -9 14503 43
rect 14503 -9 14505 43
rect 14449 -11 14505 -9
rect 14757 43 14813 45
rect 14757 -9 14759 43
rect 14759 -9 14811 43
rect 14811 -9 14813 43
rect 14757 -11 14813 -9
<< metal3 >>
rect -1496 18902 18362 18908
rect -1496 18838 -1490 18902
rect -1426 18838 -1354 18902
rect -1290 18838 -1218 18902
rect -1154 18838 18020 18902
rect 18084 18838 18156 18902
rect 18220 18838 18292 18902
rect 18356 18838 18362 18902
rect -1496 18766 18362 18838
rect -1496 18702 -1490 18766
rect -1426 18702 -1354 18766
rect -1290 18702 -1218 18766
rect -1154 18702 18020 18766
rect 18084 18702 18156 18766
rect 18220 18702 18292 18766
rect 18356 18702 18362 18766
rect -1496 18630 18362 18702
rect -1496 18566 -1490 18630
rect -1426 18566 -1354 18630
rect -1290 18566 -1218 18630
rect -1154 18566 3840 18630
rect 3904 18566 5945 18630
rect 6009 18566 10325 18630
rect 10389 18566 14172 18630
rect 14236 18566 18020 18630
rect 18084 18566 18156 18630
rect 18220 18566 18292 18630
rect 18356 18566 18362 18630
rect -1496 18560 18362 18566
rect -800 18206 17666 18212
rect -800 18142 -794 18206
rect -730 18142 -658 18206
rect -594 18142 -522 18206
rect -458 18142 17324 18206
rect 17388 18142 17460 18206
rect 17524 18142 17596 18206
rect 17660 18142 17666 18206
rect -800 18070 17666 18142
rect -800 18006 -794 18070
rect -730 18006 -658 18070
rect -594 18006 -522 18070
rect -458 18006 17324 18070
rect 17388 18006 17460 18070
rect 17524 18006 17596 18070
rect 17660 18006 17666 18070
rect -800 17934 17666 18006
rect -800 17870 -794 17934
rect -730 17870 -658 17934
rect -594 17870 -522 17934
rect -458 17870 2449 17934
rect 2513 17870 3691 17934
rect 3755 17870 5796 17934
rect 5860 17870 6921 17934
rect 6985 17870 10186 17934
rect 10250 17870 11838 17934
rect 11902 17870 13755 17934
rect 13819 17870 16537 17934
rect 16601 17870 17324 17934
rect 17388 17870 17460 17934
rect 17524 17870 17596 17934
rect 17660 17870 17666 17934
rect -800 17864 17666 17870
rect 6904 17390 7002 17401
rect 16520 17390 16618 17401
rect 6904 17384 10256 17390
rect 3685 17252 4767 17328
rect 6904 17320 6921 17384
rect 6985 17320 10186 17384
rect 10250 17320 10256 17384
rect 6904 17314 10256 17320
rect 16520 17384 17394 17390
rect 16520 17320 16537 17384
rect 16601 17320 17324 17384
rect 17388 17320 17394 17384
rect 16520 17314 17394 17320
rect 6904 17303 7002 17314
rect 16520 17303 16618 17314
rect 3685 17190 3761 17252
rect 4691 17190 4767 17252
rect -40 17176 266 17182
rect -40 17112 -25 17176
rect 39 17112 196 17176
rect 260 17112 266 17176
rect -40 17106 266 17112
rect 2434 17176 2665 17182
rect 2434 17112 2449 17176
rect 2513 17112 2595 17176
rect 2659 17112 2665 17176
rect 2434 17106 2665 17112
rect 3674 17173 3772 17190
rect 4070 17179 4168 17190
rect 4680 17179 4778 17190
rect 5928 17179 6026 17190
rect 3674 17109 3691 17173
rect 3755 17109 3772 17173
rect 3674 17092 3772 17109
rect 3834 17173 4618 17179
rect 3834 17109 3840 17173
rect 3904 17169 4618 17173
rect 3904 17113 4091 17169
rect 4147 17113 4618 17169
rect 3904 17109 4618 17113
rect 3834 17103 4618 17109
rect 4070 17092 4168 17103
rect 4081 17030 4157 17092
rect -1224 17024 4157 17030
rect -1224 16960 -1218 17024
rect -1154 16960 4157 17024
rect -1224 16954 4157 16960
rect 4542 17030 4618 17103
rect 4680 17173 5866 17179
rect 4680 17169 5796 17173
rect 4680 17113 4701 17169
rect 4757 17113 5796 17169
rect 4680 17109 5796 17113
rect 5860 17109 5866 17173
rect 4680 17103 5866 17109
rect 5928 17173 14242 17179
rect 5928 17109 5945 17173
rect 6009 17109 10325 17173
rect 10389 17109 14172 17173
rect 14236 17109 14242 17173
rect 5928 17103 14242 17109
rect 4680 17092 4778 17103
rect 5928 17092 6026 17103
rect 5939 17030 6015 17092
rect 4542 16954 6015 17030
rect 11821 16701 11919 16712
rect 11821 16695 13825 16701
rect -40 16664 266 16670
rect -40 16600 -34 16664
rect 30 16600 196 16664
rect 260 16600 266 16664
rect -40 16594 266 16600
rect 2434 16664 2665 16670
rect 2434 16600 2440 16664
rect 2504 16600 2595 16664
rect 2659 16600 2665 16664
rect 11821 16631 11838 16695
rect 11902 16631 13755 16695
rect 13819 16631 13825 16695
rect 11821 16625 13825 16631
rect 11821 16614 11919 16625
rect 2434 16594 2665 16600
rect 11821 14959 11919 14976
rect -528 14928 45 14934
rect -528 14864 -522 14928
rect -458 14864 45 14928
rect -528 14858 45 14864
rect 2434 14928 2665 14934
rect 2434 14864 2440 14928
rect 2504 14864 2595 14928
rect 2659 14864 2665 14928
rect 11821 14895 11838 14959
rect 11902 14895 11919 14959
rect 11821 14878 11919 14895
rect 2434 14858 2665 14864
rect 11821 13223 11919 13240
rect -528 13192 45 13198
rect -528 13128 -522 13192
rect -458 13128 -34 13192
rect 30 13128 45 13192
rect 2434 13128 2440 13192
rect 2504 13190 2510 13192
rect 2504 13130 2519 13190
rect 11821 13159 11838 13223
rect 11902 13159 11919 13223
rect 11821 13142 11919 13159
rect 2504 13128 2510 13130
rect -528 13122 45 13128
rect 11821 11487 11919 11504
rect -528 11456 45 11462
rect -528 11392 -522 11456
rect -458 11392 -34 11456
rect 30 11392 45 11456
rect 2434 11392 2440 11456
rect 2504 11454 2510 11456
rect 2504 11394 2519 11454
rect 11821 11423 11838 11487
rect 11902 11423 11919 11487
rect 11821 11406 11919 11423
rect 2504 11392 2510 11394
rect -528 11386 45 11392
rect 11821 9751 11919 9768
rect -528 9720 45 9726
rect -528 9656 -522 9720
rect -458 9656 -34 9720
rect 30 9656 45 9720
rect 2434 9656 2440 9720
rect 2504 9718 2510 9720
rect 2504 9658 2519 9718
rect 11821 9687 11838 9751
rect 11902 9687 11919 9751
rect 11821 9670 11919 9687
rect 2504 9656 2510 9658
rect -528 9650 45 9656
rect 3310 8080 4767 8156
rect 3310 7990 3386 8080
rect 3685 8018 3761 8080
rect 4691 8018 4767 8080
rect -528 7984 45 7990
rect 2443 7984 3386 7990
rect -528 7920 -522 7984
rect -458 7920 -34 7984
rect 30 7920 45 7984
rect 2230 7920 2236 7984
rect 2300 7920 2306 7984
rect 2434 7920 2440 7984
rect 2504 7920 3386 7984
rect 3674 7997 3772 8018
rect 4070 8007 4168 8018
rect -528 7914 45 7920
rect 2443 7914 3386 7920
rect 3448 7945 3546 7966
rect 3448 7889 3469 7945
rect 3525 7889 3546 7945
rect 3674 7941 3695 7997
rect 3751 7941 3772 7997
rect 3674 7920 3772 7941
rect 3834 7997 4168 8007
rect 3834 7941 4091 7997
rect 4147 7941 4168 7997
rect 3834 7931 4168 7941
rect 3448 7868 3546 7889
rect 3459 7806 3535 7868
rect 3834 7806 3910 7931
rect 4070 7920 4168 7931
rect 4680 7997 4778 8018
rect 5928 8007 6026 8018
rect 4680 7941 4701 7997
rect 4757 7941 4778 7997
rect 4680 7920 4778 7941
rect 4840 8001 6026 8007
rect 4840 7937 5945 8001
rect 6009 7937 6026 8001
rect 4840 7931 6026 7937
rect 11821 8015 11919 8032
rect 11821 7951 11838 8015
rect 11902 7951 11919 8015
rect 11821 7934 11919 7951
rect 3459 7730 3910 7806
rect 4081 7858 4157 7920
rect 4840 7858 4916 7931
rect 5928 7920 6026 7931
rect 4081 7782 4916 7858
rect 92 7584 190 7595
rect -1224 7578 190 7584
rect -1224 7514 -1218 7578
rect -1154 7514 109 7578
rect 173 7514 190 7578
rect -1224 7508 190 7514
rect 92 7497 190 7508
rect 2540 7159 2638 7170
rect 2230 7153 2776 7159
rect 2230 7089 2236 7153
rect 2300 7089 2408 7153
rect 2472 7149 2706 7153
rect 2472 7093 2561 7149
rect 2617 7093 2706 7149
rect 2472 7089 2706 7093
rect 2770 7089 2776 7153
rect 6802 7148 6900 7159
rect 2230 7083 2776 7089
rect 5939 7142 6900 7148
rect 2540 7072 2638 7083
rect 5939 7078 5945 7142
rect 6009 7078 6819 7142
rect 6883 7078 6900 7142
rect 5939 7072 6900 7078
rect 6802 7061 6900 7072
rect 92 6632 190 6643
rect -1224 6626 190 6632
rect -1224 6562 -1218 6626
rect -1154 6562 109 6626
rect 173 6562 190 6626
rect -1224 6556 190 6562
rect 92 6545 190 6556
rect 6798 6492 6896 6503
rect 6339 6486 6896 6492
rect 6339 6422 6345 6486
rect 6409 6422 6815 6486
rect 6879 6422 6896 6486
rect 6339 6416 6896 6422
rect 6798 6405 6896 6416
rect 16590 6492 16688 6503
rect 16590 6486 18090 6492
rect 16590 6482 18020 6486
rect 16590 6426 16611 6482
rect 16667 6426 18020 6482
rect 16590 6422 18020 6426
rect 18084 6422 18090 6486
rect 16590 6416 18090 6422
rect 16590 6405 16688 6416
rect 2540 6207 2638 6218
rect 2540 6201 2776 6207
rect 2540 6137 2557 6201
rect 2621 6137 2706 6201
rect 2770 6137 2776 6201
rect 2540 6131 2776 6137
rect 2540 6120 2638 6131
rect 92 5595 190 5606
rect -1224 5589 190 5595
rect -1224 5525 -1218 5589
rect -1154 5525 109 5589
rect 173 5525 190 5589
rect 6798 5576 6896 5587
rect -1224 5519 190 5525
rect 92 5508 190 5519
rect 5717 5570 6896 5576
rect 5717 5506 5723 5570
rect 5787 5566 6896 5570
rect 5787 5510 6819 5566
rect 6875 5510 6896 5566
rect 5787 5506 6896 5510
rect 5717 5500 6896 5506
rect 6798 5489 6896 5500
rect 16590 5576 16688 5587
rect 16590 5570 17394 5576
rect 16590 5566 17324 5570
rect 16590 5510 16611 5566
rect 16667 5510 17324 5566
rect 16590 5506 17324 5510
rect 17388 5506 17394 5570
rect 16590 5500 17394 5506
rect 16590 5489 16688 5500
rect -1496 5233 1765 5239
rect -1496 5169 1695 5233
rect 1759 5169 1765 5233
rect -1496 5163 1765 5169
rect -1496 5095 949 5101
rect -1496 5031 879 5095
rect 943 5031 949 5095
rect -1496 5025 949 5031
rect 11753 5068 11851 5085
rect 11753 5004 11770 5068
rect 11834 5004 11851 5068
rect 11753 4987 11851 5004
rect 2540 4973 2638 4984
rect 1878 4967 3662 4973
rect -1496 4887 541 4963
rect 1878 4903 1884 4967
rect 1948 4903 2557 4967
rect 2621 4903 3592 4967
rect 3656 4903 3662 4967
rect 1878 4897 3662 4903
rect 305 4814 403 4825
rect -1496 4804 403 4814
rect -1496 4748 326 4804
rect 382 4748 403 4804
rect -1496 4738 403 4748
rect 465 4814 541 4887
rect 2540 4886 2638 4897
rect 713 4814 811 4825
rect 1121 4814 1219 4825
rect 1529 4814 1627 4825
rect 1937 4814 2035 4825
rect 2345 4814 2443 4825
rect 465 4804 811 4814
rect 465 4748 734 4804
rect 790 4748 811 4804
rect 465 4738 811 4748
rect 873 4808 1219 4814
rect 873 4744 879 4808
rect 943 4804 1219 4808
rect 943 4748 1142 4804
rect 1198 4748 1219 4804
rect 943 4744 1219 4748
rect 873 4738 1219 4744
rect 1281 4808 1627 4814
rect 1281 4744 1287 4808
rect 1351 4804 1627 4808
rect 1351 4748 1550 4804
rect 1606 4748 1627 4804
rect 1351 4744 1627 4748
rect 1281 4738 1627 4744
rect 1689 4808 2035 4814
rect 1689 4744 1695 4808
rect 1759 4804 2035 4808
rect 1759 4748 1958 4804
rect 2014 4748 2035 4804
rect 1759 4744 2035 4748
rect 1689 4738 2035 4744
rect 2097 4808 2443 4814
rect 2097 4744 2103 4808
rect 2167 4804 2443 4808
rect 2167 4748 2366 4804
rect 2422 4748 2443 4804
rect 2167 4744 2443 4748
rect 2097 4738 2443 4744
rect 305 4727 403 4738
rect 713 4727 811 4738
rect 1121 4727 1219 4738
rect 1529 4727 1627 4738
rect 1937 4727 2035 4738
rect 2345 4727 2443 4738
rect 1867 4658 1965 4669
rect -528 4652 1965 4658
rect -528 4588 -522 4652
rect -458 4588 1884 4652
rect 1948 4588 1965 4652
rect -528 4582 1965 4588
rect 1867 4571 1965 4582
rect -1496 4514 1357 4520
rect -1496 4450 1287 4514
rect 1351 4450 1357 4514
rect -1496 4444 1357 4450
rect -1496 4376 2173 4382
rect -1496 4312 2103 4376
rect 2167 4312 2173 4376
rect -1496 4306 2173 4312
rect 3586 4251 3892 4257
rect 3586 4187 3592 4251
rect 3656 4187 3822 4251
rect 3886 4187 3892 4251
rect 3586 4181 3892 4187
rect 4224 4251 4504 4257
rect 4224 4187 4230 4251
rect 4294 4187 4434 4251
rect 4498 4249 4504 4251
rect 4498 4189 4513 4249
rect 5706 4248 5804 4265
rect 4498 4187 4504 4189
rect 4224 4181 4504 4187
rect 5706 4184 5723 4248
rect 5787 4184 5804 4248
rect 5706 4167 5804 4184
rect 6328 4248 6426 4265
rect 6328 4184 6345 4248
rect 6409 4184 6426 4248
rect 6328 4167 6426 4184
rect 5453 3631 6415 3707
rect 4224 3535 4513 3541
rect 3586 3471 3592 3535
rect 3656 3471 3662 3535
rect 3816 3471 3822 3535
rect 3886 3471 3892 3535
rect 4224 3471 4230 3535
rect 4294 3471 4443 3535
rect 4507 3471 4513 3535
rect 5453 3517 5529 3631
rect 6339 3569 6415 3631
rect 5706 3552 5804 3569
rect 5442 3506 5540 3517
rect 4224 3465 4513 3471
rect 4437 3357 4513 3465
rect 4583 3500 5540 3506
rect 4583 3436 4589 3500
rect 4653 3496 5540 3500
rect 4653 3440 5463 3496
rect 5519 3440 5540 3496
rect 5706 3488 5723 3552
rect 5787 3488 5804 3552
rect 5706 3471 5804 3488
rect 6328 3552 6426 3569
rect 6328 3488 6345 3552
rect 6409 3488 6426 3552
rect 6328 3471 6426 3488
rect 4653 3436 5540 3440
rect 4583 3430 5540 3436
rect 5442 3419 5540 3430
rect 5717 3357 5793 3471
rect 4437 3281 5793 3357
rect 3718 3135 3816 3146
rect 3718 3129 4659 3135
rect 3718 3065 3735 3129
rect 3799 3065 4589 3129
rect 4653 3065 4659 3129
rect 3718 3059 4659 3065
rect 3718 3048 3816 3059
rect 4534 2710 4632 2721
rect 4224 2704 4632 2710
rect 4224 2640 4230 2704
rect 4294 2640 4551 2704
rect 4615 2640 4632 2704
rect 4224 2634 4632 2640
rect 4534 2623 4632 2634
rect 1683 2539 1781 2550
rect -1224 2533 1781 2539
rect -1224 2469 -1218 2533
rect -1154 2469 1700 2533
rect 1764 2469 1781 2533
rect -1224 2463 1781 2469
rect 1683 2452 1781 2463
rect 3718 2183 3816 2194
rect 1694 2177 3816 2183
rect 1694 2113 1700 2177
rect 1764 2113 3735 2177
rect 3799 2113 3816 2177
rect 1694 2107 3816 2113
rect 3718 2096 3816 2107
rect 4534 1752 4632 1769
rect 4534 1688 4551 1752
rect 4615 1688 4632 1752
rect 4534 1671 4632 1688
rect 9948 1490 10046 1501
rect 14856 1490 14954 1501
rect 6610 1484 13825 1490
rect 488 1442 586 1453
rect -1496 1432 586 1442
rect -1496 1376 509 1432
rect 565 1376 586 1432
rect 6610 1420 6616 1484
rect 6680 1480 10186 1484
rect 6680 1424 9969 1480
rect 10025 1424 10186 1480
rect 6680 1420 10186 1424
rect 10250 1420 13755 1484
rect 13819 1420 13825 1484
rect 6610 1414 13825 1420
rect 14718 1484 17394 1490
rect 14718 1420 14724 1484
rect 14788 1480 17324 1484
rect 14788 1424 14877 1480
rect 14933 1424 17324 1480
rect 14788 1420 17324 1424
rect 17388 1420 17394 1484
rect 14718 1414 17394 1420
rect 9948 1403 10046 1414
rect 14856 1403 14954 1414
rect -1496 1366 586 1376
rect 488 1355 586 1366
rect 3718 1146 3816 1157
rect 2624 1140 6547 1146
rect 2624 1076 2630 1140
rect 2694 1076 3735 1140
rect 3799 1076 6477 1140
rect 6541 1076 6547 1140
rect 2624 1070 6547 1076
rect 3718 1059 3816 1070
rect 3088 685 3186 702
rect 3088 621 3105 685
rect 3169 621 3186 685
rect 3088 604 3186 621
rect 9948 574 10046 585
rect 14856 574 14954 585
rect 9948 568 14242 574
rect 4534 524 4632 535
rect 3041 518 6686 524
rect 3041 454 3047 518
rect 3111 454 4551 518
rect 4615 454 6616 518
rect 6680 454 6686 518
rect 9948 504 9965 568
rect 10029 504 10325 568
rect 10389 504 14172 568
rect 14236 504 14242 568
rect 9948 498 14242 504
rect 14856 568 18090 574
rect 14856 504 14873 568
rect 14937 504 18020 568
rect 18084 504 18090 568
rect 14856 498 18090 504
rect 9948 487 10046 498
rect 14856 487 14954 498
rect 3041 448 6686 454
rect 4534 437 4632 448
rect 1683 415 1781 432
rect 1683 351 1700 415
rect 1764 351 1781 415
rect 1683 334 1781 351
rect 3931 359 4029 376
rect 3931 295 3948 359
rect 4012 295 4029 359
rect 3931 278 4029 295
rect 4339 359 4437 376
rect 4339 295 4356 359
rect 4420 295 4437 359
rect 4339 278 4437 295
rect 10116 55 10214 66
rect 9821 49 10214 55
rect 9821 -15 9827 49
rect 9891 45 10214 49
rect 9891 -11 10137 45
rect 10193 -11 10214 45
rect 9891 -15 10214 -11
rect 9821 -21 10214 -15
rect 10116 -32 10214 -21
rect 10424 45 10522 66
rect 10424 -11 10445 45
rect 10501 -11 10522 45
rect 10424 -32 10522 -11
rect 10732 49 10830 66
rect 10732 -15 10749 49
rect 10813 -15 10830 49
rect 10732 -32 10830 -15
rect 11040 49 11138 66
rect 11040 -15 11057 49
rect 11121 -15 11138 49
rect 11040 -32 11138 -15
rect 11348 49 11446 66
rect 11348 -15 11365 49
rect 11429 -15 11446 49
rect 11348 -32 11446 -15
rect 11656 49 11754 66
rect 11656 -15 11673 49
rect 11737 -15 11754 49
rect 11656 -32 11754 -15
rect 11964 49 12062 66
rect 11964 -15 11981 49
rect 12045 -15 12062 49
rect 11964 -32 12062 -15
rect 12272 49 12370 66
rect 12272 -15 12289 49
rect 12353 -15 12370 49
rect 12272 -32 12370 -15
rect 12580 49 12678 66
rect 12580 -15 12597 49
rect 12661 -15 12678 49
rect 12580 -32 12678 -15
rect 12888 49 12986 66
rect 12888 -15 12905 49
rect 12969 -15 12986 49
rect 12888 -32 12986 -15
rect 13196 49 13294 66
rect 13196 -15 13213 49
rect 13277 -15 13294 49
rect 13196 -32 13294 -15
rect 13504 49 13602 66
rect 13504 -15 13521 49
rect 13585 -15 13602 49
rect 13504 -32 13602 -15
rect 13812 55 13910 66
rect 14120 55 14218 66
rect 13812 49 14048 55
rect 13812 45 13978 49
rect 13812 -11 13833 45
rect 13889 -11 13978 45
rect 13812 -15 13978 -11
rect 14042 -15 14048 49
rect 13812 -21 14048 -15
rect 14120 45 14366 55
rect 14120 -11 14141 45
rect 14197 -11 14366 45
rect 14120 -21 14366 -11
rect 13812 -32 13910 -21
rect 14120 -32 14218 -21
rect 10435 -94 10511 -32
rect 14290 -94 14366 -21
rect 14428 49 14526 66
rect 14736 55 14834 66
rect 14428 -15 14445 49
rect 14509 -15 14526 49
rect 14428 -32 14526 -15
rect 14588 45 14834 55
rect 14588 -11 14757 45
rect 14813 -11 14834 45
rect 14588 -21 14834 -11
rect 14588 -94 14664 -21
rect 14736 -32 14834 -21
rect 10435 -100 10533 -94
rect 10435 -164 10463 -100
rect 10527 -164 10533 -100
rect 10435 -170 10533 -164
rect 14290 -100 14380 -94
rect 14290 -164 14310 -100
rect 14374 -164 14380 -100
rect 14290 -170 14380 -164
rect 14580 -100 14664 -94
rect 14580 -164 14586 -100
rect 14650 -164 14664 -100
rect 14580 -170 14664 -164
rect -800 -458 17666 -452
rect -800 -522 -794 -458
rect -730 -522 -658 -458
rect -594 -522 -522 -458
rect -458 -522 1700 -458
rect 1764 -522 3047 -458
rect 3111 -522 6616 -458
rect 6680 -522 10186 -458
rect 10250 -522 13755 -458
rect 13819 -522 14724 -458
rect 14788 -522 17324 -458
rect 17388 -522 17460 -458
rect 17524 -522 17596 -458
rect 17660 -522 17666 -458
rect -800 -594 17666 -522
rect -800 -658 -794 -594
rect -730 -658 -658 -594
rect -594 -658 -522 -594
rect -458 -658 17324 -594
rect 17388 -658 17460 -594
rect 17524 -658 17596 -594
rect 17660 -658 17666 -594
rect -800 -730 17666 -658
rect -800 -794 -794 -730
rect -730 -794 -658 -730
rect -594 -794 -522 -730
rect -458 -794 17324 -730
rect 17388 -794 17460 -730
rect 17524 -794 17596 -730
rect 17660 -794 17666 -730
rect -800 -800 17666 -794
rect -1496 -1154 18362 -1148
rect -1496 -1218 -1490 -1154
rect -1426 -1218 -1354 -1154
rect -1290 -1218 -1218 -1154
rect -1154 -1218 2630 -1154
rect 2694 -1218 6477 -1154
rect 6541 -1218 9965 -1154
rect 10029 -1218 10325 -1154
rect 10389 -1218 14172 -1154
rect 14236 -1218 14873 -1154
rect 14937 -1218 18020 -1154
rect 18084 -1218 18156 -1154
rect 18220 -1218 18292 -1154
rect 18356 -1218 18362 -1154
rect -1496 -1290 18362 -1218
rect -1496 -1354 -1490 -1290
rect -1426 -1354 -1354 -1290
rect -1290 -1354 -1218 -1290
rect -1154 -1354 18020 -1290
rect 18084 -1354 18156 -1290
rect 18220 -1354 18292 -1290
rect 18356 -1354 18362 -1290
rect -1496 -1426 18362 -1354
rect -1496 -1490 -1490 -1426
rect -1426 -1490 -1354 -1426
rect -1290 -1490 -1218 -1426
rect -1154 -1490 18020 -1426
rect 18084 -1490 18156 -1426
rect 18220 -1490 18292 -1426
rect 18356 -1490 18362 -1426
rect -1496 -1496 18362 -1490
<< via3 >>
rect -1490 18838 -1426 18902
rect -1354 18838 -1290 18902
rect -1218 18838 -1154 18902
rect 18020 18838 18084 18902
rect 18156 18838 18220 18902
rect 18292 18838 18356 18902
rect -1490 18702 -1426 18766
rect -1354 18702 -1290 18766
rect -1218 18702 -1154 18766
rect 18020 18702 18084 18766
rect 18156 18702 18220 18766
rect 18292 18702 18356 18766
rect -1490 18566 -1426 18630
rect -1354 18566 -1290 18630
rect -1218 18566 -1154 18630
rect 3840 18566 3904 18630
rect 5945 18566 6009 18630
rect 10325 18566 10389 18630
rect 14172 18566 14236 18630
rect 18020 18566 18084 18630
rect 18156 18566 18220 18630
rect 18292 18566 18356 18630
rect -794 18142 -730 18206
rect -658 18142 -594 18206
rect -522 18142 -458 18206
rect 17324 18142 17388 18206
rect 17460 18142 17524 18206
rect 17596 18142 17660 18206
rect -794 18006 -730 18070
rect -658 18006 -594 18070
rect -522 18006 -458 18070
rect 17324 18006 17388 18070
rect 17460 18006 17524 18070
rect 17596 18006 17660 18070
rect -794 17870 -730 17934
rect -658 17870 -594 17934
rect -522 17870 -458 17934
rect 2449 17870 2513 17934
rect 3691 17870 3755 17934
rect 5796 17870 5860 17934
rect 6921 17870 6985 17934
rect 10186 17870 10250 17934
rect 11838 17870 11902 17934
rect 13755 17870 13819 17934
rect 16537 17870 16601 17934
rect 17324 17870 17388 17934
rect 17460 17870 17524 17934
rect 17596 17870 17660 17934
rect 6921 17380 6985 17384
rect 6921 17324 6925 17380
rect 6925 17324 6981 17380
rect 6981 17324 6985 17380
rect 6921 17320 6985 17324
rect 10186 17320 10250 17384
rect 16537 17380 16601 17384
rect 16537 17324 16541 17380
rect 16541 17324 16597 17380
rect 16597 17324 16601 17380
rect 16537 17320 16601 17324
rect 17324 17320 17388 17384
rect -25 17112 39 17176
rect 196 17112 260 17176
rect 2449 17112 2513 17176
rect 2595 17112 2659 17176
rect 3691 17169 3755 17173
rect 3691 17113 3695 17169
rect 3695 17113 3751 17169
rect 3751 17113 3755 17169
rect 3691 17109 3755 17113
rect 3840 17109 3904 17173
rect -1218 16960 -1154 17024
rect 5796 17109 5860 17173
rect 5945 17169 6009 17173
rect 5945 17113 5949 17169
rect 5949 17113 6005 17169
rect 6005 17113 6009 17169
rect 5945 17109 6009 17113
rect 10325 17109 10389 17173
rect 14172 17109 14236 17173
rect -34 16600 30 16664
rect 196 16600 260 16664
rect 2440 16600 2504 16664
rect 2595 16600 2659 16664
rect 11838 16691 11902 16695
rect 11838 16635 11842 16691
rect 11842 16635 11898 16691
rect 11898 16635 11902 16691
rect 11838 16631 11902 16635
rect 13755 16631 13819 16695
rect -522 14864 -458 14928
rect 2440 14864 2504 14928
rect 2595 14864 2659 14928
rect 11838 14955 11902 14959
rect 11838 14899 11842 14955
rect 11842 14899 11898 14955
rect 11898 14899 11902 14955
rect 11838 14895 11902 14899
rect -522 13128 -458 13192
rect -34 13128 30 13192
rect 2440 13128 2504 13192
rect 11838 13219 11902 13223
rect 11838 13163 11842 13219
rect 11842 13163 11898 13219
rect 11898 13163 11902 13219
rect 11838 13159 11902 13163
rect -522 11392 -458 11456
rect -34 11392 30 11456
rect 2440 11392 2504 11456
rect 11838 11483 11902 11487
rect 11838 11427 11842 11483
rect 11842 11427 11898 11483
rect 11898 11427 11902 11483
rect 11838 11423 11902 11427
rect -522 9656 -458 9720
rect -34 9656 30 9720
rect 2440 9656 2504 9720
rect 11838 9747 11902 9751
rect 11838 9691 11842 9747
rect 11842 9691 11898 9747
rect 11898 9691 11902 9747
rect 11838 9687 11902 9691
rect -522 7920 -458 7984
rect -34 7920 30 7984
rect 2236 7920 2300 7984
rect 2440 7920 2504 7984
rect 5945 7997 6009 8001
rect 5945 7941 5949 7997
rect 5949 7941 6005 7997
rect 6005 7941 6009 7997
rect 5945 7937 6009 7941
rect 11838 8011 11902 8015
rect 11838 7955 11842 8011
rect 11842 7955 11898 8011
rect 11898 7955 11902 8011
rect 11838 7951 11902 7955
rect -1218 7514 -1154 7578
rect 109 7574 173 7578
rect 109 7518 113 7574
rect 113 7518 169 7574
rect 169 7518 173 7574
rect 109 7514 173 7518
rect 2236 7089 2300 7153
rect 2408 7089 2472 7153
rect 2706 7089 2770 7153
rect 5945 7078 6009 7142
rect 6819 7138 6883 7142
rect 6819 7082 6823 7138
rect 6823 7082 6879 7138
rect 6879 7082 6883 7138
rect 6819 7078 6883 7082
rect -1218 6562 -1154 6626
rect 109 6622 173 6626
rect 109 6566 113 6622
rect 113 6566 169 6622
rect 169 6566 173 6622
rect 109 6562 173 6566
rect 6345 6422 6409 6486
rect 6815 6482 6879 6486
rect 6815 6426 6819 6482
rect 6819 6426 6875 6482
rect 6875 6426 6879 6482
rect 6815 6422 6879 6426
rect 18020 6422 18084 6486
rect 2557 6197 2621 6201
rect 2557 6141 2561 6197
rect 2561 6141 2617 6197
rect 2617 6141 2621 6197
rect 2557 6137 2621 6141
rect 2706 6137 2770 6201
rect -1218 5525 -1154 5589
rect 109 5585 173 5589
rect 109 5529 113 5585
rect 113 5529 169 5585
rect 169 5529 173 5585
rect 109 5525 173 5529
rect 5723 5506 5787 5570
rect 17324 5506 17388 5570
rect 1695 5169 1759 5233
rect 879 5031 943 5095
rect 11770 5064 11834 5068
rect 11770 5008 11774 5064
rect 11774 5008 11830 5064
rect 11830 5008 11834 5064
rect 11770 5004 11834 5008
rect 1884 4903 1948 4967
rect 2557 4963 2621 4967
rect 2557 4907 2561 4963
rect 2561 4907 2617 4963
rect 2617 4907 2621 4963
rect 2557 4903 2621 4907
rect 3592 4903 3656 4967
rect 879 4744 943 4808
rect 1287 4744 1351 4808
rect 1695 4744 1759 4808
rect 2103 4744 2167 4808
rect -522 4588 -458 4652
rect 1884 4588 1948 4652
rect 1287 4450 1351 4514
rect 2103 4312 2167 4376
rect 3592 4187 3656 4251
rect 3822 4187 3886 4251
rect 4230 4187 4294 4251
rect 4434 4187 4498 4251
rect 5723 4244 5787 4248
rect 5723 4188 5727 4244
rect 5727 4188 5783 4244
rect 5783 4188 5787 4244
rect 5723 4184 5787 4188
rect 6345 4244 6409 4248
rect 6345 4188 6349 4244
rect 6349 4188 6405 4244
rect 6405 4188 6409 4244
rect 6345 4184 6409 4188
rect 3592 3471 3656 3535
rect 3822 3471 3886 3535
rect 4230 3471 4294 3535
rect 4443 3471 4507 3535
rect 4589 3436 4653 3500
rect 5723 3548 5787 3552
rect 5723 3492 5727 3548
rect 5727 3492 5783 3548
rect 5783 3492 5787 3548
rect 5723 3488 5787 3492
rect 6345 3548 6409 3552
rect 6345 3492 6349 3548
rect 6349 3492 6405 3548
rect 6405 3492 6409 3548
rect 6345 3488 6409 3492
rect 3735 3125 3799 3129
rect 3735 3069 3739 3125
rect 3739 3069 3795 3125
rect 3795 3069 3799 3125
rect 3735 3065 3799 3069
rect 4589 3065 4653 3129
rect 4230 2640 4294 2704
rect 4551 2700 4615 2704
rect 4551 2644 4555 2700
rect 4555 2644 4611 2700
rect 4611 2644 4615 2700
rect 4551 2640 4615 2644
rect -1218 2469 -1154 2533
rect 1700 2469 1764 2533
rect 1700 2113 1764 2177
rect 3735 2173 3799 2177
rect 3735 2117 3739 2173
rect 3739 2117 3795 2173
rect 3795 2117 3799 2173
rect 3735 2113 3799 2117
rect 4551 1748 4615 1752
rect 4551 1692 4555 1748
rect 4555 1692 4611 1748
rect 4611 1692 4615 1748
rect 4551 1688 4615 1692
rect 6616 1420 6680 1484
rect 10186 1420 10250 1484
rect 13755 1420 13819 1484
rect 14724 1420 14788 1484
rect 17324 1420 17388 1484
rect 2630 1076 2694 1140
rect 3735 1136 3799 1140
rect 3735 1080 3739 1136
rect 3739 1080 3795 1136
rect 3795 1080 3799 1136
rect 3735 1076 3799 1080
rect 6477 1076 6541 1140
rect 3105 681 3169 685
rect 3105 625 3109 681
rect 3109 625 3165 681
rect 3165 625 3169 681
rect 3105 621 3169 625
rect 3047 454 3111 518
rect 4551 514 4615 518
rect 4551 458 4555 514
rect 4555 458 4611 514
rect 4611 458 4615 514
rect 4551 454 4615 458
rect 6616 454 6680 518
rect 9965 564 10029 568
rect 9965 508 9969 564
rect 9969 508 10025 564
rect 10025 508 10029 564
rect 9965 504 10029 508
rect 10325 504 10389 568
rect 14172 504 14236 568
rect 14873 564 14937 568
rect 14873 508 14877 564
rect 14877 508 14933 564
rect 14933 508 14937 564
rect 14873 504 14937 508
rect 18020 504 18084 568
rect 1700 351 1764 415
rect 3948 355 4012 359
rect 3948 299 3952 355
rect 3952 299 4008 355
rect 4008 299 4012 355
rect 3948 295 4012 299
rect 4356 355 4420 359
rect 4356 299 4360 355
rect 4360 299 4416 355
rect 4416 299 4420 355
rect 4356 295 4420 299
rect 9827 -15 9891 49
rect 10749 45 10813 49
rect 10749 -11 10753 45
rect 10753 -11 10809 45
rect 10809 -11 10813 45
rect 10749 -15 10813 -11
rect 11057 45 11121 49
rect 11057 -11 11061 45
rect 11061 -11 11117 45
rect 11117 -11 11121 45
rect 11057 -15 11121 -11
rect 11365 45 11429 49
rect 11365 -11 11369 45
rect 11369 -11 11425 45
rect 11425 -11 11429 45
rect 11365 -15 11429 -11
rect 11673 45 11737 49
rect 11673 -11 11677 45
rect 11677 -11 11733 45
rect 11733 -11 11737 45
rect 11673 -15 11737 -11
rect 11981 45 12045 49
rect 11981 -11 11985 45
rect 11985 -11 12041 45
rect 12041 -11 12045 45
rect 11981 -15 12045 -11
rect 12289 45 12353 49
rect 12289 -11 12293 45
rect 12293 -11 12349 45
rect 12349 -11 12353 45
rect 12289 -15 12353 -11
rect 12597 45 12661 49
rect 12597 -11 12601 45
rect 12601 -11 12657 45
rect 12657 -11 12661 45
rect 12597 -15 12661 -11
rect 12905 45 12969 49
rect 12905 -11 12909 45
rect 12909 -11 12965 45
rect 12965 -11 12969 45
rect 12905 -15 12969 -11
rect 13213 45 13277 49
rect 13213 -11 13217 45
rect 13217 -11 13273 45
rect 13273 -11 13277 45
rect 13213 -15 13277 -11
rect 13521 45 13585 49
rect 13521 -11 13525 45
rect 13525 -11 13581 45
rect 13581 -11 13585 45
rect 13521 -15 13585 -11
rect 13978 -15 14042 49
rect 14445 45 14509 49
rect 14445 -11 14449 45
rect 14449 -11 14505 45
rect 14505 -11 14509 45
rect 14445 -15 14509 -11
rect 10463 -164 10527 -100
rect 14310 -164 14374 -100
rect 14586 -164 14650 -100
rect -794 -522 -730 -458
rect -658 -522 -594 -458
rect -522 -522 -458 -458
rect 1700 -522 1764 -458
rect 3047 -522 3111 -458
rect 6616 -522 6680 -458
rect 10186 -522 10250 -458
rect 13755 -522 13819 -458
rect 14724 -522 14788 -458
rect 17324 -522 17388 -458
rect 17460 -522 17524 -458
rect 17596 -522 17660 -458
rect -794 -658 -730 -594
rect -658 -658 -594 -594
rect -522 -658 -458 -594
rect 17324 -658 17388 -594
rect 17460 -658 17524 -594
rect 17596 -658 17660 -594
rect -794 -794 -730 -730
rect -658 -794 -594 -730
rect -522 -794 -458 -730
rect 17324 -794 17388 -730
rect 17460 -794 17524 -730
rect 17596 -794 17660 -730
rect -1490 -1218 -1426 -1154
rect -1354 -1218 -1290 -1154
rect -1218 -1218 -1154 -1154
rect 2630 -1218 2694 -1154
rect 6477 -1218 6541 -1154
rect 9965 -1218 10029 -1154
rect 10325 -1218 10389 -1154
rect 14172 -1218 14236 -1154
rect 14873 -1218 14937 -1154
rect 18020 -1218 18084 -1154
rect 18156 -1218 18220 -1154
rect 18292 -1218 18356 -1154
rect -1490 -1354 -1426 -1290
rect -1354 -1354 -1290 -1290
rect -1218 -1354 -1154 -1290
rect 18020 -1354 18084 -1290
rect 18156 -1354 18220 -1290
rect 18292 -1354 18356 -1290
rect -1490 -1490 -1426 -1426
rect -1354 -1490 -1290 -1426
rect -1218 -1490 -1154 -1426
rect 18020 -1490 18084 -1426
rect 18156 -1490 18220 -1426
rect 18292 -1490 18356 -1426
<< metal4 >>
rect -1496 18902 -1148 18908
rect -1496 18838 -1490 18902
rect -1426 18838 -1354 18902
rect -1290 18838 -1218 18902
rect -1154 18838 -1148 18902
rect -1496 18766 -1148 18838
rect -1496 18702 -1490 18766
rect -1426 18702 -1354 18766
rect -1290 18702 -1218 18766
rect -1154 18702 -1148 18766
rect -1496 18630 -1148 18702
rect 18014 18902 18362 18908
rect 18014 18838 18020 18902
rect 18084 18838 18156 18902
rect 18220 18838 18292 18902
rect 18356 18838 18362 18902
rect 18014 18766 18362 18838
rect 18014 18702 18020 18766
rect 18084 18702 18156 18766
rect 18220 18702 18292 18766
rect 18356 18702 18362 18766
rect -1496 18566 -1490 18630
rect -1426 18566 -1354 18630
rect -1290 18566 -1218 18630
rect -1154 18566 -1148 18630
rect -1496 17024 -1148 18566
rect 3834 18630 3910 18636
rect 3834 18566 3840 18630
rect 3904 18566 3910 18630
rect -1496 16960 -1218 17024
rect -1154 16960 -1148 17024
rect -1496 7578 -1148 16960
rect -1496 7514 -1218 7578
rect -1154 7514 -1148 7578
rect -1496 6626 -1148 7514
rect -1496 6562 -1218 6626
rect -1154 6562 -1148 6626
rect -1496 5589 -1148 6562
rect -1496 5525 -1218 5589
rect -1154 5525 -1148 5589
rect -1496 2533 -1148 5525
rect -1496 2469 -1218 2533
rect -1154 2469 -1148 2533
rect -1496 -1154 -1148 2469
rect -800 18206 -452 18212
rect -800 18142 -794 18206
rect -730 18142 -658 18206
rect -594 18142 -522 18206
rect -458 18142 -452 18206
rect -800 18070 -452 18142
rect -800 18006 -794 18070
rect -730 18006 -658 18070
rect -594 18006 -522 18070
rect -458 18006 -452 18070
rect -800 17934 -452 18006
rect -800 17870 -794 17934
rect -730 17870 -658 17934
rect -594 17870 -522 17934
rect -458 17870 -452 17934
rect -800 14928 -452 17870
rect 2443 17934 2519 17940
rect 2443 17870 2449 17934
rect 2513 17870 2519 17934
rect -31 17176 45 17182
rect -31 17112 -25 17176
rect 39 17112 45 17176
rect -31 16670 45 17112
rect -40 16664 45 16670
rect -40 16600 -34 16664
rect 30 16600 45 16664
rect -40 16594 45 16600
rect 190 17176 266 17182
rect 190 17112 196 17176
rect 260 17112 266 17176
rect 190 16664 266 17112
rect 2443 17176 2519 17870
rect 3685 17934 3761 17940
rect 3685 17870 3691 17934
rect 3755 17870 3761 17934
rect 2443 17112 2449 17176
rect 2513 17112 2519 17176
rect 2443 16670 2519 17112
rect 190 16600 196 16664
rect 260 16600 266 16664
rect 190 16594 266 16600
rect 2434 16664 2519 16670
rect 2434 16600 2440 16664
rect 2504 16600 2519 16664
rect 2434 16594 2519 16600
rect 2589 17176 2665 17182
rect 2589 17112 2595 17176
rect 2659 17112 2665 17176
rect 2589 16664 2665 17112
rect 3685 17173 3761 17870
rect 3685 17109 3691 17173
rect 3755 17109 3761 17173
rect 3685 17103 3761 17109
rect 3834 17173 3910 18566
rect 5939 18630 6015 18636
rect 5939 18566 5945 18630
rect 6009 18566 6015 18630
rect 3834 17109 3840 17173
rect 3904 17109 3910 17173
rect 3834 17103 3910 17109
rect 5790 17934 5866 17940
rect 5790 17870 5796 17934
rect 5860 17870 5866 17934
rect 5790 17173 5866 17870
rect 5790 17109 5796 17173
rect 5860 17109 5866 17173
rect 5790 17103 5866 17109
rect 5939 17173 6015 18566
rect 10319 18630 10395 18636
rect 10319 18566 10325 18630
rect 10389 18566 10395 18630
rect 6915 17934 6991 17940
rect 6915 17870 6921 17934
rect 6985 17870 6991 17934
rect 6915 17384 6991 17870
rect 6915 17320 6921 17384
rect 6985 17320 6991 17384
rect 6915 17314 6991 17320
rect 10180 17934 10256 17940
rect 10180 17870 10186 17934
rect 10250 17870 10256 17934
rect 10180 17384 10256 17870
rect 10180 17320 10186 17384
rect 10250 17320 10256 17384
rect 10180 17314 10256 17320
rect 5939 17109 5945 17173
rect 6009 17109 6015 17173
rect 5939 17103 6015 17109
rect 10319 17173 10395 18566
rect 14166 18630 14242 18636
rect 14166 18566 14172 18630
rect 14236 18566 14242 18630
rect 10319 17109 10325 17173
rect 10389 17109 10395 17173
rect 10319 17103 10395 17109
rect 11832 17934 11908 17940
rect 11832 17870 11838 17934
rect 11902 17870 11908 17934
rect 2589 16600 2595 16664
rect 2659 16600 2665 16664
rect -800 14864 -522 14928
rect -458 14864 -452 14928
rect -800 13192 -452 14864
rect 2434 14928 2510 14934
rect 2434 14864 2440 14928
rect 2504 14864 2510 14928
rect -800 13128 -522 13192
rect -458 13128 -452 13192
rect -800 11456 -452 13128
rect -800 11392 -522 11456
rect -458 11392 -452 11456
rect -800 9720 -452 11392
rect -40 13192 36 13198
rect -40 13128 -34 13192
rect 30 13128 36 13192
rect -40 11456 36 13128
rect -40 11392 -34 11456
rect 30 11392 36 11456
rect -40 11386 36 11392
rect 2434 13192 2510 14864
rect 2589 14928 2665 16600
rect 2589 14864 2595 14928
rect 2659 14864 2665 14928
rect 2589 14858 2665 14864
rect 11832 16695 11908 17870
rect 11832 16631 11838 16695
rect 11902 16631 11908 16695
rect 11832 14959 11908 16631
rect 13749 17934 13825 17940
rect 13749 17870 13755 17934
rect 13819 17870 13825 17934
rect 13749 16695 13825 17870
rect 14166 17173 14242 18566
rect 18014 18630 18362 18702
rect 18014 18566 18020 18630
rect 18084 18566 18156 18630
rect 18220 18566 18292 18630
rect 18356 18566 18362 18630
rect 17318 18206 17666 18212
rect 17318 18142 17324 18206
rect 17388 18142 17460 18206
rect 17524 18142 17596 18206
rect 17660 18142 17666 18206
rect 17318 18070 17666 18142
rect 17318 18006 17324 18070
rect 17388 18006 17460 18070
rect 17524 18006 17596 18070
rect 17660 18006 17666 18070
rect 16531 17934 16607 17940
rect 16531 17870 16537 17934
rect 16601 17870 16607 17934
rect 16531 17384 16607 17870
rect 16531 17320 16537 17384
rect 16601 17320 16607 17384
rect 16531 17314 16607 17320
rect 17318 17934 17666 18006
rect 17318 17870 17324 17934
rect 17388 17870 17460 17934
rect 17524 17870 17596 17934
rect 17660 17870 17666 17934
rect 17318 17384 17666 17870
rect 17318 17320 17324 17384
rect 17388 17320 17666 17384
rect 14166 17109 14172 17173
rect 14236 17109 14242 17173
rect 14166 17103 14242 17109
rect 13749 16631 13755 16695
rect 13819 16631 13825 16695
rect 13749 16625 13825 16631
rect 11832 14895 11838 14959
rect 11902 14895 11908 14959
rect 2434 13128 2440 13192
rect 2504 13128 2510 13192
rect 2434 11456 2510 13128
rect 2434 11392 2440 11456
rect 2504 11392 2510 11456
rect -800 9656 -522 9720
rect -458 9656 -452 9720
rect -800 7984 -452 9656
rect -800 7920 -522 7984
rect -458 7920 -452 7984
rect -800 4652 -452 7920
rect -40 9720 36 9726
rect -40 9656 -34 9720
rect 30 9656 36 9720
rect -40 7984 36 9656
rect 2434 9720 2510 11392
rect 2434 9656 2440 9720
rect 2504 9656 2510 9720
rect -40 7920 -34 7984
rect 30 7920 36 7984
rect -40 7914 36 7920
rect 2230 7984 2306 7990
rect 2230 7920 2236 7984
rect 2300 7920 2306 7984
rect 103 7578 179 7584
rect 103 7514 109 7578
rect 173 7514 179 7578
rect 103 6626 179 7514
rect 2230 7153 2306 7920
rect 2434 7984 2510 9656
rect 11832 13223 11908 14895
rect 11832 13159 11838 13223
rect 11902 13159 11908 13223
rect 11832 11487 11908 13159
rect 11832 11423 11838 11487
rect 11902 11423 11908 11487
rect 11832 9751 11908 11423
rect 11832 9687 11838 9751
rect 11902 9687 11908 9751
rect 11832 8015 11908 9687
rect 2434 7920 2440 7984
rect 2504 7920 2510 7984
rect 2434 7159 2510 7920
rect 5939 8001 6015 8007
rect 5939 7937 5945 8001
rect 6009 7937 6015 8001
rect 2230 7089 2236 7153
rect 2300 7089 2306 7153
rect 2230 7083 2306 7089
rect 2402 7153 2510 7159
rect 2402 7089 2408 7153
rect 2472 7089 2510 7153
rect 2402 7083 2510 7089
rect 2700 7153 2776 7159
rect 2700 7089 2706 7153
rect 2770 7089 2776 7153
rect 103 6562 109 6626
rect 173 6562 179 6626
rect 103 5589 179 6562
rect 103 5525 109 5589
rect 173 5525 179 5589
rect 103 5519 179 5525
rect 2551 6201 2627 6207
rect 2551 6137 2557 6201
rect 2621 6137 2627 6201
rect 1689 5233 1765 5239
rect 1689 5169 1695 5233
rect 1759 5169 1765 5233
rect 873 5095 949 5101
rect 873 5031 879 5095
rect 943 5031 949 5095
rect 873 4808 949 5031
rect 873 4744 879 4808
rect 943 4744 949 4808
rect 873 4738 949 4744
rect 1281 4808 1357 4814
rect 1281 4744 1287 4808
rect 1351 4744 1357 4808
rect -800 4588 -522 4652
rect -458 4588 -452 4652
rect -800 -458 -452 4588
rect 1281 4514 1357 4744
rect 1689 4808 1765 5169
rect 1689 4744 1695 4808
rect 1759 4744 1765 4808
rect 1689 4738 1765 4744
rect 1878 4967 1954 4973
rect 1878 4903 1884 4967
rect 1948 4903 1954 4967
rect 1878 4652 1954 4903
rect 2551 4967 2627 6137
rect 2700 6201 2776 7089
rect 5939 7142 6015 7937
rect 11832 7951 11838 8015
rect 11902 7951 11908 8015
rect 5939 7078 5945 7142
rect 6009 7078 6015 7142
rect 5939 7072 6015 7078
rect 6809 7142 6889 7148
rect 6809 7078 6819 7142
rect 6883 7078 6889 7142
rect 6809 7072 6889 7078
rect 2700 6137 2706 6201
rect 2770 6137 2776 6201
rect 2700 6131 2776 6137
rect 6339 6486 6415 6492
rect 6339 6422 6345 6486
rect 6409 6422 6415 6486
rect 5717 5570 5793 5576
rect 5717 5506 5723 5570
rect 5787 5506 5793 5570
rect 2551 4903 2557 4967
rect 2621 4903 2627 4967
rect 2551 4897 2627 4903
rect 3586 4967 3662 4973
rect 3586 4903 3592 4967
rect 3656 4903 3662 4967
rect 1878 4588 1884 4652
rect 1948 4588 1954 4652
rect 1878 4582 1954 4588
rect 2097 4808 2173 4814
rect 2097 4744 2103 4808
rect 2167 4744 2173 4808
rect 1281 4450 1287 4514
rect 1351 4450 1357 4514
rect 1281 4444 1357 4450
rect 2097 4376 2173 4744
rect 2097 4312 2103 4376
rect 2167 4312 2173 4376
rect 2097 4306 2173 4312
rect 3586 4251 3662 4903
rect 3586 4187 3592 4251
rect 3656 4187 3662 4251
rect 3586 3535 3662 4187
rect 3586 3471 3592 3535
rect 3656 3471 3662 3535
rect 3586 3465 3662 3471
rect 3816 4251 3892 4257
rect 3816 4187 3822 4251
rect 3886 4187 3892 4251
rect 3816 3535 3892 4187
rect 3816 3471 3822 3535
rect 3886 3471 3892 3535
rect 3816 3465 3892 3471
rect 4224 4251 4300 4257
rect 4224 4187 4230 4251
rect 4294 4187 4300 4251
rect 4224 3535 4300 4187
rect 4428 4251 4513 4257
rect 4428 4187 4434 4251
rect 4498 4187 4513 4251
rect 4428 4181 4513 4187
rect 4224 3471 4230 3535
rect 4294 3471 4300 3535
rect 3729 3129 3805 3135
rect 3729 3065 3735 3129
rect 3799 3065 3805 3129
rect 1694 2533 1770 2539
rect 1694 2469 1700 2533
rect 1764 2469 1770 2533
rect 1694 2177 1770 2469
rect 1694 2113 1700 2177
rect 1764 2113 1770 2177
rect 1694 2107 1770 2113
rect 3729 2177 3805 3065
rect 4224 2704 4300 3471
rect 4437 3535 4513 4181
rect 4437 3471 4443 3535
rect 4507 3471 4513 3535
rect 5717 4248 5793 5506
rect 5717 4184 5723 4248
rect 5787 4184 5793 4248
rect 5717 3552 5793 4184
rect 4437 3465 4513 3471
rect 4583 3500 4659 3506
rect 4583 3436 4589 3500
rect 4653 3436 4659 3500
rect 5717 3488 5723 3552
rect 5787 3488 5793 3552
rect 5717 3482 5793 3488
rect 6339 4248 6415 6422
rect 6809 6486 6885 7072
rect 6809 6422 6815 6486
rect 6879 6422 6885 6486
rect 6809 6416 6885 6422
rect 11832 5074 11908 7951
rect 11764 5068 11908 5074
rect 11764 5004 11770 5068
rect 11834 5004 11908 5068
rect 11764 4998 11908 5004
rect 17318 5570 17666 17320
rect 17318 5506 17324 5570
rect 17388 5506 17666 5570
rect 6339 4184 6345 4248
rect 6409 4184 6415 4248
rect 6339 3552 6415 4184
rect 6339 3488 6345 3552
rect 6409 3488 6415 3552
rect 6339 3482 6415 3488
rect 4583 3129 4659 3436
rect 4583 3065 4589 3129
rect 4653 3065 4659 3129
rect 4583 3059 4659 3065
rect 4224 2640 4230 2704
rect 4294 2640 4300 2704
rect 4224 2634 4300 2640
rect 4545 2704 4621 2710
rect 4545 2640 4551 2704
rect 4615 2640 4621 2704
rect 3729 2113 3735 2177
rect 3799 2113 3805 2177
rect 2624 1140 2700 1146
rect 2624 1076 2630 1140
rect 2694 1076 2700 1140
rect -800 -522 -794 -458
rect -730 -522 -658 -458
rect -594 -522 -522 -458
rect -458 -522 -452 -458
rect -800 -594 -452 -522
rect 1694 415 1770 421
rect 1694 351 1700 415
rect 1764 351 1770 415
rect 1694 -458 1770 351
rect 1694 -522 1700 -458
rect 1764 -522 1770 -458
rect 1694 -528 1770 -522
rect -800 -658 -794 -594
rect -730 -658 -658 -594
rect -594 -658 -522 -594
rect -458 -658 -452 -594
rect -800 -730 -452 -658
rect -800 -794 -794 -730
rect -730 -794 -658 -730
rect -594 -794 -522 -730
rect -458 -794 -452 -730
rect -800 -800 -452 -794
rect -1496 -1218 -1490 -1154
rect -1426 -1218 -1354 -1154
rect -1290 -1218 -1218 -1154
rect -1154 -1218 -1148 -1154
rect -1496 -1290 -1148 -1218
rect 2624 -1154 2700 1076
rect 3729 1140 3805 2113
rect 3729 1076 3735 1140
rect 3799 1076 3805 1140
rect 3729 1070 3805 1076
rect 4545 1752 4621 2640
rect 4545 1688 4551 1752
rect 4615 1688 4621 1752
rect 3099 685 3175 691
rect 3099 621 3105 685
rect 3169 662 3175 685
rect 3169 621 3255 662
rect 3099 586 3255 621
rect 3041 518 3117 524
rect 3041 454 3047 518
rect 3111 454 3117 518
rect 3041 -458 3117 454
rect 3041 -522 3047 -458
rect 3111 -522 3117 -458
rect 3041 -528 3117 -522
rect 2624 -1218 2630 -1154
rect 2694 -1218 2700 -1154
rect 2624 -1224 2700 -1218
rect -1496 -1354 -1490 -1290
rect -1426 -1354 -1354 -1290
rect -1290 -1354 -1218 -1290
rect -1154 -1354 -1148 -1290
rect -1496 -1426 -1148 -1354
rect -1496 -1490 -1490 -1426
rect -1426 -1490 -1354 -1426
rect -1290 -1490 -1218 -1426
rect -1154 -1490 -1148 -1426
rect -1496 -1496 -1148 -1490
rect 3179 -1496 3255 586
rect 4545 518 4621 1688
rect 6610 1484 6686 1490
rect 6610 1420 6616 1484
rect 6680 1420 6686 1484
rect 4545 454 4551 518
rect 4615 454 4621 518
rect 4545 448 4621 454
rect 6471 1140 6547 1146
rect 6471 1076 6477 1140
rect 6541 1076 6547 1140
rect 3942 359 4018 365
rect 3942 295 3948 359
rect 4012 295 4018 359
rect 3942 -1496 4018 295
rect 4350 359 4426 365
rect 4350 295 4356 359
rect 4420 295 4426 359
rect 4350 -1496 4426 295
rect 6471 -1154 6547 1076
rect 6610 518 6686 1420
rect 10180 1484 10256 1490
rect 10180 1420 10186 1484
rect 10250 1420 10256 1484
rect 6610 454 6616 518
rect 6680 454 6686 518
rect 6610 -458 6686 454
rect 9959 568 10035 574
rect 9959 504 9965 568
rect 10029 504 10035 568
rect 6610 -522 6616 -458
rect 6680 -522 6686 -458
rect 6610 -528 6686 -522
rect 9821 49 9897 55
rect 9821 -15 9827 49
rect 9891 -15 9897 49
rect 6471 -1218 6477 -1154
rect 6541 -1218 6547 -1154
rect 6471 -1224 6547 -1218
rect 9821 -1496 9897 -15
rect 9959 -1154 10035 504
rect 10180 -458 10256 1420
rect 13749 1484 13825 1490
rect 13749 1420 13755 1484
rect 13819 1420 13825 1484
rect 10180 -522 10186 -458
rect 10250 -522 10256 -458
rect 10180 -528 10256 -522
rect 10319 568 10395 574
rect 10319 504 10325 568
rect 10389 504 10395 568
rect 9959 -1218 9965 -1154
rect 10029 -1218 10035 -1154
rect 9959 -1224 10035 -1218
rect 10319 -1154 10395 504
rect 10743 49 10819 55
rect 10743 -15 10749 49
rect 10813 -15 10819 49
rect 10319 -1218 10325 -1154
rect 10389 -1218 10395 -1154
rect 10319 -1224 10395 -1218
rect 10457 -100 10533 -94
rect 10457 -164 10463 -100
rect 10527 -164 10533 -100
rect 10457 -1496 10533 -164
rect 10743 -1496 10819 -15
rect 11051 49 11127 55
rect 11051 -15 11057 49
rect 11121 -15 11127 49
rect 11051 -1496 11127 -15
rect 11359 49 11435 55
rect 11359 -15 11365 49
rect 11429 -15 11435 49
rect 11359 -1496 11435 -15
rect 11667 49 11743 55
rect 11667 -15 11673 49
rect 11737 -15 11743 49
rect 11667 -1496 11743 -15
rect 11975 49 12051 55
rect 11975 -15 11981 49
rect 12045 -15 12051 49
rect 11975 -1496 12051 -15
rect 12283 49 12359 55
rect 12283 -15 12289 49
rect 12353 -15 12359 49
rect 12283 -1496 12359 -15
rect 12591 49 12667 55
rect 12591 -15 12597 49
rect 12661 -15 12667 49
rect 12591 -1496 12667 -15
rect 12899 49 12975 55
rect 12899 -15 12905 49
rect 12969 -15 12975 49
rect 12899 -1496 12975 -15
rect 13207 49 13283 55
rect 13207 -15 13213 49
rect 13277 -15 13283 49
rect 13207 -1496 13283 -15
rect 13515 49 13591 55
rect 13515 -15 13521 49
rect 13585 -15 13591 49
rect 13515 -1496 13591 -15
rect 13749 -458 13825 1420
rect 14718 1484 14794 1490
rect 14718 1420 14724 1484
rect 14788 1420 14794 1484
rect 14166 568 14242 574
rect 14166 504 14172 568
rect 14236 504 14242 568
rect 13749 -522 13755 -458
rect 13819 -522 13825 -458
rect 13749 -528 13825 -522
rect 13972 49 14048 55
rect 13972 -15 13978 49
rect 14042 -15 14048 49
rect 13972 -1496 14048 -15
rect 14166 -1154 14242 504
rect 14439 49 14515 55
rect 14439 -15 14445 49
rect 14509 44 14515 49
rect 14509 -15 14518 44
rect 14439 -32 14518 -15
rect 14166 -1218 14172 -1154
rect 14236 -1218 14242 -1154
rect 14166 -1224 14242 -1218
rect 14304 -100 14380 -94
rect 14304 -164 14310 -100
rect 14374 -164 14380 -100
rect 14304 -1496 14380 -164
rect 14442 -1496 14518 -32
rect 14580 -100 14656 -94
rect 14580 -164 14586 -100
rect 14650 -164 14656 -100
rect 14580 -1496 14656 -164
rect 14718 -458 14794 1420
rect 17318 1484 17666 5506
rect 17318 1420 17324 1484
rect 17388 1420 17666 1484
rect 14718 -522 14724 -458
rect 14788 -522 14794 -458
rect 14718 -528 14794 -522
rect 14867 568 14943 574
rect 14867 504 14873 568
rect 14937 504 14943 568
rect 14867 -1154 14943 504
rect 17318 -458 17666 1420
rect 17318 -522 17324 -458
rect 17388 -522 17460 -458
rect 17524 -522 17596 -458
rect 17660 -522 17666 -458
rect 17318 -594 17666 -522
rect 17318 -658 17324 -594
rect 17388 -658 17460 -594
rect 17524 -658 17596 -594
rect 17660 -658 17666 -594
rect 17318 -730 17666 -658
rect 17318 -794 17324 -730
rect 17388 -794 17460 -730
rect 17524 -794 17596 -730
rect 17660 -794 17666 -730
rect 17318 -800 17666 -794
rect 18014 6486 18362 18566
rect 18014 6422 18020 6486
rect 18084 6422 18362 6486
rect 18014 568 18362 6422
rect 18014 504 18020 568
rect 18084 504 18362 568
rect 14867 -1218 14873 -1154
rect 14937 -1218 14943 -1154
rect 14867 -1224 14943 -1218
rect 18014 -1154 18362 504
rect 18014 -1218 18020 -1154
rect 18084 -1218 18156 -1154
rect 18220 -1218 18292 -1154
rect 18356 -1218 18362 -1154
rect 18014 -1290 18362 -1218
rect 18014 -1354 18020 -1290
rect 18084 -1354 18156 -1290
rect 18220 -1354 18292 -1290
rect 18356 -1354 18362 -1290
rect 18014 -1426 18362 -1354
rect 18014 -1490 18020 -1426
rect 18084 -1490 18156 -1426
rect 18220 -1490 18292 -1426
rect 18356 -1490 18362 -1426
rect 18014 -1496 18362 -1490
use sky130_rom_krom_rom_base_array  sky130_rom_krom_rom_base_array_0
timestamp 1581321262
transform 1 0 6825 0 1 7110
box 0 -84 10041 10269
use sky130_rom_krom_rom_bitline_inverter  sky130_rom_krom_rom_bitline_inverter_0
timestamp 1581321264
transform 0 -1 16639 1 0 5208
box 136 -79 1879 9887
use sky130_rom_krom_rom_column_decode  sky130_rom_krom_rom_column_decode_0
timestamp 1581321264
transform 1 0 3626 0 1 250
box -39 44 3105 4237
use sky130_rom_krom_rom_column_mux_array  sky130_rom_krom_rom_column_mux_array_0
timestamp 1581321264
transform 1 0 6873 0 1 3062
box 0 382 9843 2041
use sky130_rom_krom_rom_control_logic  sky130_rom_krom_rom_control_logic_0
timestamp 1581321264
transform 1 0 456 0 1 383
box -36 -49 2966 4286
use sky130_rom_krom_rom_output_buffer  sky130_rom_krom_rom_output_buffer_0
timestamp 1581321264
transform 0 1 9977 -1 0 1782
box 44 -50 1800 5023
use sky130_rom_krom_rom_row_decode  sky130_rom_krom_rom_row_decode_0
timestamp 1581321264
transform 1 0 0 0 1 4699
box -39 44 6731 12713
<< labels >>
rlabel metal4 s 3179 -1496 3255 -1420 4 cs0
port 3 nsew
rlabel metal3 s -1496 1366 -1420 1442 4 clk0
port 5 nsew
rlabel metal4 s 9821 -1496 9897 -1420 4 dout0[0]
port 7 nsew
rlabel metal4 s 10457 -1496 10533 -1420 4 dout0[1]
port 9 nsew
rlabel metal4 s 10743 -1496 10819 -1420 4 dout0[2]
port 11 nsew
rlabel metal4 s 11051 -1496 11127 -1420 4 dout0[3]
port 13 nsew
rlabel metal4 s 11359 -1496 11435 -1420 4 dout0[4]
port 15 nsew
rlabel metal4 s 11667 -1496 11743 -1420 4 dout0[5]
port 17 nsew
rlabel metal4 s 11975 -1496 12051 -1420 4 dout0[6]
port 19 nsew
rlabel metal4 s 12283 -1496 12359 -1420 4 dout0[7]
port 21 nsew
rlabel metal4 s 12591 -1496 12667 -1420 4 dout0[8]
port 23 nsew
rlabel metal4 s 12899 -1496 12975 -1420 4 dout0[9]
port 25 nsew
rlabel metal4 s 13207 -1496 13283 -1420 4 dout0[10]
port 27 nsew
rlabel metal4 s 13515 -1496 13591 -1420 4 dout0[11]
port 29 nsew
rlabel metal4 s 13972 -1496 14048 -1420 4 dout0[12]
port 31 nsew
rlabel metal4 s 14304 -1496 14380 -1420 4 dout0[13]
port 33 nsew
rlabel metal4 s 14442 -1496 14518 -1420 4 dout0[14]
port 35 nsew
rlabel metal4 s 14580 -1496 14656 -1420 4 dout0[15]
port 37 nsew
rlabel metal4 s 3942 -1496 4018 -1420 4 addr0[0]
port 39 nsew
rlabel metal4 s 4350 -1496 4426 -1420 4 addr0[1]
port 41 nsew
rlabel metal3 s -1496 4738 -1420 4814 4 addr0[2]
port 43 nsew
rlabel metal3 s -1496 4887 -1420 4963 4 addr0[3]
port 45 nsew
rlabel metal3 s -1496 5025 -1420 5101 4 addr0[4]
port 47 nsew
rlabel metal3 s -1496 4444 -1420 4520 4 addr0[5]
port 49 nsew
rlabel metal3 s -1496 5163 -1420 5239 4 addr0[6]
port 51 nsew
rlabel metal3 s -1496 4306 -1420 4382 4 addr0[7]
port 53 nsew
rlabel metal3 s -1496 18560 18362 18908 4 vccd1
port 55 nsew
rlabel metal4 s -1496 -1496 -1148 18908 4 vccd1
port 55 nsew
rlabel metal3 s -1496 -1496 18362 -1148 4 vccd1
port 55 nsew
rlabel metal4 s 18014 -1496 18362 18908 4 vccd1
port 55 nsew
rlabel metal4 s -800 -800 -452 18212 4 vssd1
port 57 nsew
rlabel metal4 s 17318 -800 17666 18212 4 vssd1
port 57 nsew
rlabel metal3 s -800 -800 17666 -452 4 vssd1
port 57 nsew
rlabel metal3 s -800 17864 17666 18212 4 vssd1
port 57 nsew
<< properties >>
string FIXED_BBOX 18286 -1491 18362 -1425
<< end >>
