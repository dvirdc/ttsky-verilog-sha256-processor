magic
tech sky130A
magscale 1 2
timestamp 1581398725
<< checkpaint >>
rect -1299 -1216 9271 6517
<< locali >>
rect 2361 4883 2395 4899
rect 7959 4849 7993 4883
rect 2361 4833 2395 4849
rect 2361 4679 2395 4695
rect 7959 4645 7993 4679
rect 2361 4629 2395 4645
rect 2361 4475 2395 4491
rect 7959 4441 7993 4475
rect 2361 4425 2395 4441
rect 2361 4271 2395 4287
rect 7959 4237 7993 4271
rect 2361 4221 2395 4237
rect 2361 4067 2395 4083
rect 7959 4033 7993 4067
rect 2361 4017 2395 4033
rect 2361 3863 2395 3879
rect 7959 3829 7993 3863
rect 2361 3813 2395 3829
rect 2361 3659 2395 3675
rect 7959 3625 7993 3659
rect 2361 3609 2395 3625
rect 2361 3455 2395 3471
rect 7959 3421 7993 3455
rect 2361 3405 2395 3421
rect 321 60 387 94
rect 729 60 795 94
rect 1137 60 1203 94
<< viali >>
rect 2361 4849 2395 4883
rect 2361 4645 2395 4679
rect 2361 4441 2395 4475
rect 2361 4237 2395 4271
rect 2361 4033 2395 4067
rect 2361 3829 2395 3863
rect 2361 3625 2395 3659
rect 2361 3421 2395 3455
<< metal1 >>
rect 1877 5229 1905 5257
rect 2749 4972 2777 5000
rect 3997 4972 4025 5000
rect 5595 4972 5623 5000
rect 7243 4972 7271 5000
rect 2349 4883 2407 4889
rect 2349 4880 2361 4883
rect 2259 4852 2361 4880
rect 2349 4849 2361 4852
rect 2395 4849 2407 4883
rect 2349 4843 2407 4849
rect 2349 4679 2407 4685
rect 2349 4676 2361 4679
rect 2259 4648 2361 4676
rect 2349 4645 2361 4648
rect 2395 4645 2407 4679
rect 2349 4639 2407 4645
rect 2349 4475 2407 4481
rect 2349 4472 2361 4475
rect 2259 4444 2361 4472
rect 2349 4441 2361 4444
rect 2395 4441 2407 4475
rect 2349 4435 2407 4441
rect 2349 4271 2407 4277
rect 2349 4268 2361 4271
rect 2259 4240 2361 4268
rect 2349 4237 2361 4240
rect 2395 4237 2407 4271
rect 2349 4231 2407 4237
rect 2349 4067 2407 4073
rect 2349 4064 2361 4067
rect 2259 4036 2361 4064
rect 2349 4033 2361 4036
rect 2395 4033 2407 4067
rect 2349 4027 2407 4033
rect 2349 3863 2407 3869
rect 2349 3860 2361 3863
rect 2259 3832 2361 3860
rect 2349 3829 2361 3832
rect 2395 3829 2407 3863
rect 2349 3823 2407 3829
rect 2349 3659 2407 3665
rect 2349 3656 2361 3659
rect 2259 3628 2361 3656
rect 2349 3625 2361 3628
rect 2395 3625 2407 3659
rect 2349 3619 2407 3625
rect 2349 3455 2407 3461
rect 2349 3452 2361 3455
rect 2259 3424 2361 3452
rect 2349 3421 2361 3424
rect 2395 3421 2407 3455
rect 2349 3415 2407 3421
rect 2749 3256 2777 3284
rect 3997 3256 4025 3284
rect 5595 3256 5623 3284
rect 7243 3256 7271 3284
rect 298 3199 304 3251
rect 356 3199 362 3251
rect 502 3199 508 3251
rect 560 3199 566 3251
rect 706 3199 712 3251
rect 764 3199 770 3251
rect 910 3199 916 3251
rect 968 3199 974 3251
rect 1114 3199 1120 3251
rect 1172 3199 1178 3251
rect 1318 3199 1324 3251
rect 1376 3199 1382 3251
rect 316 3138 344 3199
rect 298 3086 304 3138
rect 356 3086 362 3138
rect 438 3086 444 3138
rect 496 3126 502 3138
rect 520 3126 548 3199
rect 724 3138 752 3199
rect 496 3098 548 3126
rect 496 3086 502 3098
rect 706 3086 712 3138
rect 764 3086 770 3138
rect 846 3086 852 3138
rect 904 3126 910 3138
rect 928 3126 956 3199
rect 1132 3138 1160 3199
rect 904 3098 956 3126
rect 904 3086 910 3098
rect 1114 3086 1120 3138
rect 1172 3086 1178 3138
rect 1254 3086 1260 3138
rect 1312 3126 1318 3138
rect 1336 3126 1364 3199
rect 1312 3098 1364 3126
rect 1312 3086 1318 3098
rect 127 2833 155 2861
rect 1351 2408 1379 2436
rect 127 2160 1351 2188
rect 127 1881 155 1909
rect 1351 1456 1379 1484
rect 127 844 155 872
rect 1351 222 1379 250
<< via1 >>
rect 304 3199 356 3251
rect 508 3199 560 3251
rect 712 3199 764 3251
rect 916 3199 968 3251
rect 1120 3199 1172 3251
rect 1324 3199 1376 3251
rect 304 3086 356 3138
rect 444 3086 496 3138
rect 712 3086 764 3138
rect 852 3086 904 3138
rect 1120 3086 1172 3138
rect 1260 3086 1312 3138
<< metal2 >>
rect 304 3251 356 3257
rect 304 3193 356 3199
rect 508 3251 560 3257
rect 508 3193 560 3199
rect 712 3251 764 3257
rect 712 3193 764 3199
rect 916 3251 968 3257
rect 916 3193 968 3199
rect 1120 3251 1172 3257
rect 1120 3193 1172 3199
rect 1324 3251 1376 3257
rect 1877 3253 1905 3281
rect 2241 3204 2305 3232
rect 1324 3193 1376 3199
rect 304 3138 356 3144
rect 304 3080 356 3086
rect 444 3138 496 3144
rect 444 3080 496 3086
rect 712 3138 764 3144
rect 712 3080 764 3086
rect 852 3138 904 3144
rect 852 3080 904 3086
rect 1120 3138 1172 3144
rect 1120 3080 1172 3086
rect 1260 3138 1312 3144
rect 1260 3080 1312 3086
<< metal3 >>
rect -31 4959 29 5019
rect 1235 4959 1295 5019
rect -31 3223 29 3283
rect 1235 3223 1295 3283
use sky130_rom_krom_rom_address_control_array  sky130_rom_krom_rom_address_control_array_0
timestamp 1581398725
transform 1 0 127 0 1 0
box -48 44 1319 3128
use sky130_rom_krom_rom_row_decode_array  sky130_rom_krom_rom_row_decode_array_0
timestamp 1581398725
transform 0 -1 2273 1 0 3192
box -6 -84 2065 2312
use sky130_rom_krom_rom_row_decode_wordline_buffer  sky130_rom_krom_rom_row_decode_wordline_buffer_0
timestamp 1581398725
transform 1 0 2301 0 1 3250
box 44 -50 5710 1831
<< labels >>
rlabel metal1 s 127 2160 1351 2188 4 clk
port 3 nsew
rlabel locali s 7976 3438 7976 3438 4 wl_0
port 4 nsew
rlabel locali s 7976 3642 7976 3642 4 wl_1
port 5 nsew
rlabel locali s 7976 3846 7976 3846 4 wl_2
port 6 nsew
rlabel locali s 7976 4050 7976 4050 4 wl_3
port 7 nsew
rlabel locali s 7976 4254 7976 4254 4 wl_4
port 8 nsew
rlabel locali s 7976 4458 7976 4458 4 wl_5
port 9 nsew
rlabel locali s 7976 4662 7976 4662 4 wl_6
port 10 nsew
rlabel locali s 7976 4866 7976 4866 4 wl_7
port 11 nsew
rlabel metal2 s 1877 3253 1905 3281 4 precharge
port 13 nsew
rlabel metal1 s 1877 5229 1905 5257 4 precharge_r
port 15 nsew
rlabel locali s 354 77 354 77 4 A0
port 16 nsew
rlabel locali s 762 77 762 77 4 A1
port 17 nsew
rlabel locali s 1170 77 1170 77 4 A2
port 18 nsew
rlabel metal1 s 127 1881 155 1909 4 vdd
port 20 nsew
rlabel metal1 s 3997 3256 4025 3284 4 vdd
port 20 nsew
rlabel metal2 s 2241 3204 2305 3232 4 vdd
port 20 nsew
rlabel metal1 s 127 844 155 872 4 vdd
port 20 nsew
rlabel metal1 s 7243 4972 7271 5000 4 vdd
port 20 nsew
rlabel metal1 s 3997 4972 4025 5000 4 vdd
port 20 nsew
rlabel metal1 s 7243 3256 7271 3284 4 vdd
port 20 nsew
rlabel metal1 s 127 2833 155 2861 4 vdd
port 20 nsew
rlabel metal1 s 2749 4972 2777 5000 4 gnd
port 22 nsew
rlabel metal1 s 5595 3256 5623 3284 4 gnd
port 22 nsew
rlabel metal3 s 1235 3223 1295 3283 4 gnd
port 22 nsew
rlabel metal3 s 1235 4959 1295 5019 4 gnd
port 22 nsew
rlabel metal1 s 1351 1456 1379 1484 4 gnd
port 22 nsew
rlabel metal1 s 1351 2408 1379 2436 4 gnd
port 22 nsew
rlabel metal3 s -31 3223 29 3283 4 gnd
port 22 nsew
rlabel metal1 s 2749 3256 2777 3284 4 gnd
port 22 nsew
rlabel metal3 s -31 4959 29 5019 4 gnd
port 22 nsew
rlabel metal1 s 1351 222 1379 250 4 gnd
port 22 nsew
rlabel metal1 s 5595 4972 5623 5000 4 gnd
port 22 nsew
<< properties >>
string FIXED_BBOX -31 0 7993 5257
<< end >>
