magic
tech sky130A
magscale 1 2
timestamp 1581320207
<< checkpaint >>
rect -1296 -1277 2204 3946
<< nwell >>
rect -36 1262 944 2686
<< pwell >>
rect 28 159 770 1077
rect 28 25 874 159
<< scnmos >>
rect 114 51 144 1051
rect 222 51 252 1051
rect 330 51 360 1051
rect 438 51 468 1051
rect 546 51 576 1051
rect 654 51 684 1051
<< scpmos >>
rect 114 1578 144 2578
rect 222 1578 252 2578
rect 330 1578 360 2578
rect 438 1578 468 2578
rect 546 1578 576 2578
rect 654 1578 684 2578
<< ndiff >>
rect 54 568 114 1051
rect 54 534 62 568
rect 96 534 114 568
rect 54 51 114 534
rect 144 568 222 1051
rect 144 534 166 568
rect 200 534 222 568
rect 144 51 222 534
rect 252 568 330 1051
rect 252 534 274 568
rect 308 534 330 568
rect 252 51 330 534
rect 360 568 438 1051
rect 360 534 382 568
rect 416 534 438 568
rect 360 51 438 534
rect 468 568 546 1051
rect 468 534 490 568
rect 524 534 546 568
rect 468 51 546 534
rect 576 568 654 1051
rect 576 534 598 568
rect 632 534 654 568
rect 576 51 654 534
rect 684 568 744 1051
rect 684 534 702 568
rect 736 534 744 568
rect 684 51 744 534
<< pdiff >>
rect 54 2095 114 2578
rect 54 2061 62 2095
rect 96 2061 114 2095
rect 54 1578 114 2061
rect 144 2095 222 2578
rect 144 2061 166 2095
rect 200 2061 222 2095
rect 144 1578 222 2061
rect 252 2095 330 2578
rect 252 2061 274 2095
rect 308 2061 330 2095
rect 252 1578 330 2061
rect 360 2095 438 2578
rect 360 2061 382 2095
rect 416 2061 438 2095
rect 360 1578 438 2061
rect 468 2095 546 2578
rect 468 2061 490 2095
rect 524 2061 546 2095
rect 468 1578 546 2061
rect 576 2095 654 2578
rect 576 2061 598 2095
rect 632 2061 654 2095
rect 576 1578 654 2061
rect 684 2095 744 2578
rect 684 2061 702 2095
rect 736 2061 744 2095
rect 684 1578 744 2061
<< ndiffc >>
rect 62 534 96 568
rect 166 534 200 568
rect 274 534 308 568
rect 382 534 416 568
rect 490 534 524 568
rect 598 534 632 568
rect 702 534 736 568
<< pdiffc >>
rect 62 2061 96 2095
rect 166 2061 200 2095
rect 274 2061 308 2095
rect 382 2061 416 2095
rect 490 2061 524 2095
rect 598 2061 632 2095
rect 702 2061 736 2095
<< psubdiff >>
rect 798 109 848 133
rect 798 75 806 109
rect 840 75 848 109
rect 798 51 848 75
<< nsubdiff >>
rect 798 2541 848 2565
rect 798 2507 806 2541
rect 840 2507 848 2541
rect 798 2483 848 2507
<< psubdiffcont >>
rect 806 75 840 109
<< nsubdiffcont >>
rect 806 2507 840 2541
<< poly >>
rect 114 2578 144 2604
rect 222 2578 252 2604
rect 330 2578 360 2604
rect 438 2578 468 2604
rect 546 2578 576 2604
rect 654 2578 684 2604
rect 114 1552 144 1578
rect 222 1552 252 1578
rect 330 1552 360 1578
rect 438 1552 468 1578
rect 546 1552 576 1578
rect 654 1552 684 1578
rect 114 1522 684 1552
rect 114 1348 144 1522
rect 48 1332 144 1348
rect 48 1298 64 1332
rect 98 1298 144 1332
rect 48 1282 144 1298
rect 114 1107 144 1282
rect 114 1077 684 1107
rect 114 1051 144 1077
rect 222 1051 252 1077
rect 330 1051 360 1077
rect 438 1051 468 1077
rect 546 1051 576 1077
rect 654 1051 684 1077
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
rect 438 25 468 51
rect 546 25 576 51
rect 654 25 684 51
<< polycont >>
rect 64 1298 98 1332
<< locali >>
rect 0 2612 908 2646
rect 62 2095 96 2612
rect 62 2045 96 2061
rect 166 2095 200 2111
rect 166 2011 200 2061
rect 274 2095 308 2612
rect 274 2045 308 2061
rect 382 2095 416 2111
rect 382 2011 416 2061
rect 490 2095 524 2612
rect 490 2045 524 2061
rect 598 2095 632 2111
rect 598 2011 632 2061
rect 702 2095 736 2612
rect 806 2541 840 2612
rect 806 2491 840 2507
rect 702 2045 736 2061
rect 166 1977 632 2011
rect 64 1332 98 1348
rect 64 1282 98 1298
rect 382 1332 416 1977
rect 382 1298 433 1332
rect 382 652 416 1298
rect 166 618 632 652
rect 62 568 96 584
rect 62 17 96 534
rect 166 568 200 618
rect 166 518 200 534
rect 274 568 308 584
rect 274 17 308 534
rect 382 568 416 618
rect 382 518 416 534
rect 490 568 524 584
rect 490 17 524 534
rect 598 568 632 618
rect 598 518 632 534
rect 702 568 736 584
rect 702 17 736 534
rect 806 109 840 125
rect 806 17 840 75
rect 0 -17 908 17
<< labels >>
rlabel locali s 81 1315 81 1315 4 A
port 1 nsew
rlabel locali s 416 1315 416 1315 4 Z
port 2 nsew
rlabel locali s 454 0 454 0 4 gnd
port 3 nsew
rlabel locali s 454 2629 454 2629 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 908 1994
<< end >>
