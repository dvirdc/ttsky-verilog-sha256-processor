magic
tech sky130A
magscale 1 2
timestamp 1581320207
<< checkpaint >>
rect -1296 -1277 1772 3946
<< nwell >>
rect -36 1262 512 2686
<< pwell >>
rect 28 159 338 477
rect 28 25 442 159
<< scnmos >>
rect 114 51 144 451
rect 222 51 252 451
<< scpmos >>
rect 114 1578 144 2578
rect 222 1578 252 2578
<< ndiff >>
rect 54 268 114 451
rect 54 234 62 268
rect 96 234 114 268
rect 54 51 114 234
rect 144 268 222 451
rect 144 234 166 268
rect 200 234 222 268
rect 144 51 222 234
rect 252 268 312 451
rect 252 234 270 268
rect 304 234 312 268
rect 252 51 312 234
<< pdiff >>
rect 54 2095 114 2578
rect 54 2061 62 2095
rect 96 2061 114 2095
rect 54 1578 114 2061
rect 144 2095 222 2578
rect 144 2061 166 2095
rect 200 2061 222 2095
rect 144 1578 222 2061
rect 252 2095 312 2578
rect 252 2061 270 2095
rect 304 2061 312 2095
rect 252 1578 312 2061
<< ndiffc >>
rect 62 234 96 268
rect 166 234 200 268
rect 270 234 304 268
<< pdiffc >>
rect 62 2061 96 2095
rect 166 2061 200 2095
rect 270 2061 304 2095
<< psubdiff >>
rect 366 109 416 133
rect 366 75 374 109
rect 408 75 416 109
rect 366 51 416 75
<< nsubdiff >>
rect 366 2541 416 2565
rect 366 2507 374 2541
rect 408 2507 416 2541
rect 366 2483 416 2507
<< psubdiffcont >>
rect 374 75 408 109
<< nsubdiffcont >>
rect 374 2507 408 2541
<< poly >>
rect 114 2578 144 2604
rect 222 2578 252 2604
rect 114 1552 144 1578
rect 222 1552 252 1578
rect 114 1522 252 1552
rect 114 1198 144 1522
rect 48 1182 144 1198
rect 48 1148 64 1182
rect 98 1148 144 1182
rect 48 1132 144 1148
rect 114 507 144 1132
rect 114 477 252 507
rect 114 451 144 477
rect 222 451 252 477
rect 114 25 144 51
rect 222 25 252 51
<< polycont >>
rect 64 1148 98 1182
<< locali >>
rect 0 2612 476 2646
rect 62 2095 96 2612
rect 62 2045 96 2061
rect 166 2095 200 2111
rect 64 1182 98 1198
rect 64 1132 98 1148
rect 166 1182 200 2061
rect 270 2095 304 2612
rect 374 2541 408 2612
rect 374 2491 408 2507
rect 270 2045 304 2061
rect 166 1148 217 1182
rect 62 268 96 284
rect 62 17 96 234
rect 166 268 200 1148
rect 166 218 200 234
rect 270 268 304 284
rect 270 17 304 234
rect 374 109 408 125
rect 374 17 408 75
rect 0 -17 476 17
<< labels >>
rlabel locali s 81 1165 81 1165 4 A
port 1 nsew
rlabel locali s 200 1165 200 1165 4 Z
port 2 nsew
rlabel locali s 238 0 238 0 4 gnd
port 3 nsew
rlabel locali s 238 2629 238 2629 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 476 1994
<< end >>
