magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1216 -1310 2020 1559
<< nwell >>
rect 428 -45 760 299
rect 510 -50 678 -45
<< pwell >>
rect 136 -17 260 185
<< scnmos >>
rect 162 69 234 99
<< scpmos >>
rect 482 69 706 99
<< ndiff >>
rect 162 151 234 159
rect 162 117 181 151
rect 215 117 234 151
rect 162 99 234 117
rect 162 51 234 69
rect 162 17 181 51
rect 215 17 234 51
rect 162 9 234 17
<< pdiff >>
rect 482 151 706 159
rect 482 117 577 151
rect 611 117 706 151
rect 482 99 706 117
rect 482 51 706 69
rect 482 17 577 51
rect 611 17 706 51
rect 482 9 706 17
<< ndiffc >>
rect 181 117 215 151
rect 181 17 215 51
<< pdiffc >>
rect 577 117 611 151
rect 577 17 611 51
<< poly >>
rect 44 101 110 117
rect 44 67 60 101
rect 94 99 110 101
rect 94 69 162 99
rect 234 69 482 99
rect 706 69 732 99
rect 94 67 110 69
rect 44 51 110 67
<< polycont >>
rect 60 67 94 101
<< locali >>
rect 181 151 215 167
rect 577 151 611 167
rect 165 117 181 151
rect 215 117 231 151
rect 561 117 577 151
rect 611 117 627 151
rect 60 101 94 117
rect 181 101 215 117
rect 577 101 611 117
rect 60 51 94 67
rect 165 17 181 51
rect 215 17 577 51
rect 611 17 742 51
<< viali >>
rect 181 117 215 151
rect 577 117 611 151
<< metal1 >>
rect 184 157 212 204
rect 580 157 608 204
rect 169 151 227 157
rect 169 117 181 151
rect 215 117 227 151
rect 169 111 227 117
rect 565 151 623 157
rect 565 117 577 151
rect 611 117 623 151
rect 565 111 623 117
rect 184 0 212 111
rect 580 0 608 111
<< labels >>
rlabel locali s 77 84 77 84 4 A
port 2 nsew
rlabel locali s 453 34 453 34 4 Z
port 3 nsew
rlabel metal1 s 184 0 212 204 4 gnd
port 5 nsew
rlabel metal1 s 580 0 608 204 4 vdd
port 7 nsew
<< properties >>
string FIXED_BBOX 510 -50 678 -45
<< end >>
