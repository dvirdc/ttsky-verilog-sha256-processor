magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1124 -1339 3139 11147
<< locali >>
rect 226 9639 260 9689
rect 1821 9639 1855 9705
rect 226 9605 297 9639
rect 226 9435 260 9485
rect 1821 9435 1855 9501
rect 226 9401 297 9435
rect 226 9231 260 9281
rect 1821 9231 1855 9297
rect 226 9197 297 9231
rect 226 9027 260 9077
rect 1821 9027 1855 9093
rect 226 8993 297 9027
rect 226 8823 260 8873
rect 1821 8823 1855 8889
rect 226 8789 297 8823
rect 226 8619 260 8669
rect 1821 8619 1855 8685
rect 226 8585 297 8619
rect 226 8415 260 8465
rect 1821 8415 1855 8481
rect 226 8381 297 8415
rect 226 8211 260 8261
rect 1821 8211 1855 8277
rect 226 8177 297 8211
rect 226 8007 260 8057
rect 1821 8007 1855 8073
rect 226 7973 297 8007
rect 226 7803 260 7853
rect 1821 7803 1855 7869
rect 226 7769 297 7803
rect 226 7599 260 7649
rect 1821 7599 1855 7665
rect 226 7565 297 7599
rect 226 7395 260 7445
rect 1821 7395 1855 7461
rect 226 7361 297 7395
rect 226 7191 260 7241
rect 1821 7191 1855 7257
rect 226 7157 297 7191
rect 226 6987 260 7037
rect 1821 6987 1855 7053
rect 226 6953 297 6987
rect 226 6783 260 6833
rect 1821 6783 1855 6849
rect 226 6749 297 6783
rect 226 6579 260 6629
rect 1821 6579 1855 6645
rect 226 6545 297 6579
rect 226 6375 260 6425
rect 1821 6375 1855 6441
rect 226 6341 297 6375
rect 226 6171 260 6221
rect 1821 6171 1855 6237
rect 226 6137 297 6171
rect 226 5967 260 6017
rect 1821 5967 1855 6033
rect 226 5933 297 5967
rect 226 5763 260 5813
rect 1821 5763 1855 5829
rect 226 5729 297 5763
rect 226 5559 260 5609
rect 1821 5559 1855 5625
rect 226 5525 297 5559
rect 226 5355 260 5405
rect 1821 5355 1855 5421
rect 226 5321 297 5355
rect 226 5151 260 5201
rect 1821 5151 1855 5217
rect 226 5117 297 5151
rect 226 4947 260 4997
rect 1821 4947 1855 5013
rect 226 4913 297 4947
rect 226 4743 260 4793
rect 1821 4743 1855 4809
rect 226 4709 297 4743
rect 226 4539 260 4589
rect 1821 4539 1855 4605
rect 226 4505 297 4539
rect 226 4335 260 4385
rect 1821 4335 1855 4401
rect 226 4301 297 4335
rect 226 4131 260 4181
rect 1821 4131 1855 4197
rect 226 4097 297 4131
rect 226 3927 260 3977
rect 1821 3927 1855 3993
rect 226 3893 297 3927
rect 226 3723 260 3773
rect 1821 3723 1855 3789
rect 226 3689 297 3723
rect 226 3519 260 3569
rect 1821 3519 1855 3585
rect 226 3485 297 3519
rect 226 3315 260 3365
rect 1821 3315 1855 3381
rect 226 3281 297 3315
rect 226 3111 260 3161
rect 1821 3111 1855 3177
rect 226 3077 297 3111
rect 226 2907 260 2957
rect 1821 2907 1855 2973
rect 226 2873 297 2907
rect 226 2703 260 2753
rect 1821 2703 1855 2769
rect 226 2669 297 2703
rect 226 2499 260 2549
rect 1821 2499 1855 2565
rect 226 2465 297 2499
rect 226 2295 260 2345
rect 1821 2295 1855 2361
rect 226 2261 297 2295
rect 226 2091 260 2141
rect 1821 2091 1855 2157
rect 226 2057 297 2091
rect 226 1887 260 1937
rect 1821 1887 1855 1953
rect 226 1853 297 1887
rect 226 1683 260 1733
rect 1821 1683 1855 1749
rect 226 1649 297 1683
rect 226 1479 260 1529
rect 1821 1479 1855 1545
rect 226 1445 297 1479
rect 226 1275 260 1325
rect 1821 1275 1855 1341
rect 226 1241 297 1275
rect 226 1071 260 1121
rect 1821 1071 1855 1137
rect 226 1037 297 1071
rect 226 867 260 917
rect 1821 867 1855 933
rect 226 833 297 867
rect 226 663 260 713
rect 1821 663 1855 729
rect 226 629 297 663
rect 226 459 260 509
rect 1821 459 1855 525
rect 226 425 297 459
rect 226 255 260 305
rect 1821 255 1855 321
rect 226 221 297 255
rect 226 51 260 101
rect 1821 51 1855 117
rect 226 17 297 51
<< metal1 >>
rect 316 -14 344 9806
rect 1232 -14 1260 9806
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_0
timestamp 1581321264
transform 1 0 0 0 1 9588
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_1
timestamp 1581321264
transform 1 0 0 0 1 9384
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_2
timestamp 1581321264
transform 1 0 0 0 1 9180
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_3
timestamp 1581321264
transform 1 0 0 0 1 8976
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_4
timestamp 1581321264
transform 1 0 0 0 1 8772
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_5
timestamp 1581321264
transform 1 0 0 0 1 8568
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_6
timestamp 1581321264
transform 1 0 0 0 1 8364
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_7
timestamp 1581321264
transform 1 0 0 0 1 8160
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_8
timestamp 1581321264
transform 1 0 0 0 1 7956
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_9
timestamp 1581321264
transform 1 0 0 0 1 7752
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_10
timestamp 1581321264
transform 1 0 0 0 1 7548
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_11
timestamp 1581321264
transform 1 0 0 0 1 7344
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_12
timestamp 1581321264
transform 1 0 0 0 1 7140
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_13
timestamp 1581321264
transform 1 0 0 0 1 6936
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_14
timestamp 1581321264
transform 1 0 0 0 1 6732
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_15
timestamp 1581321264
transform 1 0 0 0 1 6528
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_16
timestamp 1581321264
transform 1 0 0 0 1 6324
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_17
timestamp 1581321264
transform 1 0 0 0 1 6120
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_18
timestamp 1581321264
transform 1 0 0 0 1 5916
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_19
timestamp 1581321264
transform 1 0 0 0 1 5712
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_20
timestamp 1581321264
transform 1 0 0 0 1 5508
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_21
timestamp 1581321264
transform 1 0 0 0 1 5304
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_22
timestamp 1581321264
transform 1 0 0 0 1 5100
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_23
timestamp 1581321264
transform 1 0 0 0 1 4896
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_24
timestamp 1581321264
transform 1 0 0 0 1 4692
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_25
timestamp 1581321264
transform 1 0 0 0 1 4488
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_26
timestamp 1581321264
transform 1 0 0 0 1 4284
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_27
timestamp 1581321264
transform 1 0 0 0 1 4080
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_28
timestamp 1581321264
transform 1 0 0 0 1 3876
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_29
timestamp 1581321264
transform 1 0 0 0 1 3672
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_30
timestamp 1581321264
transform 1 0 0 0 1 3468
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_31
timestamp 1581321264
transform 1 0 0 0 1 3264
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_32
timestamp 1581321264
transform 1 0 0 0 1 3060
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_33
timestamp 1581321264
transform 1 0 0 0 1 2856
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_34
timestamp 1581321264
transform 1 0 0 0 1 2652
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_35
timestamp 1581321264
transform 1 0 0 0 1 2448
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_36
timestamp 1581321264
transform 1 0 0 0 1 2244
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_37
timestamp 1581321264
transform 1 0 0 0 1 2040
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_38
timestamp 1581321264
transform 1 0 0 0 1 1836
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_39
timestamp 1581321264
transform 1 0 0 0 1 1632
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_40
timestamp 1581321264
transform 1 0 0 0 1 1428
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_41
timestamp 1581321264
transform 1 0 0 0 1 1224
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_42
timestamp 1581321264
transform 1 0 0 0 1 1020
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_43
timestamp 1581321264
transform 1 0 0 0 1 816
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_44
timestamp 1581321264
transform 1 0 0 0 1 612
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_45
timestamp 1581321264
transform 1 0 0 0 1 408
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_46
timestamp 1581321264
transform 1 0 0 0 1 204
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_47
timestamp 1581321264
transform 1 0 0 0 1 0
box 136 -79 1879 299
<< labels >>
rlabel locali s 1838 9672 1838 9672 4 in_0
port 2 nsew
rlabel locali s 243 9672 243 9672 4 out_0
port 3 nsew
rlabel locali s 1838 9468 1838 9468 4 in_1
port 4 nsew
rlabel locali s 243 9468 243 9468 4 out_1
port 5 nsew
rlabel locali s 1838 9264 1838 9264 4 in_2
port 6 nsew
rlabel locali s 243 9264 243 9264 4 out_2
port 7 nsew
rlabel locali s 1838 9060 1838 9060 4 in_3
port 8 nsew
rlabel locali s 243 9060 243 9060 4 out_3
port 9 nsew
rlabel locali s 1838 8856 1838 8856 4 in_4
port 10 nsew
rlabel locali s 243 8856 243 8856 4 out_4
port 11 nsew
rlabel locali s 1838 8652 1838 8652 4 in_5
port 12 nsew
rlabel locali s 243 8652 243 8652 4 out_5
port 13 nsew
rlabel locali s 1838 8448 1838 8448 4 in_6
port 14 nsew
rlabel locali s 243 8448 243 8448 4 out_6
port 15 nsew
rlabel locali s 1838 8244 1838 8244 4 in_7
port 16 nsew
rlabel locali s 243 8244 243 8244 4 out_7
port 17 nsew
rlabel locali s 1838 8040 1838 8040 4 in_8
port 18 nsew
rlabel locali s 243 8040 243 8040 4 out_8
port 19 nsew
rlabel locali s 1838 7836 1838 7836 4 in_9
port 20 nsew
rlabel locali s 243 7836 243 7836 4 out_9
port 21 nsew
rlabel locali s 1838 7632 1838 7632 4 in_10
port 22 nsew
rlabel locali s 243 7632 243 7632 4 out_10
port 23 nsew
rlabel locali s 1838 7428 1838 7428 4 in_11
port 24 nsew
rlabel locali s 243 7428 243 7428 4 out_11
port 25 nsew
rlabel locali s 1838 7224 1838 7224 4 in_12
port 26 nsew
rlabel locali s 243 7224 243 7224 4 out_12
port 27 nsew
rlabel locali s 1838 7020 1838 7020 4 in_13
port 28 nsew
rlabel locali s 243 7020 243 7020 4 out_13
port 29 nsew
rlabel locali s 1838 6816 1838 6816 4 in_14
port 30 nsew
rlabel locali s 243 6816 243 6816 4 out_14
port 31 nsew
rlabel locali s 1838 6612 1838 6612 4 in_15
port 32 nsew
rlabel locali s 243 6612 243 6612 4 out_15
port 33 nsew
rlabel locali s 1838 6408 1838 6408 4 in_16
port 34 nsew
rlabel locali s 243 6408 243 6408 4 out_16
port 35 nsew
rlabel locali s 1838 6204 1838 6204 4 in_17
port 36 nsew
rlabel locali s 243 6204 243 6204 4 out_17
port 37 nsew
rlabel locali s 1838 6000 1838 6000 4 in_18
port 38 nsew
rlabel locali s 243 6000 243 6000 4 out_18
port 39 nsew
rlabel locali s 1838 5796 1838 5796 4 in_19
port 40 nsew
rlabel locali s 243 5796 243 5796 4 out_19
port 41 nsew
rlabel locali s 1838 5592 1838 5592 4 in_20
port 42 nsew
rlabel locali s 243 5592 243 5592 4 out_20
port 43 nsew
rlabel locali s 1838 5388 1838 5388 4 in_21
port 44 nsew
rlabel locali s 243 5388 243 5388 4 out_21
port 45 nsew
rlabel locali s 1838 5184 1838 5184 4 in_22
port 46 nsew
rlabel locali s 243 5184 243 5184 4 out_22
port 47 nsew
rlabel locali s 1838 4980 1838 4980 4 in_23
port 48 nsew
rlabel locali s 243 4980 243 4980 4 out_23
port 49 nsew
rlabel locali s 1838 4776 1838 4776 4 in_24
port 50 nsew
rlabel locali s 243 4776 243 4776 4 out_24
port 51 nsew
rlabel locali s 1838 4572 1838 4572 4 in_25
port 52 nsew
rlabel locali s 243 4572 243 4572 4 out_25
port 53 nsew
rlabel locali s 1838 4368 1838 4368 4 in_26
port 54 nsew
rlabel locali s 243 4368 243 4368 4 out_26
port 55 nsew
rlabel locali s 1838 4164 1838 4164 4 in_27
port 56 nsew
rlabel locali s 243 4164 243 4164 4 out_27
port 57 nsew
rlabel locali s 1838 3960 1838 3960 4 in_28
port 58 nsew
rlabel locali s 243 3960 243 3960 4 out_28
port 59 nsew
rlabel locali s 1838 3756 1838 3756 4 in_29
port 60 nsew
rlabel locali s 243 3756 243 3756 4 out_29
port 61 nsew
rlabel locali s 1838 3552 1838 3552 4 in_30
port 62 nsew
rlabel locali s 243 3552 243 3552 4 out_30
port 63 nsew
rlabel locali s 1838 3348 1838 3348 4 in_31
port 64 nsew
rlabel locali s 243 3348 243 3348 4 out_31
port 65 nsew
rlabel locali s 1838 3144 1838 3144 4 in_32
port 66 nsew
rlabel locali s 243 3144 243 3144 4 out_32
port 67 nsew
rlabel locali s 1838 2940 1838 2940 4 in_33
port 68 nsew
rlabel locali s 243 2940 243 2940 4 out_33
port 69 nsew
rlabel locali s 1838 2736 1838 2736 4 in_34
port 70 nsew
rlabel locali s 243 2736 243 2736 4 out_34
port 71 nsew
rlabel locali s 1838 2532 1838 2532 4 in_35
port 72 nsew
rlabel locali s 243 2532 243 2532 4 out_35
port 73 nsew
rlabel locali s 1838 2328 1838 2328 4 in_36
port 74 nsew
rlabel locali s 243 2328 243 2328 4 out_36
port 75 nsew
rlabel locali s 1838 2124 1838 2124 4 in_37
port 76 nsew
rlabel locali s 243 2124 243 2124 4 out_37
port 77 nsew
rlabel locali s 1838 1920 1838 1920 4 in_38
port 78 nsew
rlabel locali s 243 1920 243 1920 4 out_38
port 79 nsew
rlabel locali s 1838 1716 1838 1716 4 in_39
port 80 nsew
rlabel locali s 243 1716 243 1716 4 out_39
port 81 nsew
rlabel locali s 1838 1512 1838 1512 4 in_40
port 82 nsew
rlabel locali s 243 1512 243 1512 4 out_40
port 83 nsew
rlabel locali s 1838 1308 1838 1308 4 in_41
port 84 nsew
rlabel locali s 243 1308 243 1308 4 out_41
port 85 nsew
rlabel locali s 1838 1104 1838 1104 4 in_42
port 86 nsew
rlabel locali s 243 1104 243 1104 4 out_42
port 87 nsew
rlabel locali s 1838 900 1838 900 4 in_43
port 88 nsew
rlabel locali s 243 900 243 900 4 out_43
port 89 nsew
rlabel locali s 1838 696 1838 696 4 in_44
port 90 nsew
rlabel locali s 243 696 243 696 4 out_44
port 91 nsew
rlabel locali s 1838 492 1838 492 4 in_45
port 92 nsew
rlabel locali s 243 492 243 492 4 out_45
port 93 nsew
rlabel locali s 1838 288 1838 288 4 in_46
port 94 nsew
rlabel locali s 243 288 243 288 4 out_46
port 95 nsew
rlabel locali s 1838 84 1838 84 4 in_47
port 96 nsew
rlabel locali s 243 84 243 84 4 out_47
port 97 nsew
rlabel metal1 s 316 -14 344 14 4 gnd
port 99 nsew
rlabel metal1 s 316 9778 344 9806 4 gnd
port 99 nsew
rlabel metal1 s 1232 9778 1260 9806 4 vdd
port 101 nsew
rlabel metal1 s 1232 -14 1260 14 4 vdd
port 101 nsew
<< properties >>
string FIXED_BBOX 0 0 1782 9792
<< end >>
