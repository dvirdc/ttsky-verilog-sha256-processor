magic
tech sky130A
magscale 1 2
timestamp 1581320207
<< checkpaint >>
rect -1299 -1216 8035 11725
<< locali >>
rect 3177 10091 3211 10107
rect 6723 10057 6757 10091
rect 3177 10041 3211 10057
rect 3177 9887 3211 9903
rect 6723 9853 6757 9887
rect 3177 9837 3211 9853
rect 3177 9683 3211 9699
rect 6723 9649 6757 9683
rect 3177 9633 3211 9649
rect 3177 9479 3211 9495
rect 6723 9445 6757 9479
rect 3177 9429 3211 9445
rect 3177 9275 3211 9291
rect 6723 9241 6757 9275
rect 3177 9225 3211 9241
rect 3177 9071 3211 9087
rect 6723 9037 6757 9071
rect 3177 9021 3211 9037
rect 3177 8867 3211 8883
rect 6723 8833 6757 8867
rect 3177 8817 3211 8833
rect 3177 8663 3211 8679
rect 6723 8629 6757 8663
rect 3177 8613 3211 8629
rect 3177 8355 3211 8371
rect 6723 8321 6757 8355
rect 3177 8305 3211 8321
rect 3177 8151 3211 8167
rect 6723 8117 6757 8151
rect 3177 8101 3211 8117
rect 3177 7947 3211 7963
rect 6723 7913 6757 7947
rect 3177 7897 3211 7913
rect 3177 7743 3211 7759
rect 6723 7709 6757 7743
rect 3177 7693 3211 7709
rect 3177 7539 3211 7555
rect 6723 7505 6757 7539
rect 3177 7489 3211 7505
rect 3177 7335 3211 7351
rect 6723 7301 6757 7335
rect 3177 7285 3211 7301
rect 3177 7131 3211 7147
rect 6723 7097 6757 7131
rect 3177 7081 3211 7097
rect 3177 6927 3211 6943
rect 6723 6893 6757 6927
rect 3177 6877 3211 6893
rect 3177 6619 3211 6635
rect 6723 6585 6757 6619
rect 3177 6569 3211 6585
rect 3177 6415 3211 6431
rect 6723 6381 6757 6415
rect 3177 6365 3211 6381
rect 3177 6211 3211 6227
rect 6723 6177 6757 6211
rect 3177 6161 3211 6177
rect 3177 6007 3211 6023
rect 6723 5973 6757 6007
rect 3177 5957 3211 5973
rect 3177 5803 3211 5819
rect 6723 5769 6757 5803
rect 3177 5753 3211 5769
rect 3177 5599 3211 5615
rect 6723 5565 6757 5599
rect 3177 5549 3211 5565
rect 3177 5395 3211 5411
rect 6723 5361 6757 5395
rect 3177 5345 3211 5361
rect 3177 5191 3211 5207
rect 6723 5157 6757 5191
rect 3177 5141 3211 5157
rect 3177 4883 3211 4899
rect 6723 4849 6757 4883
rect 3177 4833 3211 4849
rect 3177 4679 3211 4695
rect 6723 4645 6757 4679
rect 3177 4629 3211 4645
rect 3177 4475 3211 4491
rect 6723 4441 6757 4475
rect 3177 4425 3211 4441
rect 3177 4271 3211 4287
rect 6723 4237 6757 4271
rect 3177 4221 3211 4237
rect 3177 4067 3211 4083
rect 6723 4033 6757 4067
rect 3177 4017 3211 4033
rect 3177 3863 3211 3879
rect 6723 3829 6757 3863
rect 3177 3813 3211 3829
rect 3177 3659 3211 3675
rect 6723 3625 6757 3659
rect 3177 3609 3211 3625
rect 3177 3455 3211 3471
rect 6723 3421 6757 3455
rect 3177 3405 3211 3421
rect 321 60 387 94
rect 729 60 795 94
rect 1137 60 1203 94
rect 1545 60 1611 94
rect 1953 60 2019 94
<< viali >>
rect 3177 10057 3211 10091
rect 3177 9853 3211 9887
rect 3177 9649 3211 9683
rect 3177 9445 3211 9479
rect 3177 9241 3211 9275
rect 3177 9037 3211 9071
rect 3177 8833 3211 8867
rect 3177 8629 3211 8663
rect 3177 8321 3211 8355
rect 3177 8117 3211 8151
rect 3177 7913 3211 7947
rect 3177 7709 3211 7743
rect 3177 7505 3211 7539
rect 3177 7301 3211 7335
rect 3177 7097 3211 7131
rect 3177 6893 3211 6927
rect 3177 6585 3211 6619
rect 3177 6381 3211 6415
rect 3177 6177 3211 6211
rect 3177 5973 3211 6007
rect 3177 5769 3211 5803
rect 3177 5565 3211 5599
rect 3177 5361 3211 5395
rect 3177 5157 3211 5191
rect 3177 4849 3211 4883
rect 3177 4645 3211 4679
rect 3177 4441 3211 4475
rect 3177 4237 3211 4271
rect 3177 4033 3211 4067
rect 3177 3829 3211 3863
rect 3177 3625 3211 3659
rect 3177 3421 3211 3455
<< metal1 >>
rect 2693 10437 2721 10465
rect 3339 10180 3367 10208
rect 3961 10180 3989 10208
rect 4759 10180 4787 10208
rect 6007 10180 6035 10208
rect 3165 10091 3223 10097
rect 3165 10088 3177 10091
rect 3075 10060 3177 10088
rect 3165 10057 3177 10060
rect 3211 10057 3223 10091
rect 3165 10051 3223 10057
rect 3165 9887 3223 9893
rect 3165 9884 3177 9887
rect 3075 9856 3177 9884
rect 3165 9853 3177 9856
rect 3211 9853 3223 9887
rect 3165 9847 3223 9853
rect 3165 9683 3223 9689
rect 3165 9680 3177 9683
rect 3075 9652 3177 9680
rect 3165 9649 3177 9652
rect 3211 9649 3223 9683
rect 3165 9643 3223 9649
rect 3165 9479 3223 9485
rect 3165 9476 3177 9479
rect 3075 9448 3177 9476
rect 3165 9445 3177 9448
rect 3211 9445 3223 9479
rect 3165 9439 3223 9445
rect 3165 9275 3223 9281
rect 3165 9272 3177 9275
rect 3075 9244 3177 9272
rect 3165 9241 3177 9244
rect 3211 9241 3223 9275
rect 3165 9235 3223 9241
rect 3165 9071 3223 9077
rect 3165 9068 3177 9071
rect 3075 9040 3177 9068
rect 3165 9037 3177 9040
rect 3211 9037 3223 9071
rect 3165 9031 3223 9037
rect 3165 8867 3223 8873
rect 3165 8864 3177 8867
rect 3075 8836 3177 8864
rect 3165 8833 3177 8836
rect 3211 8833 3223 8867
rect 3165 8827 3223 8833
rect 3165 8663 3223 8669
rect 3165 8660 3177 8663
rect 3075 8632 3177 8660
rect 3165 8629 3177 8632
rect 3211 8629 3223 8663
rect 3165 8623 3223 8629
rect 3165 8355 3223 8361
rect 3165 8352 3177 8355
rect 3075 8324 3177 8352
rect 3165 8321 3177 8324
rect 3211 8321 3223 8355
rect 3165 8315 3223 8321
rect 3165 8151 3223 8157
rect 3165 8148 3177 8151
rect 3075 8120 3177 8148
rect 3165 8117 3177 8120
rect 3211 8117 3223 8151
rect 3165 8111 3223 8117
rect 3165 7947 3223 7953
rect 3165 7944 3177 7947
rect 3075 7916 3177 7944
rect 3165 7913 3177 7916
rect 3211 7913 3223 7947
rect 3165 7907 3223 7913
rect 3165 7743 3223 7749
rect 3165 7740 3177 7743
rect 3075 7712 3177 7740
rect 3165 7709 3177 7712
rect 3211 7709 3223 7743
rect 3165 7703 3223 7709
rect 3165 7539 3223 7545
rect 3165 7536 3177 7539
rect 3075 7508 3177 7536
rect 3165 7505 3177 7508
rect 3211 7505 3223 7539
rect 3165 7499 3223 7505
rect 3165 7335 3223 7341
rect 3165 7332 3177 7335
rect 3075 7304 3177 7332
rect 3165 7301 3177 7304
rect 3211 7301 3223 7335
rect 3165 7295 3223 7301
rect 3165 7131 3223 7137
rect 3165 7128 3177 7131
rect 3075 7100 3177 7128
rect 3165 7097 3177 7100
rect 3211 7097 3223 7131
rect 3165 7091 3223 7097
rect 3165 6927 3223 6933
rect 3165 6924 3177 6927
rect 3075 6896 3177 6924
rect 3165 6893 3177 6896
rect 3211 6893 3223 6927
rect 3165 6887 3223 6893
rect 3165 6619 3223 6625
rect 3165 6616 3177 6619
rect 3075 6588 3177 6616
rect 3165 6585 3177 6588
rect 3211 6585 3223 6619
rect 3165 6579 3223 6585
rect 3165 6415 3223 6421
rect 3165 6412 3177 6415
rect 3075 6384 3177 6412
rect 3165 6381 3177 6384
rect 3211 6381 3223 6415
rect 3165 6375 3223 6381
rect 3165 6211 3223 6217
rect 3165 6208 3177 6211
rect 3075 6180 3177 6208
rect 3165 6177 3177 6180
rect 3211 6177 3223 6211
rect 3165 6171 3223 6177
rect 3165 6007 3223 6013
rect 3165 6004 3177 6007
rect 3075 5976 3177 6004
rect 3165 5973 3177 5976
rect 3211 5973 3223 6007
rect 3165 5967 3223 5973
rect 3165 5803 3223 5809
rect 3165 5800 3177 5803
rect 3075 5772 3177 5800
rect 3165 5769 3177 5772
rect 3211 5769 3223 5803
rect 3165 5763 3223 5769
rect 3165 5599 3223 5605
rect 3165 5596 3177 5599
rect 3075 5568 3177 5596
rect 3165 5565 3177 5568
rect 3211 5565 3223 5599
rect 3165 5559 3223 5565
rect 3165 5395 3223 5401
rect 3165 5392 3177 5395
rect 3075 5364 3177 5392
rect 3165 5361 3177 5364
rect 3211 5361 3223 5395
rect 3165 5355 3223 5361
rect 3165 5191 3223 5197
rect 3165 5188 3177 5191
rect 3075 5160 3177 5188
rect 3165 5157 3177 5160
rect 3211 5157 3223 5191
rect 3165 5151 3223 5157
rect 3165 4883 3223 4889
rect 3165 4880 3177 4883
rect 3075 4852 3177 4880
rect 3165 4849 3177 4852
rect 3211 4849 3223 4883
rect 3165 4843 3223 4849
rect 3165 4679 3223 4685
rect 3165 4676 3177 4679
rect 3075 4648 3177 4676
rect 3165 4645 3177 4648
rect 3211 4645 3223 4679
rect 3165 4639 3223 4645
rect 3165 4475 3223 4481
rect 3165 4472 3177 4475
rect 3075 4444 3177 4472
rect 3165 4441 3177 4444
rect 3211 4441 3223 4475
rect 3165 4435 3223 4441
rect 3165 4271 3223 4277
rect 3165 4268 3177 4271
rect 3075 4240 3177 4268
rect 3165 4237 3177 4240
rect 3211 4237 3223 4271
rect 3165 4231 3223 4237
rect 3165 4067 3223 4073
rect 3165 4064 3177 4067
rect 3075 4036 3177 4064
rect 3165 4033 3177 4036
rect 3211 4033 3223 4067
rect 3165 4027 3223 4033
rect 3165 3863 3223 3869
rect 3165 3860 3177 3863
rect 3075 3832 3177 3860
rect 3165 3829 3177 3832
rect 3211 3829 3223 3863
rect 3165 3823 3223 3829
rect 3165 3659 3223 3665
rect 3165 3656 3177 3659
rect 3075 3628 3177 3656
rect 3165 3625 3177 3628
rect 3211 3625 3223 3659
rect 3165 3619 3223 3625
rect 3165 3455 3223 3461
rect 3165 3452 3177 3455
rect 3075 3424 3177 3452
rect 3165 3421 3177 3424
rect 3211 3421 3223 3455
rect 3165 3415 3223 3421
rect 3339 3256 3367 3284
rect 3961 3256 3989 3284
rect 4759 3256 4787 3284
rect 6007 3256 6035 3284
rect 298 3199 304 3251
rect 356 3199 362 3251
rect 502 3199 508 3251
rect 560 3199 566 3251
rect 706 3199 712 3251
rect 764 3199 770 3251
rect 910 3199 916 3251
rect 968 3199 974 3251
rect 1114 3199 1120 3251
rect 1172 3199 1178 3251
rect 1318 3199 1324 3251
rect 1376 3199 1382 3251
rect 1522 3199 1528 3251
rect 1580 3199 1586 3251
rect 1726 3199 1732 3251
rect 1784 3199 1790 3251
rect 1930 3199 1936 3251
rect 1988 3199 1994 3251
rect 2134 3199 2140 3251
rect 2192 3199 2198 3251
rect 316 3138 344 3199
rect 298 3086 304 3138
rect 356 3086 362 3138
rect 438 3086 444 3138
rect 496 3126 502 3138
rect 520 3126 548 3199
rect 724 3138 752 3199
rect 496 3098 548 3126
rect 496 3086 502 3098
rect 706 3086 712 3138
rect 764 3086 770 3138
rect 846 3086 852 3138
rect 904 3126 910 3138
rect 928 3126 956 3199
rect 1132 3138 1160 3199
rect 904 3098 956 3126
rect 904 3086 910 3098
rect 1114 3086 1120 3138
rect 1172 3086 1178 3138
rect 1254 3086 1260 3138
rect 1312 3126 1318 3138
rect 1336 3126 1364 3199
rect 1540 3138 1568 3199
rect 1312 3098 1364 3126
rect 1312 3086 1318 3098
rect 1522 3086 1528 3138
rect 1580 3086 1586 3138
rect 1662 3086 1668 3138
rect 1720 3126 1726 3138
rect 1744 3126 1772 3199
rect 1948 3138 1976 3199
rect 1720 3098 1772 3126
rect 1720 3086 1726 3098
rect 1930 3086 1936 3138
rect 1988 3086 1994 3138
rect 2070 3086 2076 3138
rect 2128 3126 2134 3138
rect 2152 3126 2180 3199
rect 2128 3098 2180 3126
rect 2128 3086 2134 3098
rect 127 2833 155 2861
rect 2167 2408 2195 2436
rect 127 2160 2167 2188
rect 127 1881 155 1909
rect 2167 1456 2195 1484
rect 127 844 155 872
rect 2167 222 2195 250
<< via1 >>
rect 304 3199 356 3251
rect 508 3199 560 3251
rect 712 3199 764 3251
rect 916 3199 968 3251
rect 1120 3199 1172 3251
rect 1324 3199 1376 3251
rect 1528 3199 1580 3251
rect 1732 3199 1784 3251
rect 1936 3199 1988 3251
rect 2140 3199 2192 3251
rect 304 3086 356 3138
rect 444 3086 496 3138
rect 712 3086 764 3138
rect 852 3086 904 3138
rect 1120 3086 1172 3138
rect 1260 3086 1312 3138
rect 1528 3086 1580 3138
rect 1668 3086 1720 3138
rect 1936 3086 1988 3138
rect 2076 3086 2128 3138
<< metal2 >>
rect 304 3251 356 3257
rect 304 3193 356 3199
rect 508 3251 560 3257
rect 508 3193 560 3199
rect 712 3251 764 3257
rect 712 3193 764 3199
rect 916 3251 968 3257
rect 916 3193 968 3199
rect 1120 3251 1172 3257
rect 1120 3193 1172 3199
rect 1324 3251 1376 3257
rect 1324 3193 1376 3199
rect 1528 3251 1580 3257
rect 1528 3193 1580 3199
rect 1732 3251 1784 3257
rect 1732 3193 1784 3199
rect 1936 3251 1988 3257
rect 1936 3193 1988 3199
rect 2140 3251 2192 3257
rect 2693 3253 2721 3281
rect 3057 3204 3121 3232
rect 2140 3193 2192 3199
rect 304 3138 356 3144
rect 304 3080 356 3086
rect 444 3138 496 3144
rect 444 3080 496 3086
rect 712 3138 764 3144
rect 712 3080 764 3086
rect 852 3138 904 3144
rect 852 3080 904 3086
rect 1120 3138 1172 3144
rect 1120 3080 1172 3086
rect 1260 3138 1312 3144
rect 1260 3080 1312 3086
rect 1528 3138 1580 3144
rect 1528 3080 1580 3086
rect 1668 3138 1720 3144
rect 1668 3080 1720 3086
rect 1936 3138 1988 3144
rect 1936 3080 1988 3086
rect 2076 3138 2128 3144
rect 2076 3080 2128 3086
<< metal3 >>
rect -31 10167 29 10227
rect 2051 10167 2111 10227
rect -31 8431 29 8491
rect 2051 8431 2111 8491
rect -31 6695 29 6755
rect 2051 6695 2111 6755
rect -31 4959 29 5019
rect 2051 4959 2111 5019
rect -31 3223 29 3283
rect 2051 3223 2111 3283
use sky130_rom_krom_rom_address_control_array  sky130_rom_krom_rom_address_control_array_0
timestamp 1581320207
transform 1 0 127 0 1 0
box -48 44 2135 3128
use sky130_rom_krom_rom_row_decode_array  sky130_rom_krom_rom_row_decode_array_0
timestamp 1581320207
transform 0 -1 3089 1 0 3192
box -6 -84 7273 3128
use sky130_rom_krom_rom_row_decode_wordline_buffer  sky130_rom_krom_rom_row_decode_wordline_buffer_0
timestamp 1581320207
transform 1 0 3117 0 1 3250
box 44 -50 3658 7039
<< labels >>
rlabel metal1 s 127 2160 2167 2188 4 clk
port 3 nsew
rlabel locali s 6740 3438 6740 3438 4 wl_0
port 4 nsew
rlabel locali s 6740 3642 6740 3642 4 wl_1
port 5 nsew
rlabel locali s 6740 3846 6740 3846 4 wl_2
port 6 nsew
rlabel locali s 6740 4050 6740 4050 4 wl_3
port 7 nsew
rlabel locali s 6740 4254 6740 4254 4 wl_4
port 8 nsew
rlabel locali s 6740 4458 6740 4458 4 wl_5
port 9 nsew
rlabel locali s 6740 4662 6740 4662 4 wl_6
port 10 nsew
rlabel locali s 6740 4866 6740 4866 4 wl_7
port 11 nsew
rlabel locali s 6740 5174 6740 5174 4 wl_8
port 12 nsew
rlabel locali s 6740 5378 6740 5378 4 wl_9
port 13 nsew
rlabel locali s 6740 5582 6740 5582 4 wl_10
port 14 nsew
rlabel locali s 6740 5786 6740 5786 4 wl_11
port 15 nsew
rlabel locali s 6740 5990 6740 5990 4 wl_12
port 16 nsew
rlabel locali s 6740 6194 6740 6194 4 wl_13
port 17 nsew
rlabel locali s 6740 6398 6740 6398 4 wl_14
port 18 nsew
rlabel locali s 6740 6602 6740 6602 4 wl_15
port 19 nsew
rlabel locali s 6740 6910 6740 6910 4 wl_16
port 20 nsew
rlabel locali s 6740 7114 6740 7114 4 wl_17
port 21 nsew
rlabel locali s 6740 7318 6740 7318 4 wl_18
port 22 nsew
rlabel locali s 6740 7522 6740 7522 4 wl_19
port 23 nsew
rlabel locali s 6740 7726 6740 7726 4 wl_20
port 24 nsew
rlabel locali s 6740 7930 6740 7930 4 wl_21
port 25 nsew
rlabel locali s 6740 8134 6740 8134 4 wl_22
port 26 nsew
rlabel locali s 6740 8338 6740 8338 4 wl_23
port 27 nsew
rlabel locali s 6740 8646 6740 8646 4 wl_24
port 28 nsew
rlabel locali s 6740 8850 6740 8850 4 wl_25
port 29 nsew
rlabel locali s 6740 9054 6740 9054 4 wl_26
port 30 nsew
rlabel locali s 6740 9258 6740 9258 4 wl_27
port 31 nsew
rlabel locali s 6740 9462 6740 9462 4 wl_28
port 32 nsew
rlabel locali s 6740 9666 6740 9666 4 wl_29
port 33 nsew
rlabel locali s 6740 9870 6740 9870 4 wl_30
port 34 nsew
rlabel locali s 6740 10074 6740 10074 4 wl_31
port 35 nsew
rlabel metal2 s 2693 3253 2721 3281 4 precharge
port 37 nsew
rlabel metal1 s 2693 10437 2721 10465 4 precharge_r
port 39 nsew
rlabel locali s 354 77 354 77 4 A0
port 40 nsew
rlabel locali s 762 77 762 77 4 A1
port 41 nsew
rlabel locali s 1170 77 1170 77 4 A2
port 42 nsew
rlabel locali s 1578 77 1578 77 4 A3
port 43 nsew
rlabel locali s 1986 77 1986 77 4 A4
port 44 nsew
rlabel metal1 s 3961 10180 3989 10208 4 vdd
port 46 nsew
rlabel metal1 s 3961 3256 3989 3284 4 vdd
port 46 nsew
rlabel metal1 s 127 844 155 872 4 vdd
port 46 nsew
rlabel metal1 s 127 1881 155 1909 4 vdd
port 46 nsew
rlabel metal1 s 6007 3256 6035 3284 4 vdd
port 46 nsew
rlabel metal1 s 127 2833 155 2861 4 vdd
port 46 nsew
rlabel metal1 s 6007 10180 6035 10208 4 vdd
port 46 nsew
rlabel metal2 s 3057 3204 3121 3232 4 vdd
port 46 nsew
rlabel metal3 s 2051 3223 2111 3283 4 gnd
port 48 nsew
rlabel metal1 s 3339 10180 3367 10208 4 gnd
port 48 nsew
rlabel metal3 s -31 3223 29 3283 4 gnd
port 48 nsew
rlabel metal1 s 2167 2408 2195 2436 4 gnd
port 48 nsew
rlabel metal3 s 2051 8431 2111 8491 4 gnd
port 48 nsew
rlabel metal1 s 2167 222 2195 250 4 gnd
port 48 nsew
rlabel metal3 s 2051 6695 2111 6755 4 gnd
port 48 nsew
rlabel metal3 s -31 6695 29 6755 4 gnd
port 48 nsew
rlabel metal3 s -31 4959 29 5019 4 gnd
port 48 nsew
rlabel metal1 s 3339 3256 3367 3284 4 gnd
port 48 nsew
rlabel metal3 s 2051 10167 2111 10227 4 gnd
port 48 nsew
rlabel metal3 s -31 10167 29 10227 4 gnd
port 48 nsew
rlabel metal1 s 4759 3256 4787 3284 4 gnd
port 48 nsew
rlabel metal1 s 2167 1456 2195 1484 4 gnd
port 48 nsew
rlabel metal1 s 4759 10180 4787 10208 4 gnd
port 48 nsew
rlabel metal3 s -31 8431 29 8491 4 gnd
port 48 nsew
rlabel metal3 s 2051 4959 2111 5019 4 gnd
port 48 nsew
<< properties >>
string FIXED_BBOX -31 0 6757 10465
<< end >>
