magic
tech sky130A
magscale 1 2
timestamp 1581449086
<< checkpaint >>
rect -1260 -1344 53733 4073
<< pwell >>
rect 177 822 52345 924
<< psubdiff >>
rect 203 890 285 898
rect 203 856 227 890
rect 261 856 285 890
rect 203 848 285 856
rect 407 890 489 898
rect 407 856 431 890
rect 465 856 489 890
rect 407 848 489 856
rect 611 890 693 898
rect 611 856 635 890
rect 669 856 693 890
rect 611 848 693 856
rect 815 890 897 898
rect 815 856 839 890
rect 873 856 897 890
rect 815 848 897 856
rect 1019 890 1101 898
rect 1019 856 1043 890
rect 1077 856 1101 890
rect 1019 848 1101 856
rect 1223 890 1305 898
rect 1223 856 1247 890
rect 1281 856 1305 890
rect 1223 848 1305 856
rect 1427 890 1509 898
rect 1427 856 1451 890
rect 1485 856 1509 890
rect 1427 848 1509 856
rect 1631 890 1713 898
rect 1631 856 1655 890
rect 1689 856 1713 890
rect 1631 848 1713 856
rect 1835 890 1917 898
rect 1835 856 1859 890
rect 1893 856 1917 890
rect 1835 848 1917 856
rect 2039 890 2121 898
rect 2039 856 2063 890
rect 2097 856 2121 890
rect 2039 848 2121 856
rect 2243 890 2325 898
rect 2243 856 2267 890
rect 2301 856 2325 890
rect 2243 848 2325 856
rect 2447 890 2529 898
rect 2447 856 2471 890
rect 2505 856 2529 890
rect 2447 848 2529 856
rect 2651 890 2733 898
rect 2651 856 2675 890
rect 2709 856 2733 890
rect 2651 848 2733 856
rect 2855 890 2937 898
rect 2855 856 2879 890
rect 2913 856 2937 890
rect 2855 848 2937 856
rect 3059 890 3141 898
rect 3059 856 3083 890
rect 3117 856 3141 890
rect 3059 848 3141 856
rect 3263 890 3345 898
rect 3263 856 3287 890
rect 3321 856 3345 890
rect 3263 848 3345 856
rect 3467 890 3549 898
rect 3467 856 3491 890
rect 3525 856 3549 890
rect 3467 848 3549 856
rect 3671 890 3753 898
rect 3671 856 3695 890
rect 3729 856 3753 890
rect 3671 848 3753 856
rect 3875 890 3957 898
rect 3875 856 3899 890
rect 3933 856 3957 890
rect 3875 848 3957 856
rect 4079 890 4161 898
rect 4079 856 4103 890
rect 4137 856 4161 890
rect 4079 848 4161 856
rect 4283 890 4365 898
rect 4283 856 4307 890
rect 4341 856 4365 890
rect 4283 848 4365 856
rect 4487 890 4569 898
rect 4487 856 4511 890
rect 4545 856 4569 890
rect 4487 848 4569 856
rect 4691 890 4773 898
rect 4691 856 4715 890
rect 4749 856 4773 890
rect 4691 848 4773 856
rect 4895 890 4977 898
rect 4895 856 4919 890
rect 4953 856 4977 890
rect 4895 848 4977 856
rect 5099 890 5181 898
rect 5099 856 5123 890
rect 5157 856 5181 890
rect 5099 848 5181 856
rect 5303 890 5385 898
rect 5303 856 5327 890
rect 5361 856 5385 890
rect 5303 848 5385 856
rect 5507 890 5589 898
rect 5507 856 5531 890
rect 5565 856 5589 890
rect 5507 848 5589 856
rect 5711 890 5793 898
rect 5711 856 5735 890
rect 5769 856 5793 890
rect 5711 848 5793 856
rect 5915 890 5997 898
rect 5915 856 5939 890
rect 5973 856 5997 890
rect 5915 848 5997 856
rect 6119 890 6201 898
rect 6119 856 6143 890
rect 6177 856 6201 890
rect 6119 848 6201 856
rect 6323 890 6405 898
rect 6323 856 6347 890
rect 6381 856 6405 890
rect 6323 848 6405 856
rect 6527 890 6609 898
rect 6527 856 6551 890
rect 6585 856 6609 890
rect 6527 848 6609 856
rect 6731 890 6813 898
rect 6731 856 6755 890
rect 6789 856 6813 890
rect 6731 848 6813 856
rect 6935 890 7017 898
rect 6935 856 6959 890
rect 6993 856 7017 890
rect 6935 848 7017 856
rect 7139 890 7221 898
rect 7139 856 7163 890
rect 7197 856 7221 890
rect 7139 848 7221 856
rect 7343 890 7425 898
rect 7343 856 7367 890
rect 7401 856 7425 890
rect 7343 848 7425 856
rect 7547 890 7629 898
rect 7547 856 7571 890
rect 7605 856 7629 890
rect 7547 848 7629 856
rect 7751 890 7833 898
rect 7751 856 7775 890
rect 7809 856 7833 890
rect 7751 848 7833 856
rect 7955 890 8037 898
rect 7955 856 7979 890
rect 8013 856 8037 890
rect 7955 848 8037 856
rect 8159 890 8241 898
rect 8159 856 8183 890
rect 8217 856 8241 890
rect 8159 848 8241 856
rect 8363 890 8445 898
rect 8363 856 8387 890
rect 8421 856 8445 890
rect 8363 848 8445 856
rect 8567 890 8649 898
rect 8567 856 8591 890
rect 8625 856 8649 890
rect 8567 848 8649 856
rect 8771 890 8853 898
rect 8771 856 8795 890
rect 8829 856 8853 890
rect 8771 848 8853 856
rect 8975 890 9057 898
rect 8975 856 8999 890
rect 9033 856 9057 890
rect 8975 848 9057 856
rect 9179 890 9261 898
rect 9179 856 9203 890
rect 9237 856 9261 890
rect 9179 848 9261 856
rect 9383 890 9465 898
rect 9383 856 9407 890
rect 9441 856 9465 890
rect 9383 848 9465 856
rect 9587 890 9669 898
rect 9587 856 9611 890
rect 9645 856 9669 890
rect 9587 848 9669 856
rect 9791 890 9873 898
rect 9791 856 9815 890
rect 9849 856 9873 890
rect 9791 848 9873 856
rect 9995 890 10077 898
rect 9995 856 10019 890
rect 10053 856 10077 890
rect 9995 848 10077 856
rect 10199 890 10281 898
rect 10199 856 10223 890
rect 10257 856 10281 890
rect 10199 848 10281 856
rect 10403 890 10485 898
rect 10403 856 10427 890
rect 10461 856 10485 890
rect 10403 848 10485 856
rect 10607 890 10689 898
rect 10607 856 10631 890
rect 10665 856 10689 890
rect 10607 848 10689 856
rect 10811 890 10893 898
rect 10811 856 10835 890
rect 10869 856 10893 890
rect 10811 848 10893 856
rect 11015 890 11097 898
rect 11015 856 11039 890
rect 11073 856 11097 890
rect 11015 848 11097 856
rect 11219 890 11301 898
rect 11219 856 11243 890
rect 11277 856 11301 890
rect 11219 848 11301 856
rect 11423 890 11505 898
rect 11423 856 11447 890
rect 11481 856 11505 890
rect 11423 848 11505 856
rect 11627 890 11709 898
rect 11627 856 11651 890
rect 11685 856 11709 890
rect 11627 848 11709 856
rect 11831 890 11913 898
rect 11831 856 11855 890
rect 11889 856 11913 890
rect 11831 848 11913 856
rect 12035 890 12117 898
rect 12035 856 12059 890
rect 12093 856 12117 890
rect 12035 848 12117 856
rect 12239 890 12321 898
rect 12239 856 12263 890
rect 12297 856 12321 890
rect 12239 848 12321 856
rect 12443 890 12525 898
rect 12443 856 12467 890
rect 12501 856 12525 890
rect 12443 848 12525 856
rect 12647 890 12729 898
rect 12647 856 12671 890
rect 12705 856 12729 890
rect 12647 848 12729 856
rect 12851 890 12933 898
rect 12851 856 12875 890
rect 12909 856 12933 890
rect 12851 848 12933 856
rect 13055 890 13137 898
rect 13055 856 13079 890
rect 13113 856 13137 890
rect 13055 848 13137 856
rect 13259 890 13341 898
rect 13259 856 13283 890
rect 13317 856 13341 890
rect 13259 848 13341 856
rect 13463 890 13545 898
rect 13463 856 13487 890
rect 13521 856 13545 890
rect 13463 848 13545 856
rect 13667 890 13749 898
rect 13667 856 13691 890
rect 13725 856 13749 890
rect 13667 848 13749 856
rect 13871 890 13953 898
rect 13871 856 13895 890
rect 13929 856 13953 890
rect 13871 848 13953 856
rect 14075 890 14157 898
rect 14075 856 14099 890
rect 14133 856 14157 890
rect 14075 848 14157 856
rect 14279 890 14361 898
rect 14279 856 14303 890
rect 14337 856 14361 890
rect 14279 848 14361 856
rect 14483 890 14565 898
rect 14483 856 14507 890
rect 14541 856 14565 890
rect 14483 848 14565 856
rect 14687 890 14769 898
rect 14687 856 14711 890
rect 14745 856 14769 890
rect 14687 848 14769 856
rect 14891 890 14973 898
rect 14891 856 14915 890
rect 14949 856 14973 890
rect 14891 848 14973 856
rect 15095 890 15177 898
rect 15095 856 15119 890
rect 15153 856 15177 890
rect 15095 848 15177 856
rect 15299 890 15381 898
rect 15299 856 15323 890
rect 15357 856 15381 890
rect 15299 848 15381 856
rect 15503 890 15585 898
rect 15503 856 15527 890
rect 15561 856 15585 890
rect 15503 848 15585 856
rect 15707 890 15789 898
rect 15707 856 15731 890
rect 15765 856 15789 890
rect 15707 848 15789 856
rect 15911 890 15993 898
rect 15911 856 15935 890
rect 15969 856 15993 890
rect 15911 848 15993 856
rect 16115 890 16197 898
rect 16115 856 16139 890
rect 16173 856 16197 890
rect 16115 848 16197 856
rect 16319 890 16401 898
rect 16319 856 16343 890
rect 16377 856 16401 890
rect 16319 848 16401 856
rect 16523 890 16605 898
rect 16523 856 16547 890
rect 16581 856 16605 890
rect 16523 848 16605 856
rect 16727 890 16809 898
rect 16727 856 16751 890
rect 16785 856 16809 890
rect 16727 848 16809 856
rect 16931 890 17013 898
rect 16931 856 16955 890
rect 16989 856 17013 890
rect 16931 848 17013 856
rect 17135 890 17217 898
rect 17135 856 17159 890
rect 17193 856 17217 890
rect 17135 848 17217 856
rect 17339 890 17421 898
rect 17339 856 17363 890
rect 17397 856 17421 890
rect 17339 848 17421 856
rect 17543 890 17625 898
rect 17543 856 17567 890
rect 17601 856 17625 890
rect 17543 848 17625 856
rect 17747 890 17829 898
rect 17747 856 17771 890
rect 17805 856 17829 890
rect 17747 848 17829 856
rect 17951 890 18033 898
rect 17951 856 17975 890
rect 18009 856 18033 890
rect 17951 848 18033 856
rect 18155 890 18237 898
rect 18155 856 18179 890
rect 18213 856 18237 890
rect 18155 848 18237 856
rect 18359 890 18441 898
rect 18359 856 18383 890
rect 18417 856 18441 890
rect 18359 848 18441 856
rect 18563 890 18645 898
rect 18563 856 18587 890
rect 18621 856 18645 890
rect 18563 848 18645 856
rect 18767 890 18849 898
rect 18767 856 18791 890
rect 18825 856 18849 890
rect 18767 848 18849 856
rect 18971 890 19053 898
rect 18971 856 18995 890
rect 19029 856 19053 890
rect 18971 848 19053 856
rect 19175 890 19257 898
rect 19175 856 19199 890
rect 19233 856 19257 890
rect 19175 848 19257 856
rect 19379 890 19461 898
rect 19379 856 19403 890
rect 19437 856 19461 890
rect 19379 848 19461 856
rect 19583 890 19665 898
rect 19583 856 19607 890
rect 19641 856 19665 890
rect 19583 848 19665 856
rect 19787 890 19869 898
rect 19787 856 19811 890
rect 19845 856 19869 890
rect 19787 848 19869 856
rect 19991 890 20073 898
rect 19991 856 20015 890
rect 20049 856 20073 890
rect 19991 848 20073 856
rect 20195 890 20277 898
rect 20195 856 20219 890
rect 20253 856 20277 890
rect 20195 848 20277 856
rect 20399 890 20481 898
rect 20399 856 20423 890
rect 20457 856 20481 890
rect 20399 848 20481 856
rect 20603 890 20685 898
rect 20603 856 20627 890
rect 20661 856 20685 890
rect 20603 848 20685 856
rect 20807 890 20889 898
rect 20807 856 20831 890
rect 20865 856 20889 890
rect 20807 848 20889 856
rect 21011 890 21093 898
rect 21011 856 21035 890
rect 21069 856 21093 890
rect 21011 848 21093 856
rect 21215 890 21297 898
rect 21215 856 21239 890
rect 21273 856 21297 890
rect 21215 848 21297 856
rect 21419 890 21501 898
rect 21419 856 21443 890
rect 21477 856 21501 890
rect 21419 848 21501 856
rect 21623 890 21705 898
rect 21623 856 21647 890
rect 21681 856 21705 890
rect 21623 848 21705 856
rect 21827 890 21909 898
rect 21827 856 21851 890
rect 21885 856 21909 890
rect 21827 848 21909 856
rect 22031 890 22113 898
rect 22031 856 22055 890
rect 22089 856 22113 890
rect 22031 848 22113 856
rect 22235 890 22317 898
rect 22235 856 22259 890
rect 22293 856 22317 890
rect 22235 848 22317 856
rect 22439 890 22521 898
rect 22439 856 22463 890
rect 22497 856 22521 890
rect 22439 848 22521 856
rect 22643 890 22725 898
rect 22643 856 22667 890
rect 22701 856 22725 890
rect 22643 848 22725 856
rect 22847 890 22929 898
rect 22847 856 22871 890
rect 22905 856 22929 890
rect 22847 848 22929 856
rect 23051 890 23133 898
rect 23051 856 23075 890
rect 23109 856 23133 890
rect 23051 848 23133 856
rect 23255 890 23337 898
rect 23255 856 23279 890
rect 23313 856 23337 890
rect 23255 848 23337 856
rect 23459 890 23541 898
rect 23459 856 23483 890
rect 23517 856 23541 890
rect 23459 848 23541 856
rect 23663 890 23745 898
rect 23663 856 23687 890
rect 23721 856 23745 890
rect 23663 848 23745 856
rect 23867 890 23949 898
rect 23867 856 23891 890
rect 23925 856 23949 890
rect 23867 848 23949 856
rect 24071 890 24153 898
rect 24071 856 24095 890
rect 24129 856 24153 890
rect 24071 848 24153 856
rect 24275 890 24357 898
rect 24275 856 24299 890
rect 24333 856 24357 890
rect 24275 848 24357 856
rect 24479 890 24561 898
rect 24479 856 24503 890
rect 24537 856 24561 890
rect 24479 848 24561 856
rect 24683 890 24765 898
rect 24683 856 24707 890
rect 24741 856 24765 890
rect 24683 848 24765 856
rect 24887 890 24969 898
rect 24887 856 24911 890
rect 24945 856 24969 890
rect 24887 848 24969 856
rect 25091 890 25173 898
rect 25091 856 25115 890
rect 25149 856 25173 890
rect 25091 848 25173 856
rect 25295 890 25377 898
rect 25295 856 25319 890
rect 25353 856 25377 890
rect 25295 848 25377 856
rect 25499 890 25581 898
rect 25499 856 25523 890
rect 25557 856 25581 890
rect 25499 848 25581 856
rect 25703 890 25785 898
rect 25703 856 25727 890
rect 25761 856 25785 890
rect 25703 848 25785 856
rect 25907 890 25989 898
rect 25907 856 25931 890
rect 25965 856 25989 890
rect 25907 848 25989 856
rect 26111 890 26193 898
rect 26111 856 26135 890
rect 26169 856 26193 890
rect 26111 848 26193 856
rect 26315 890 26397 898
rect 26315 856 26339 890
rect 26373 856 26397 890
rect 26315 848 26397 856
rect 26519 890 26601 898
rect 26519 856 26543 890
rect 26577 856 26601 890
rect 26519 848 26601 856
rect 26723 890 26805 898
rect 26723 856 26747 890
rect 26781 856 26805 890
rect 26723 848 26805 856
rect 26927 890 27009 898
rect 26927 856 26951 890
rect 26985 856 27009 890
rect 26927 848 27009 856
rect 27131 890 27213 898
rect 27131 856 27155 890
rect 27189 856 27213 890
rect 27131 848 27213 856
rect 27335 890 27417 898
rect 27335 856 27359 890
rect 27393 856 27417 890
rect 27335 848 27417 856
rect 27539 890 27621 898
rect 27539 856 27563 890
rect 27597 856 27621 890
rect 27539 848 27621 856
rect 27743 890 27825 898
rect 27743 856 27767 890
rect 27801 856 27825 890
rect 27743 848 27825 856
rect 27947 890 28029 898
rect 27947 856 27971 890
rect 28005 856 28029 890
rect 27947 848 28029 856
rect 28151 890 28233 898
rect 28151 856 28175 890
rect 28209 856 28233 890
rect 28151 848 28233 856
rect 28355 890 28437 898
rect 28355 856 28379 890
rect 28413 856 28437 890
rect 28355 848 28437 856
rect 28559 890 28641 898
rect 28559 856 28583 890
rect 28617 856 28641 890
rect 28559 848 28641 856
rect 28763 890 28845 898
rect 28763 856 28787 890
rect 28821 856 28845 890
rect 28763 848 28845 856
rect 28967 890 29049 898
rect 28967 856 28991 890
rect 29025 856 29049 890
rect 28967 848 29049 856
rect 29171 890 29253 898
rect 29171 856 29195 890
rect 29229 856 29253 890
rect 29171 848 29253 856
rect 29375 890 29457 898
rect 29375 856 29399 890
rect 29433 856 29457 890
rect 29375 848 29457 856
rect 29579 890 29661 898
rect 29579 856 29603 890
rect 29637 856 29661 890
rect 29579 848 29661 856
rect 29783 890 29865 898
rect 29783 856 29807 890
rect 29841 856 29865 890
rect 29783 848 29865 856
rect 29987 890 30069 898
rect 29987 856 30011 890
rect 30045 856 30069 890
rect 29987 848 30069 856
rect 30191 890 30273 898
rect 30191 856 30215 890
rect 30249 856 30273 890
rect 30191 848 30273 856
rect 30395 890 30477 898
rect 30395 856 30419 890
rect 30453 856 30477 890
rect 30395 848 30477 856
rect 30599 890 30681 898
rect 30599 856 30623 890
rect 30657 856 30681 890
rect 30599 848 30681 856
rect 30803 890 30885 898
rect 30803 856 30827 890
rect 30861 856 30885 890
rect 30803 848 30885 856
rect 31007 890 31089 898
rect 31007 856 31031 890
rect 31065 856 31089 890
rect 31007 848 31089 856
rect 31211 890 31293 898
rect 31211 856 31235 890
rect 31269 856 31293 890
rect 31211 848 31293 856
rect 31415 890 31497 898
rect 31415 856 31439 890
rect 31473 856 31497 890
rect 31415 848 31497 856
rect 31619 890 31701 898
rect 31619 856 31643 890
rect 31677 856 31701 890
rect 31619 848 31701 856
rect 31823 890 31905 898
rect 31823 856 31847 890
rect 31881 856 31905 890
rect 31823 848 31905 856
rect 32027 890 32109 898
rect 32027 856 32051 890
rect 32085 856 32109 890
rect 32027 848 32109 856
rect 32231 890 32313 898
rect 32231 856 32255 890
rect 32289 856 32313 890
rect 32231 848 32313 856
rect 32435 890 32517 898
rect 32435 856 32459 890
rect 32493 856 32517 890
rect 32435 848 32517 856
rect 32639 890 32721 898
rect 32639 856 32663 890
rect 32697 856 32721 890
rect 32639 848 32721 856
rect 32843 890 32925 898
rect 32843 856 32867 890
rect 32901 856 32925 890
rect 32843 848 32925 856
rect 33047 890 33129 898
rect 33047 856 33071 890
rect 33105 856 33129 890
rect 33047 848 33129 856
rect 33251 890 33333 898
rect 33251 856 33275 890
rect 33309 856 33333 890
rect 33251 848 33333 856
rect 33455 890 33537 898
rect 33455 856 33479 890
rect 33513 856 33537 890
rect 33455 848 33537 856
rect 33659 890 33741 898
rect 33659 856 33683 890
rect 33717 856 33741 890
rect 33659 848 33741 856
rect 33863 890 33945 898
rect 33863 856 33887 890
rect 33921 856 33945 890
rect 33863 848 33945 856
rect 34067 890 34149 898
rect 34067 856 34091 890
rect 34125 856 34149 890
rect 34067 848 34149 856
rect 34271 890 34353 898
rect 34271 856 34295 890
rect 34329 856 34353 890
rect 34271 848 34353 856
rect 34475 890 34557 898
rect 34475 856 34499 890
rect 34533 856 34557 890
rect 34475 848 34557 856
rect 34679 890 34761 898
rect 34679 856 34703 890
rect 34737 856 34761 890
rect 34679 848 34761 856
rect 34883 890 34965 898
rect 34883 856 34907 890
rect 34941 856 34965 890
rect 34883 848 34965 856
rect 35087 890 35169 898
rect 35087 856 35111 890
rect 35145 856 35169 890
rect 35087 848 35169 856
rect 35291 890 35373 898
rect 35291 856 35315 890
rect 35349 856 35373 890
rect 35291 848 35373 856
rect 35495 890 35577 898
rect 35495 856 35519 890
rect 35553 856 35577 890
rect 35495 848 35577 856
rect 35699 890 35781 898
rect 35699 856 35723 890
rect 35757 856 35781 890
rect 35699 848 35781 856
rect 35903 890 35985 898
rect 35903 856 35927 890
rect 35961 856 35985 890
rect 35903 848 35985 856
rect 36107 890 36189 898
rect 36107 856 36131 890
rect 36165 856 36189 890
rect 36107 848 36189 856
rect 36311 890 36393 898
rect 36311 856 36335 890
rect 36369 856 36393 890
rect 36311 848 36393 856
rect 36515 890 36597 898
rect 36515 856 36539 890
rect 36573 856 36597 890
rect 36515 848 36597 856
rect 36719 890 36801 898
rect 36719 856 36743 890
rect 36777 856 36801 890
rect 36719 848 36801 856
rect 36923 890 37005 898
rect 36923 856 36947 890
rect 36981 856 37005 890
rect 36923 848 37005 856
rect 37127 890 37209 898
rect 37127 856 37151 890
rect 37185 856 37209 890
rect 37127 848 37209 856
rect 37331 890 37413 898
rect 37331 856 37355 890
rect 37389 856 37413 890
rect 37331 848 37413 856
rect 37535 890 37617 898
rect 37535 856 37559 890
rect 37593 856 37617 890
rect 37535 848 37617 856
rect 37739 890 37821 898
rect 37739 856 37763 890
rect 37797 856 37821 890
rect 37739 848 37821 856
rect 37943 890 38025 898
rect 37943 856 37967 890
rect 38001 856 38025 890
rect 37943 848 38025 856
rect 38147 890 38229 898
rect 38147 856 38171 890
rect 38205 856 38229 890
rect 38147 848 38229 856
rect 38351 890 38433 898
rect 38351 856 38375 890
rect 38409 856 38433 890
rect 38351 848 38433 856
rect 38555 890 38637 898
rect 38555 856 38579 890
rect 38613 856 38637 890
rect 38555 848 38637 856
rect 38759 890 38841 898
rect 38759 856 38783 890
rect 38817 856 38841 890
rect 38759 848 38841 856
rect 38963 890 39045 898
rect 38963 856 38987 890
rect 39021 856 39045 890
rect 38963 848 39045 856
rect 39167 890 39249 898
rect 39167 856 39191 890
rect 39225 856 39249 890
rect 39167 848 39249 856
rect 39371 890 39453 898
rect 39371 856 39395 890
rect 39429 856 39453 890
rect 39371 848 39453 856
rect 39575 890 39657 898
rect 39575 856 39599 890
rect 39633 856 39657 890
rect 39575 848 39657 856
rect 39779 890 39861 898
rect 39779 856 39803 890
rect 39837 856 39861 890
rect 39779 848 39861 856
rect 39983 890 40065 898
rect 39983 856 40007 890
rect 40041 856 40065 890
rect 39983 848 40065 856
rect 40187 890 40269 898
rect 40187 856 40211 890
rect 40245 856 40269 890
rect 40187 848 40269 856
rect 40391 890 40473 898
rect 40391 856 40415 890
rect 40449 856 40473 890
rect 40391 848 40473 856
rect 40595 890 40677 898
rect 40595 856 40619 890
rect 40653 856 40677 890
rect 40595 848 40677 856
rect 40799 890 40881 898
rect 40799 856 40823 890
rect 40857 856 40881 890
rect 40799 848 40881 856
rect 41003 890 41085 898
rect 41003 856 41027 890
rect 41061 856 41085 890
rect 41003 848 41085 856
rect 41207 890 41289 898
rect 41207 856 41231 890
rect 41265 856 41289 890
rect 41207 848 41289 856
rect 41411 890 41493 898
rect 41411 856 41435 890
rect 41469 856 41493 890
rect 41411 848 41493 856
rect 41615 890 41697 898
rect 41615 856 41639 890
rect 41673 856 41697 890
rect 41615 848 41697 856
rect 41819 890 41901 898
rect 41819 856 41843 890
rect 41877 856 41901 890
rect 41819 848 41901 856
rect 42023 890 42105 898
rect 42023 856 42047 890
rect 42081 856 42105 890
rect 42023 848 42105 856
rect 42227 890 42309 898
rect 42227 856 42251 890
rect 42285 856 42309 890
rect 42227 848 42309 856
rect 42431 890 42513 898
rect 42431 856 42455 890
rect 42489 856 42513 890
rect 42431 848 42513 856
rect 42635 890 42717 898
rect 42635 856 42659 890
rect 42693 856 42717 890
rect 42635 848 42717 856
rect 42839 890 42921 898
rect 42839 856 42863 890
rect 42897 856 42921 890
rect 42839 848 42921 856
rect 43043 890 43125 898
rect 43043 856 43067 890
rect 43101 856 43125 890
rect 43043 848 43125 856
rect 43247 890 43329 898
rect 43247 856 43271 890
rect 43305 856 43329 890
rect 43247 848 43329 856
rect 43451 890 43533 898
rect 43451 856 43475 890
rect 43509 856 43533 890
rect 43451 848 43533 856
rect 43655 890 43737 898
rect 43655 856 43679 890
rect 43713 856 43737 890
rect 43655 848 43737 856
rect 43859 890 43941 898
rect 43859 856 43883 890
rect 43917 856 43941 890
rect 43859 848 43941 856
rect 44063 890 44145 898
rect 44063 856 44087 890
rect 44121 856 44145 890
rect 44063 848 44145 856
rect 44267 890 44349 898
rect 44267 856 44291 890
rect 44325 856 44349 890
rect 44267 848 44349 856
rect 44471 890 44553 898
rect 44471 856 44495 890
rect 44529 856 44553 890
rect 44471 848 44553 856
rect 44675 890 44757 898
rect 44675 856 44699 890
rect 44733 856 44757 890
rect 44675 848 44757 856
rect 44879 890 44961 898
rect 44879 856 44903 890
rect 44937 856 44961 890
rect 44879 848 44961 856
rect 45083 890 45165 898
rect 45083 856 45107 890
rect 45141 856 45165 890
rect 45083 848 45165 856
rect 45287 890 45369 898
rect 45287 856 45311 890
rect 45345 856 45369 890
rect 45287 848 45369 856
rect 45491 890 45573 898
rect 45491 856 45515 890
rect 45549 856 45573 890
rect 45491 848 45573 856
rect 45695 890 45777 898
rect 45695 856 45719 890
rect 45753 856 45777 890
rect 45695 848 45777 856
rect 45899 890 45981 898
rect 45899 856 45923 890
rect 45957 856 45981 890
rect 45899 848 45981 856
rect 46103 890 46185 898
rect 46103 856 46127 890
rect 46161 856 46185 890
rect 46103 848 46185 856
rect 46307 890 46389 898
rect 46307 856 46331 890
rect 46365 856 46389 890
rect 46307 848 46389 856
rect 46511 890 46593 898
rect 46511 856 46535 890
rect 46569 856 46593 890
rect 46511 848 46593 856
rect 46715 890 46797 898
rect 46715 856 46739 890
rect 46773 856 46797 890
rect 46715 848 46797 856
rect 46919 890 47001 898
rect 46919 856 46943 890
rect 46977 856 47001 890
rect 46919 848 47001 856
rect 47123 890 47205 898
rect 47123 856 47147 890
rect 47181 856 47205 890
rect 47123 848 47205 856
rect 47327 890 47409 898
rect 47327 856 47351 890
rect 47385 856 47409 890
rect 47327 848 47409 856
rect 47531 890 47613 898
rect 47531 856 47555 890
rect 47589 856 47613 890
rect 47531 848 47613 856
rect 47735 890 47817 898
rect 47735 856 47759 890
rect 47793 856 47817 890
rect 47735 848 47817 856
rect 47939 890 48021 898
rect 47939 856 47963 890
rect 47997 856 48021 890
rect 47939 848 48021 856
rect 48143 890 48225 898
rect 48143 856 48167 890
rect 48201 856 48225 890
rect 48143 848 48225 856
rect 48347 890 48429 898
rect 48347 856 48371 890
rect 48405 856 48429 890
rect 48347 848 48429 856
rect 48551 890 48633 898
rect 48551 856 48575 890
rect 48609 856 48633 890
rect 48551 848 48633 856
rect 48755 890 48837 898
rect 48755 856 48779 890
rect 48813 856 48837 890
rect 48755 848 48837 856
rect 48959 890 49041 898
rect 48959 856 48983 890
rect 49017 856 49041 890
rect 48959 848 49041 856
rect 49163 890 49245 898
rect 49163 856 49187 890
rect 49221 856 49245 890
rect 49163 848 49245 856
rect 49367 890 49449 898
rect 49367 856 49391 890
rect 49425 856 49449 890
rect 49367 848 49449 856
rect 49571 890 49653 898
rect 49571 856 49595 890
rect 49629 856 49653 890
rect 49571 848 49653 856
rect 49775 890 49857 898
rect 49775 856 49799 890
rect 49833 856 49857 890
rect 49775 848 49857 856
rect 49979 890 50061 898
rect 49979 856 50003 890
rect 50037 856 50061 890
rect 49979 848 50061 856
rect 50183 890 50265 898
rect 50183 856 50207 890
rect 50241 856 50265 890
rect 50183 848 50265 856
rect 50387 890 50469 898
rect 50387 856 50411 890
rect 50445 856 50469 890
rect 50387 848 50469 856
rect 50591 890 50673 898
rect 50591 856 50615 890
rect 50649 856 50673 890
rect 50591 848 50673 856
rect 50795 890 50877 898
rect 50795 856 50819 890
rect 50853 856 50877 890
rect 50795 848 50877 856
rect 50999 890 51081 898
rect 50999 856 51023 890
rect 51057 856 51081 890
rect 50999 848 51081 856
rect 51203 890 51285 898
rect 51203 856 51227 890
rect 51261 856 51285 890
rect 51203 848 51285 856
rect 51407 890 51489 898
rect 51407 856 51431 890
rect 51465 856 51489 890
rect 51407 848 51489 856
rect 51611 890 51693 898
rect 51611 856 51635 890
rect 51669 856 51693 890
rect 51611 848 51693 856
rect 51815 890 51897 898
rect 51815 856 51839 890
rect 51873 856 51897 890
rect 51815 848 51897 856
rect 52019 890 52101 898
rect 52019 856 52043 890
rect 52077 856 52101 890
rect 52019 848 52101 856
rect 52237 890 52319 898
rect 52237 856 52261 890
rect 52295 856 52319 890
rect 52237 848 52319 856
<< psubdiffcont >>
rect 227 856 261 890
rect 431 856 465 890
rect 635 856 669 890
rect 839 856 873 890
rect 1043 856 1077 890
rect 1247 856 1281 890
rect 1451 856 1485 890
rect 1655 856 1689 890
rect 1859 856 1893 890
rect 2063 856 2097 890
rect 2267 856 2301 890
rect 2471 856 2505 890
rect 2675 856 2709 890
rect 2879 856 2913 890
rect 3083 856 3117 890
rect 3287 856 3321 890
rect 3491 856 3525 890
rect 3695 856 3729 890
rect 3899 856 3933 890
rect 4103 856 4137 890
rect 4307 856 4341 890
rect 4511 856 4545 890
rect 4715 856 4749 890
rect 4919 856 4953 890
rect 5123 856 5157 890
rect 5327 856 5361 890
rect 5531 856 5565 890
rect 5735 856 5769 890
rect 5939 856 5973 890
rect 6143 856 6177 890
rect 6347 856 6381 890
rect 6551 856 6585 890
rect 6755 856 6789 890
rect 6959 856 6993 890
rect 7163 856 7197 890
rect 7367 856 7401 890
rect 7571 856 7605 890
rect 7775 856 7809 890
rect 7979 856 8013 890
rect 8183 856 8217 890
rect 8387 856 8421 890
rect 8591 856 8625 890
rect 8795 856 8829 890
rect 8999 856 9033 890
rect 9203 856 9237 890
rect 9407 856 9441 890
rect 9611 856 9645 890
rect 9815 856 9849 890
rect 10019 856 10053 890
rect 10223 856 10257 890
rect 10427 856 10461 890
rect 10631 856 10665 890
rect 10835 856 10869 890
rect 11039 856 11073 890
rect 11243 856 11277 890
rect 11447 856 11481 890
rect 11651 856 11685 890
rect 11855 856 11889 890
rect 12059 856 12093 890
rect 12263 856 12297 890
rect 12467 856 12501 890
rect 12671 856 12705 890
rect 12875 856 12909 890
rect 13079 856 13113 890
rect 13283 856 13317 890
rect 13487 856 13521 890
rect 13691 856 13725 890
rect 13895 856 13929 890
rect 14099 856 14133 890
rect 14303 856 14337 890
rect 14507 856 14541 890
rect 14711 856 14745 890
rect 14915 856 14949 890
rect 15119 856 15153 890
rect 15323 856 15357 890
rect 15527 856 15561 890
rect 15731 856 15765 890
rect 15935 856 15969 890
rect 16139 856 16173 890
rect 16343 856 16377 890
rect 16547 856 16581 890
rect 16751 856 16785 890
rect 16955 856 16989 890
rect 17159 856 17193 890
rect 17363 856 17397 890
rect 17567 856 17601 890
rect 17771 856 17805 890
rect 17975 856 18009 890
rect 18179 856 18213 890
rect 18383 856 18417 890
rect 18587 856 18621 890
rect 18791 856 18825 890
rect 18995 856 19029 890
rect 19199 856 19233 890
rect 19403 856 19437 890
rect 19607 856 19641 890
rect 19811 856 19845 890
rect 20015 856 20049 890
rect 20219 856 20253 890
rect 20423 856 20457 890
rect 20627 856 20661 890
rect 20831 856 20865 890
rect 21035 856 21069 890
rect 21239 856 21273 890
rect 21443 856 21477 890
rect 21647 856 21681 890
rect 21851 856 21885 890
rect 22055 856 22089 890
rect 22259 856 22293 890
rect 22463 856 22497 890
rect 22667 856 22701 890
rect 22871 856 22905 890
rect 23075 856 23109 890
rect 23279 856 23313 890
rect 23483 856 23517 890
rect 23687 856 23721 890
rect 23891 856 23925 890
rect 24095 856 24129 890
rect 24299 856 24333 890
rect 24503 856 24537 890
rect 24707 856 24741 890
rect 24911 856 24945 890
rect 25115 856 25149 890
rect 25319 856 25353 890
rect 25523 856 25557 890
rect 25727 856 25761 890
rect 25931 856 25965 890
rect 26135 856 26169 890
rect 26339 856 26373 890
rect 26543 856 26577 890
rect 26747 856 26781 890
rect 26951 856 26985 890
rect 27155 856 27189 890
rect 27359 856 27393 890
rect 27563 856 27597 890
rect 27767 856 27801 890
rect 27971 856 28005 890
rect 28175 856 28209 890
rect 28379 856 28413 890
rect 28583 856 28617 890
rect 28787 856 28821 890
rect 28991 856 29025 890
rect 29195 856 29229 890
rect 29399 856 29433 890
rect 29603 856 29637 890
rect 29807 856 29841 890
rect 30011 856 30045 890
rect 30215 856 30249 890
rect 30419 856 30453 890
rect 30623 856 30657 890
rect 30827 856 30861 890
rect 31031 856 31065 890
rect 31235 856 31269 890
rect 31439 856 31473 890
rect 31643 856 31677 890
rect 31847 856 31881 890
rect 32051 856 32085 890
rect 32255 856 32289 890
rect 32459 856 32493 890
rect 32663 856 32697 890
rect 32867 856 32901 890
rect 33071 856 33105 890
rect 33275 856 33309 890
rect 33479 856 33513 890
rect 33683 856 33717 890
rect 33887 856 33921 890
rect 34091 856 34125 890
rect 34295 856 34329 890
rect 34499 856 34533 890
rect 34703 856 34737 890
rect 34907 856 34941 890
rect 35111 856 35145 890
rect 35315 856 35349 890
rect 35519 856 35553 890
rect 35723 856 35757 890
rect 35927 856 35961 890
rect 36131 856 36165 890
rect 36335 856 36369 890
rect 36539 856 36573 890
rect 36743 856 36777 890
rect 36947 856 36981 890
rect 37151 856 37185 890
rect 37355 856 37389 890
rect 37559 856 37593 890
rect 37763 856 37797 890
rect 37967 856 38001 890
rect 38171 856 38205 890
rect 38375 856 38409 890
rect 38579 856 38613 890
rect 38783 856 38817 890
rect 38987 856 39021 890
rect 39191 856 39225 890
rect 39395 856 39429 890
rect 39599 856 39633 890
rect 39803 856 39837 890
rect 40007 856 40041 890
rect 40211 856 40245 890
rect 40415 856 40449 890
rect 40619 856 40653 890
rect 40823 856 40857 890
rect 41027 856 41061 890
rect 41231 856 41265 890
rect 41435 856 41469 890
rect 41639 856 41673 890
rect 41843 856 41877 890
rect 42047 856 42081 890
rect 42251 856 42285 890
rect 42455 856 42489 890
rect 42659 856 42693 890
rect 42863 856 42897 890
rect 43067 856 43101 890
rect 43271 856 43305 890
rect 43475 856 43509 890
rect 43679 856 43713 890
rect 43883 856 43917 890
rect 44087 856 44121 890
rect 44291 856 44325 890
rect 44495 856 44529 890
rect 44699 856 44733 890
rect 44903 856 44937 890
rect 45107 856 45141 890
rect 45311 856 45345 890
rect 45515 856 45549 890
rect 45719 856 45753 890
rect 45923 856 45957 890
rect 46127 856 46161 890
rect 46331 856 46365 890
rect 46535 856 46569 890
rect 46739 856 46773 890
rect 46943 856 46977 890
rect 47147 856 47181 890
rect 47351 856 47385 890
rect 47555 856 47589 890
rect 47759 856 47793 890
rect 47963 856 47997 890
rect 48167 856 48201 890
rect 48371 856 48405 890
rect 48575 856 48609 890
rect 48779 856 48813 890
rect 48983 856 49017 890
rect 49187 856 49221 890
rect 49391 856 49425 890
rect 49595 856 49629 890
rect 49799 856 49833 890
rect 50003 856 50037 890
rect 50207 856 50241 890
rect 50411 856 50445 890
rect 50615 856 50649 890
rect 50819 856 50853 890
rect 51023 856 51057 890
rect 51227 856 51261 890
rect 51431 856 51465 890
rect 51635 856 51669 890
rect 51839 856 51873 890
rect 52043 856 52077 890
rect 52261 856 52295 890
<< poly >>
rect 0 2676 66 2692
rect 0 2642 16 2676
rect 50 2674 66 2676
rect 1632 2676 1698 2692
rect 1632 2674 1648 2676
rect 50 2644 1648 2674
rect 50 2642 66 2644
rect 0 2626 66 2642
rect 1632 2642 1648 2644
rect 1682 2674 1698 2676
rect 3264 2676 3330 2692
rect 3264 2674 3280 2676
rect 1682 2644 3280 2674
rect 1682 2642 1698 2644
rect 1632 2626 1698 2642
rect 3264 2642 3280 2644
rect 3314 2674 3330 2676
rect 4896 2676 4962 2692
rect 4896 2674 4912 2676
rect 3314 2644 4912 2674
rect 3314 2642 3330 2644
rect 3264 2626 3330 2642
rect 4896 2642 4912 2644
rect 4946 2674 4962 2676
rect 6528 2676 6594 2692
rect 6528 2674 6544 2676
rect 4946 2644 6544 2674
rect 4946 2642 4962 2644
rect 4896 2626 4962 2642
rect 6528 2642 6544 2644
rect 6578 2674 6594 2676
rect 8160 2676 8226 2692
rect 8160 2674 8176 2676
rect 6578 2644 8176 2674
rect 6578 2642 6594 2644
rect 6528 2626 6594 2642
rect 8160 2642 8176 2644
rect 8210 2674 8226 2676
rect 9792 2676 9858 2692
rect 9792 2674 9808 2676
rect 8210 2644 9808 2674
rect 8210 2642 8226 2644
rect 8160 2626 8226 2642
rect 9792 2642 9808 2644
rect 9842 2674 9858 2676
rect 11424 2676 11490 2692
rect 11424 2674 11440 2676
rect 9842 2644 11440 2674
rect 9842 2642 9858 2644
rect 9792 2626 9858 2642
rect 11424 2642 11440 2644
rect 11474 2674 11490 2676
rect 13056 2676 13122 2692
rect 13056 2674 13072 2676
rect 11474 2644 13072 2674
rect 11474 2642 11490 2644
rect 11424 2626 11490 2642
rect 13056 2642 13072 2644
rect 13106 2674 13122 2676
rect 14688 2676 14754 2692
rect 14688 2674 14704 2676
rect 13106 2644 14704 2674
rect 13106 2642 13122 2644
rect 13056 2626 13122 2642
rect 14688 2642 14704 2644
rect 14738 2674 14754 2676
rect 16320 2676 16386 2692
rect 16320 2674 16336 2676
rect 14738 2644 16336 2674
rect 14738 2642 14754 2644
rect 14688 2626 14754 2642
rect 16320 2642 16336 2644
rect 16370 2674 16386 2676
rect 17952 2676 18018 2692
rect 17952 2674 17968 2676
rect 16370 2644 17968 2674
rect 16370 2642 16386 2644
rect 16320 2626 16386 2642
rect 17952 2642 17968 2644
rect 18002 2674 18018 2676
rect 19584 2676 19650 2692
rect 19584 2674 19600 2676
rect 18002 2644 19600 2674
rect 18002 2642 18018 2644
rect 17952 2626 18018 2642
rect 19584 2642 19600 2644
rect 19634 2674 19650 2676
rect 21216 2676 21282 2692
rect 21216 2674 21232 2676
rect 19634 2644 21232 2674
rect 19634 2642 19650 2644
rect 19584 2626 19650 2642
rect 21216 2642 21232 2644
rect 21266 2674 21282 2676
rect 22848 2676 22914 2692
rect 22848 2674 22864 2676
rect 21266 2644 22864 2674
rect 21266 2642 21282 2644
rect 21216 2626 21282 2642
rect 22848 2642 22864 2644
rect 22898 2674 22914 2676
rect 24480 2676 24546 2692
rect 24480 2674 24496 2676
rect 22898 2644 24496 2674
rect 22898 2642 22914 2644
rect 22848 2626 22914 2642
rect 24480 2642 24496 2644
rect 24530 2674 24546 2676
rect 26112 2676 26178 2692
rect 26112 2674 26128 2676
rect 24530 2644 26128 2674
rect 24530 2642 24546 2644
rect 24480 2626 24546 2642
rect 26112 2642 26128 2644
rect 26162 2674 26178 2676
rect 27744 2676 27810 2692
rect 27744 2674 27760 2676
rect 26162 2644 27760 2674
rect 26162 2642 26178 2644
rect 26112 2626 26178 2642
rect 27744 2642 27760 2644
rect 27794 2674 27810 2676
rect 29376 2676 29442 2692
rect 29376 2674 29392 2676
rect 27794 2644 29392 2674
rect 27794 2642 27810 2644
rect 27744 2626 27810 2642
rect 29376 2642 29392 2644
rect 29426 2674 29442 2676
rect 31008 2676 31074 2692
rect 31008 2674 31024 2676
rect 29426 2644 31024 2674
rect 29426 2642 29442 2644
rect 29376 2626 29442 2642
rect 31008 2642 31024 2644
rect 31058 2674 31074 2676
rect 32640 2676 32706 2692
rect 32640 2674 32656 2676
rect 31058 2644 32656 2674
rect 31058 2642 31074 2644
rect 31008 2626 31074 2642
rect 32640 2642 32656 2644
rect 32690 2674 32706 2676
rect 34272 2676 34338 2692
rect 34272 2674 34288 2676
rect 32690 2644 34288 2674
rect 32690 2642 32706 2644
rect 32640 2626 32706 2642
rect 34272 2642 34288 2644
rect 34322 2674 34338 2676
rect 35904 2676 35970 2692
rect 35904 2674 35920 2676
rect 34322 2644 35920 2674
rect 34322 2642 34338 2644
rect 34272 2626 34338 2642
rect 35904 2642 35920 2644
rect 35954 2674 35970 2676
rect 37536 2676 37602 2692
rect 37536 2674 37552 2676
rect 35954 2644 37552 2674
rect 35954 2642 35970 2644
rect 35904 2626 35970 2642
rect 37536 2642 37552 2644
rect 37586 2674 37602 2676
rect 39168 2676 39234 2692
rect 39168 2674 39184 2676
rect 37586 2644 39184 2674
rect 37586 2642 37602 2644
rect 37536 2626 37602 2642
rect 39168 2642 39184 2644
rect 39218 2674 39234 2676
rect 40800 2676 40866 2692
rect 40800 2674 40816 2676
rect 39218 2644 40816 2674
rect 39218 2642 39234 2644
rect 39168 2626 39234 2642
rect 40800 2642 40816 2644
rect 40850 2674 40866 2676
rect 42432 2676 42498 2692
rect 42432 2674 42448 2676
rect 40850 2644 42448 2674
rect 40850 2642 40866 2644
rect 40800 2626 40866 2642
rect 42432 2642 42448 2644
rect 42482 2674 42498 2676
rect 44064 2676 44130 2692
rect 44064 2674 44080 2676
rect 42482 2644 44080 2674
rect 42482 2642 42498 2644
rect 42432 2626 42498 2642
rect 44064 2642 44080 2644
rect 44114 2674 44130 2676
rect 45696 2676 45762 2692
rect 45696 2674 45712 2676
rect 44114 2644 45712 2674
rect 44114 2642 44130 2644
rect 44064 2626 44130 2642
rect 45696 2642 45712 2644
rect 45746 2674 45762 2676
rect 47328 2676 47394 2692
rect 47328 2674 47344 2676
rect 45746 2644 47344 2674
rect 45746 2642 45762 2644
rect 45696 2626 45762 2642
rect 47328 2642 47344 2644
rect 47378 2674 47394 2676
rect 48960 2676 49026 2692
rect 48960 2674 48976 2676
rect 47378 2644 48976 2674
rect 47378 2642 47394 2644
rect 47328 2626 47394 2642
rect 48960 2642 48976 2644
rect 49010 2674 49026 2676
rect 50592 2676 50658 2692
rect 50592 2674 50608 2676
rect 49010 2644 50608 2674
rect 49010 2642 49026 2644
rect 48960 2626 49026 2642
rect 50592 2642 50608 2644
rect 50642 2674 50658 2676
rect 52224 2676 52290 2692
rect 52224 2674 52240 2676
rect 50642 2644 52240 2674
rect 50642 2642 50658 2644
rect 50592 2626 50658 2642
rect 52224 2642 52240 2644
rect 52274 2642 52290 2676
rect 52224 2626 52290 2642
rect 0 2472 66 2488
rect 0 2438 16 2472
rect 50 2470 66 2472
rect 1632 2472 1698 2488
rect 1632 2470 1648 2472
rect 50 2440 1648 2470
rect 50 2438 66 2440
rect 0 2422 66 2438
rect 1632 2438 1648 2440
rect 1682 2470 1698 2472
rect 3264 2472 3330 2488
rect 3264 2470 3280 2472
rect 1682 2440 3280 2470
rect 1682 2438 1698 2440
rect 1632 2422 1698 2438
rect 3264 2438 3280 2440
rect 3314 2470 3330 2472
rect 4896 2472 4962 2488
rect 4896 2470 4912 2472
rect 3314 2440 4912 2470
rect 3314 2438 3330 2440
rect 3264 2422 3330 2438
rect 4896 2438 4912 2440
rect 4946 2470 4962 2472
rect 6528 2472 6594 2488
rect 6528 2470 6544 2472
rect 4946 2440 6544 2470
rect 4946 2438 4962 2440
rect 4896 2422 4962 2438
rect 6528 2438 6544 2440
rect 6578 2470 6594 2472
rect 8160 2472 8226 2488
rect 8160 2470 8176 2472
rect 6578 2440 8176 2470
rect 6578 2438 6594 2440
rect 6528 2422 6594 2438
rect 8160 2438 8176 2440
rect 8210 2470 8226 2472
rect 9792 2472 9858 2488
rect 9792 2470 9808 2472
rect 8210 2440 9808 2470
rect 8210 2438 8226 2440
rect 8160 2422 8226 2438
rect 9792 2438 9808 2440
rect 9842 2470 9858 2472
rect 11424 2472 11490 2488
rect 11424 2470 11440 2472
rect 9842 2440 11440 2470
rect 9842 2438 9858 2440
rect 9792 2422 9858 2438
rect 11424 2438 11440 2440
rect 11474 2470 11490 2472
rect 13056 2472 13122 2488
rect 13056 2470 13072 2472
rect 11474 2440 13072 2470
rect 11474 2438 11490 2440
rect 11424 2422 11490 2438
rect 13056 2438 13072 2440
rect 13106 2470 13122 2472
rect 14688 2472 14754 2488
rect 14688 2470 14704 2472
rect 13106 2440 14704 2470
rect 13106 2438 13122 2440
rect 13056 2422 13122 2438
rect 14688 2438 14704 2440
rect 14738 2470 14754 2472
rect 16320 2472 16386 2488
rect 16320 2470 16336 2472
rect 14738 2440 16336 2470
rect 14738 2438 14754 2440
rect 14688 2422 14754 2438
rect 16320 2438 16336 2440
rect 16370 2470 16386 2472
rect 17952 2472 18018 2488
rect 17952 2470 17968 2472
rect 16370 2440 17968 2470
rect 16370 2438 16386 2440
rect 16320 2422 16386 2438
rect 17952 2438 17968 2440
rect 18002 2470 18018 2472
rect 19584 2472 19650 2488
rect 19584 2470 19600 2472
rect 18002 2440 19600 2470
rect 18002 2438 18018 2440
rect 17952 2422 18018 2438
rect 19584 2438 19600 2440
rect 19634 2470 19650 2472
rect 21216 2472 21282 2488
rect 21216 2470 21232 2472
rect 19634 2440 21232 2470
rect 19634 2438 19650 2440
rect 19584 2422 19650 2438
rect 21216 2438 21232 2440
rect 21266 2470 21282 2472
rect 22848 2472 22914 2488
rect 22848 2470 22864 2472
rect 21266 2440 22864 2470
rect 21266 2438 21282 2440
rect 21216 2422 21282 2438
rect 22848 2438 22864 2440
rect 22898 2470 22914 2472
rect 24480 2472 24546 2488
rect 24480 2470 24496 2472
rect 22898 2440 24496 2470
rect 22898 2438 22914 2440
rect 22848 2422 22914 2438
rect 24480 2438 24496 2440
rect 24530 2470 24546 2472
rect 26112 2472 26178 2488
rect 26112 2470 26128 2472
rect 24530 2440 26128 2470
rect 24530 2438 24546 2440
rect 24480 2422 24546 2438
rect 26112 2438 26128 2440
rect 26162 2470 26178 2472
rect 27744 2472 27810 2488
rect 27744 2470 27760 2472
rect 26162 2440 27760 2470
rect 26162 2438 26178 2440
rect 26112 2422 26178 2438
rect 27744 2438 27760 2440
rect 27794 2470 27810 2472
rect 29376 2472 29442 2488
rect 29376 2470 29392 2472
rect 27794 2440 29392 2470
rect 27794 2438 27810 2440
rect 27744 2422 27810 2438
rect 29376 2438 29392 2440
rect 29426 2470 29442 2472
rect 31008 2472 31074 2488
rect 31008 2470 31024 2472
rect 29426 2440 31024 2470
rect 29426 2438 29442 2440
rect 29376 2422 29442 2438
rect 31008 2438 31024 2440
rect 31058 2470 31074 2472
rect 32640 2472 32706 2488
rect 32640 2470 32656 2472
rect 31058 2440 32656 2470
rect 31058 2438 31074 2440
rect 31008 2422 31074 2438
rect 32640 2438 32656 2440
rect 32690 2470 32706 2472
rect 34272 2472 34338 2488
rect 34272 2470 34288 2472
rect 32690 2440 34288 2470
rect 32690 2438 32706 2440
rect 32640 2422 32706 2438
rect 34272 2438 34288 2440
rect 34322 2470 34338 2472
rect 35904 2472 35970 2488
rect 35904 2470 35920 2472
rect 34322 2440 35920 2470
rect 34322 2438 34338 2440
rect 34272 2422 34338 2438
rect 35904 2438 35920 2440
rect 35954 2470 35970 2472
rect 37536 2472 37602 2488
rect 37536 2470 37552 2472
rect 35954 2440 37552 2470
rect 35954 2438 35970 2440
rect 35904 2422 35970 2438
rect 37536 2438 37552 2440
rect 37586 2470 37602 2472
rect 39168 2472 39234 2488
rect 39168 2470 39184 2472
rect 37586 2440 39184 2470
rect 37586 2438 37602 2440
rect 37536 2422 37602 2438
rect 39168 2438 39184 2440
rect 39218 2470 39234 2472
rect 40800 2472 40866 2488
rect 40800 2470 40816 2472
rect 39218 2440 40816 2470
rect 39218 2438 39234 2440
rect 39168 2422 39234 2438
rect 40800 2438 40816 2440
rect 40850 2470 40866 2472
rect 42432 2472 42498 2488
rect 42432 2470 42448 2472
rect 40850 2440 42448 2470
rect 40850 2438 40866 2440
rect 40800 2422 40866 2438
rect 42432 2438 42448 2440
rect 42482 2470 42498 2472
rect 44064 2472 44130 2488
rect 44064 2470 44080 2472
rect 42482 2440 44080 2470
rect 42482 2438 42498 2440
rect 42432 2422 42498 2438
rect 44064 2438 44080 2440
rect 44114 2470 44130 2472
rect 45696 2472 45762 2488
rect 45696 2470 45712 2472
rect 44114 2440 45712 2470
rect 44114 2438 44130 2440
rect 44064 2422 44130 2438
rect 45696 2438 45712 2440
rect 45746 2470 45762 2472
rect 47328 2472 47394 2488
rect 47328 2470 47344 2472
rect 45746 2440 47344 2470
rect 45746 2438 45762 2440
rect 45696 2422 45762 2438
rect 47328 2438 47344 2440
rect 47378 2470 47394 2472
rect 48960 2472 49026 2488
rect 48960 2470 48976 2472
rect 47378 2440 48976 2470
rect 47378 2438 47394 2440
rect 47328 2422 47394 2438
rect 48960 2438 48976 2440
rect 49010 2470 49026 2472
rect 50592 2472 50658 2488
rect 50592 2470 50608 2472
rect 49010 2440 50608 2470
rect 49010 2438 49026 2440
rect 48960 2422 49026 2438
rect 50592 2438 50608 2440
rect 50642 2470 50658 2472
rect 52224 2472 52290 2488
rect 52224 2470 52240 2472
rect 50642 2440 52240 2470
rect 50642 2438 50658 2440
rect 50592 2422 50658 2438
rect 52224 2438 52240 2440
rect 52274 2438 52290 2472
rect 52224 2422 52290 2438
rect 0 2268 66 2284
rect 0 2234 16 2268
rect 50 2266 66 2268
rect 1632 2268 1698 2284
rect 1632 2266 1648 2268
rect 50 2236 1648 2266
rect 50 2234 66 2236
rect 0 2218 66 2234
rect 1632 2234 1648 2236
rect 1682 2266 1698 2268
rect 3264 2268 3330 2284
rect 3264 2266 3280 2268
rect 1682 2236 3280 2266
rect 1682 2234 1698 2236
rect 1632 2218 1698 2234
rect 3264 2234 3280 2236
rect 3314 2266 3330 2268
rect 4896 2268 4962 2284
rect 4896 2266 4912 2268
rect 3314 2236 4912 2266
rect 3314 2234 3330 2236
rect 3264 2218 3330 2234
rect 4896 2234 4912 2236
rect 4946 2266 4962 2268
rect 6528 2268 6594 2284
rect 6528 2266 6544 2268
rect 4946 2236 6544 2266
rect 4946 2234 4962 2236
rect 4896 2218 4962 2234
rect 6528 2234 6544 2236
rect 6578 2266 6594 2268
rect 8160 2268 8226 2284
rect 8160 2266 8176 2268
rect 6578 2236 8176 2266
rect 6578 2234 6594 2236
rect 6528 2218 6594 2234
rect 8160 2234 8176 2236
rect 8210 2266 8226 2268
rect 9792 2268 9858 2284
rect 9792 2266 9808 2268
rect 8210 2236 9808 2266
rect 8210 2234 8226 2236
rect 8160 2218 8226 2234
rect 9792 2234 9808 2236
rect 9842 2266 9858 2268
rect 11424 2268 11490 2284
rect 11424 2266 11440 2268
rect 9842 2236 11440 2266
rect 9842 2234 9858 2236
rect 9792 2218 9858 2234
rect 11424 2234 11440 2236
rect 11474 2266 11490 2268
rect 13056 2268 13122 2284
rect 13056 2266 13072 2268
rect 11474 2236 13072 2266
rect 11474 2234 11490 2236
rect 11424 2218 11490 2234
rect 13056 2234 13072 2236
rect 13106 2266 13122 2268
rect 14688 2268 14754 2284
rect 14688 2266 14704 2268
rect 13106 2236 14704 2266
rect 13106 2234 13122 2236
rect 13056 2218 13122 2234
rect 14688 2234 14704 2236
rect 14738 2266 14754 2268
rect 16320 2268 16386 2284
rect 16320 2266 16336 2268
rect 14738 2236 16336 2266
rect 14738 2234 14754 2236
rect 14688 2218 14754 2234
rect 16320 2234 16336 2236
rect 16370 2266 16386 2268
rect 17952 2268 18018 2284
rect 17952 2266 17968 2268
rect 16370 2236 17968 2266
rect 16370 2234 16386 2236
rect 16320 2218 16386 2234
rect 17952 2234 17968 2236
rect 18002 2266 18018 2268
rect 19584 2268 19650 2284
rect 19584 2266 19600 2268
rect 18002 2236 19600 2266
rect 18002 2234 18018 2236
rect 17952 2218 18018 2234
rect 19584 2234 19600 2236
rect 19634 2266 19650 2268
rect 21216 2268 21282 2284
rect 21216 2266 21232 2268
rect 19634 2236 21232 2266
rect 19634 2234 19650 2236
rect 19584 2218 19650 2234
rect 21216 2234 21232 2236
rect 21266 2266 21282 2268
rect 22848 2268 22914 2284
rect 22848 2266 22864 2268
rect 21266 2236 22864 2266
rect 21266 2234 21282 2236
rect 21216 2218 21282 2234
rect 22848 2234 22864 2236
rect 22898 2266 22914 2268
rect 24480 2268 24546 2284
rect 24480 2266 24496 2268
rect 22898 2236 24496 2266
rect 22898 2234 22914 2236
rect 22848 2218 22914 2234
rect 24480 2234 24496 2236
rect 24530 2266 24546 2268
rect 26112 2268 26178 2284
rect 26112 2266 26128 2268
rect 24530 2236 26128 2266
rect 24530 2234 24546 2236
rect 24480 2218 24546 2234
rect 26112 2234 26128 2236
rect 26162 2266 26178 2268
rect 27744 2268 27810 2284
rect 27744 2266 27760 2268
rect 26162 2236 27760 2266
rect 26162 2234 26178 2236
rect 26112 2218 26178 2234
rect 27744 2234 27760 2236
rect 27794 2266 27810 2268
rect 29376 2268 29442 2284
rect 29376 2266 29392 2268
rect 27794 2236 29392 2266
rect 27794 2234 27810 2236
rect 27744 2218 27810 2234
rect 29376 2234 29392 2236
rect 29426 2266 29442 2268
rect 31008 2268 31074 2284
rect 31008 2266 31024 2268
rect 29426 2236 31024 2266
rect 29426 2234 29442 2236
rect 29376 2218 29442 2234
rect 31008 2234 31024 2236
rect 31058 2266 31074 2268
rect 32640 2268 32706 2284
rect 32640 2266 32656 2268
rect 31058 2236 32656 2266
rect 31058 2234 31074 2236
rect 31008 2218 31074 2234
rect 32640 2234 32656 2236
rect 32690 2266 32706 2268
rect 34272 2268 34338 2284
rect 34272 2266 34288 2268
rect 32690 2236 34288 2266
rect 32690 2234 32706 2236
rect 32640 2218 32706 2234
rect 34272 2234 34288 2236
rect 34322 2266 34338 2268
rect 35904 2268 35970 2284
rect 35904 2266 35920 2268
rect 34322 2236 35920 2266
rect 34322 2234 34338 2236
rect 34272 2218 34338 2234
rect 35904 2234 35920 2236
rect 35954 2266 35970 2268
rect 37536 2268 37602 2284
rect 37536 2266 37552 2268
rect 35954 2236 37552 2266
rect 35954 2234 35970 2236
rect 35904 2218 35970 2234
rect 37536 2234 37552 2236
rect 37586 2266 37602 2268
rect 39168 2268 39234 2284
rect 39168 2266 39184 2268
rect 37586 2236 39184 2266
rect 37586 2234 37602 2236
rect 37536 2218 37602 2234
rect 39168 2234 39184 2236
rect 39218 2266 39234 2268
rect 40800 2268 40866 2284
rect 40800 2266 40816 2268
rect 39218 2236 40816 2266
rect 39218 2234 39234 2236
rect 39168 2218 39234 2234
rect 40800 2234 40816 2236
rect 40850 2266 40866 2268
rect 42432 2268 42498 2284
rect 42432 2266 42448 2268
rect 40850 2236 42448 2266
rect 40850 2234 40866 2236
rect 40800 2218 40866 2234
rect 42432 2234 42448 2236
rect 42482 2266 42498 2268
rect 44064 2268 44130 2284
rect 44064 2266 44080 2268
rect 42482 2236 44080 2266
rect 42482 2234 42498 2236
rect 42432 2218 42498 2234
rect 44064 2234 44080 2236
rect 44114 2266 44130 2268
rect 45696 2268 45762 2284
rect 45696 2266 45712 2268
rect 44114 2236 45712 2266
rect 44114 2234 44130 2236
rect 44064 2218 44130 2234
rect 45696 2234 45712 2236
rect 45746 2266 45762 2268
rect 47328 2268 47394 2284
rect 47328 2266 47344 2268
rect 45746 2236 47344 2266
rect 45746 2234 45762 2236
rect 45696 2218 45762 2234
rect 47328 2234 47344 2236
rect 47378 2266 47394 2268
rect 48960 2268 49026 2284
rect 48960 2266 48976 2268
rect 47378 2236 48976 2266
rect 47378 2234 47394 2236
rect 47328 2218 47394 2234
rect 48960 2234 48976 2236
rect 49010 2266 49026 2268
rect 50592 2268 50658 2284
rect 50592 2266 50608 2268
rect 49010 2236 50608 2266
rect 49010 2234 49026 2236
rect 48960 2218 49026 2234
rect 50592 2234 50608 2236
rect 50642 2266 50658 2268
rect 52224 2268 52290 2284
rect 52224 2266 52240 2268
rect 50642 2236 52240 2266
rect 50642 2234 50658 2236
rect 50592 2218 50658 2234
rect 52224 2234 52240 2236
rect 52274 2234 52290 2268
rect 52224 2218 52290 2234
rect 0 2064 66 2080
rect 0 2030 16 2064
rect 50 2062 66 2064
rect 1632 2064 1698 2080
rect 1632 2062 1648 2064
rect 50 2032 1648 2062
rect 50 2030 66 2032
rect 0 2014 66 2030
rect 1632 2030 1648 2032
rect 1682 2062 1698 2064
rect 3264 2064 3330 2080
rect 3264 2062 3280 2064
rect 1682 2032 3280 2062
rect 1682 2030 1698 2032
rect 1632 2014 1698 2030
rect 3264 2030 3280 2032
rect 3314 2062 3330 2064
rect 4896 2064 4962 2080
rect 4896 2062 4912 2064
rect 3314 2032 4912 2062
rect 3314 2030 3330 2032
rect 3264 2014 3330 2030
rect 4896 2030 4912 2032
rect 4946 2062 4962 2064
rect 6528 2064 6594 2080
rect 6528 2062 6544 2064
rect 4946 2032 6544 2062
rect 4946 2030 4962 2032
rect 4896 2014 4962 2030
rect 6528 2030 6544 2032
rect 6578 2062 6594 2064
rect 8160 2064 8226 2080
rect 8160 2062 8176 2064
rect 6578 2032 8176 2062
rect 6578 2030 6594 2032
rect 6528 2014 6594 2030
rect 8160 2030 8176 2032
rect 8210 2062 8226 2064
rect 9792 2064 9858 2080
rect 9792 2062 9808 2064
rect 8210 2032 9808 2062
rect 8210 2030 8226 2032
rect 8160 2014 8226 2030
rect 9792 2030 9808 2032
rect 9842 2062 9858 2064
rect 11424 2064 11490 2080
rect 11424 2062 11440 2064
rect 9842 2032 11440 2062
rect 9842 2030 9858 2032
rect 9792 2014 9858 2030
rect 11424 2030 11440 2032
rect 11474 2062 11490 2064
rect 13056 2064 13122 2080
rect 13056 2062 13072 2064
rect 11474 2032 13072 2062
rect 11474 2030 11490 2032
rect 11424 2014 11490 2030
rect 13056 2030 13072 2032
rect 13106 2062 13122 2064
rect 14688 2064 14754 2080
rect 14688 2062 14704 2064
rect 13106 2032 14704 2062
rect 13106 2030 13122 2032
rect 13056 2014 13122 2030
rect 14688 2030 14704 2032
rect 14738 2062 14754 2064
rect 16320 2064 16386 2080
rect 16320 2062 16336 2064
rect 14738 2032 16336 2062
rect 14738 2030 14754 2032
rect 14688 2014 14754 2030
rect 16320 2030 16336 2032
rect 16370 2062 16386 2064
rect 17952 2064 18018 2080
rect 17952 2062 17968 2064
rect 16370 2032 17968 2062
rect 16370 2030 16386 2032
rect 16320 2014 16386 2030
rect 17952 2030 17968 2032
rect 18002 2062 18018 2064
rect 19584 2064 19650 2080
rect 19584 2062 19600 2064
rect 18002 2032 19600 2062
rect 18002 2030 18018 2032
rect 17952 2014 18018 2030
rect 19584 2030 19600 2032
rect 19634 2062 19650 2064
rect 21216 2064 21282 2080
rect 21216 2062 21232 2064
rect 19634 2032 21232 2062
rect 19634 2030 19650 2032
rect 19584 2014 19650 2030
rect 21216 2030 21232 2032
rect 21266 2062 21282 2064
rect 22848 2064 22914 2080
rect 22848 2062 22864 2064
rect 21266 2032 22864 2062
rect 21266 2030 21282 2032
rect 21216 2014 21282 2030
rect 22848 2030 22864 2032
rect 22898 2062 22914 2064
rect 24480 2064 24546 2080
rect 24480 2062 24496 2064
rect 22898 2032 24496 2062
rect 22898 2030 22914 2032
rect 22848 2014 22914 2030
rect 24480 2030 24496 2032
rect 24530 2062 24546 2064
rect 26112 2064 26178 2080
rect 26112 2062 26128 2064
rect 24530 2032 26128 2062
rect 24530 2030 24546 2032
rect 24480 2014 24546 2030
rect 26112 2030 26128 2032
rect 26162 2062 26178 2064
rect 27744 2064 27810 2080
rect 27744 2062 27760 2064
rect 26162 2032 27760 2062
rect 26162 2030 26178 2032
rect 26112 2014 26178 2030
rect 27744 2030 27760 2032
rect 27794 2062 27810 2064
rect 29376 2064 29442 2080
rect 29376 2062 29392 2064
rect 27794 2032 29392 2062
rect 27794 2030 27810 2032
rect 27744 2014 27810 2030
rect 29376 2030 29392 2032
rect 29426 2062 29442 2064
rect 31008 2064 31074 2080
rect 31008 2062 31024 2064
rect 29426 2032 31024 2062
rect 29426 2030 29442 2032
rect 29376 2014 29442 2030
rect 31008 2030 31024 2032
rect 31058 2062 31074 2064
rect 32640 2064 32706 2080
rect 32640 2062 32656 2064
rect 31058 2032 32656 2062
rect 31058 2030 31074 2032
rect 31008 2014 31074 2030
rect 32640 2030 32656 2032
rect 32690 2062 32706 2064
rect 34272 2064 34338 2080
rect 34272 2062 34288 2064
rect 32690 2032 34288 2062
rect 32690 2030 32706 2032
rect 32640 2014 32706 2030
rect 34272 2030 34288 2032
rect 34322 2062 34338 2064
rect 35904 2064 35970 2080
rect 35904 2062 35920 2064
rect 34322 2032 35920 2062
rect 34322 2030 34338 2032
rect 34272 2014 34338 2030
rect 35904 2030 35920 2032
rect 35954 2062 35970 2064
rect 37536 2064 37602 2080
rect 37536 2062 37552 2064
rect 35954 2032 37552 2062
rect 35954 2030 35970 2032
rect 35904 2014 35970 2030
rect 37536 2030 37552 2032
rect 37586 2062 37602 2064
rect 39168 2064 39234 2080
rect 39168 2062 39184 2064
rect 37586 2032 39184 2062
rect 37586 2030 37602 2032
rect 37536 2014 37602 2030
rect 39168 2030 39184 2032
rect 39218 2062 39234 2064
rect 40800 2064 40866 2080
rect 40800 2062 40816 2064
rect 39218 2032 40816 2062
rect 39218 2030 39234 2032
rect 39168 2014 39234 2030
rect 40800 2030 40816 2032
rect 40850 2062 40866 2064
rect 42432 2064 42498 2080
rect 42432 2062 42448 2064
rect 40850 2032 42448 2062
rect 40850 2030 40866 2032
rect 40800 2014 40866 2030
rect 42432 2030 42448 2032
rect 42482 2062 42498 2064
rect 44064 2064 44130 2080
rect 44064 2062 44080 2064
rect 42482 2032 44080 2062
rect 42482 2030 42498 2032
rect 42432 2014 42498 2030
rect 44064 2030 44080 2032
rect 44114 2062 44130 2064
rect 45696 2064 45762 2080
rect 45696 2062 45712 2064
rect 44114 2032 45712 2062
rect 44114 2030 44130 2032
rect 44064 2014 44130 2030
rect 45696 2030 45712 2032
rect 45746 2062 45762 2064
rect 47328 2064 47394 2080
rect 47328 2062 47344 2064
rect 45746 2032 47344 2062
rect 45746 2030 45762 2032
rect 45696 2014 45762 2030
rect 47328 2030 47344 2032
rect 47378 2062 47394 2064
rect 48960 2064 49026 2080
rect 48960 2062 48976 2064
rect 47378 2032 48976 2062
rect 47378 2030 47394 2032
rect 47328 2014 47394 2030
rect 48960 2030 48976 2032
rect 49010 2062 49026 2064
rect 50592 2064 50658 2080
rect 50592 2062 50608 2064
rect 49010 2032 50608 2062
rect 49010 2030 49026 2032
rect 48960 2014 49026 2030
rect 50592 2030 50608 2032
rect 50642 2062 50658 2064
rect 52224 2064 52290 2080
rect 52224 2062 52240 2064
rect 50642 2032 52240 2062
rect 50642 2030 50658 2032
rect 50592 2014 50658 2030
rect 52224 2030 52240 2032
rect 52274 2030 52290 2064
rect 52224 2014 52290 2030
rect 0 1860 66 1876
rect 0 1826 16 1860
rect 50 1858 66 1860
rect 1632 1860 1698 1876
rect 1632 1858 1648 1860
rect 50 1828 1648 1858
rect 50 1826 66 1828
rect 0 1810 66 1826
rect 1632 1826 1648 1828
rect 1682 1858 1698 1860
rect 3264 1860 3330 1876
rect 3264 1858 3280 1860
rect 1682 1828 3280 1858
rect 1682 1826 1698 1828
rect 1632 1810 1698 1826
rect 3264 1826 3280 1828
rect 3314 1858 3330 1860
rect 4896 1860 4962 1876
rect 4896 1858 4912 1860
rect 3314 1828 4912 1858
rect 3314 1826 3330 1828
rect 3264 1810 3330 1826
rect 4896 1826 4912 1828
rect 4946 1858 4962 1860
rect 6528 1860 6594 1876
rect 6528 1858 6544 1860
rect 4946 1828 6544 1858
rect 4946 1826 4962 1828
rect 4896 1810 4962 1826
rect 6528 1826 6544 1828
rect 6578 1858 6594 1860
rect 8160 1860 8226 1876
rect 8160 1858 8176 1860
rect 6578 1828 8176 1858
rect 6578 1826 6594 1828
rect 6528 1810 6594 1826
rect 8160 1826 8176 1828
rect 8210 1858 8226 1860
rect 9792 1860 9858 1876
rect 9792 1858 9808 1860
rect 8210 1828 9808 1858
rect 8210 1826 8226 1828
rect 8160 1810 8226 1826
rect 9792 1826 9808 1828
rect 9842 1858 9858 1860
rect 11424 1860 11490 1876
rect 11424 1858 11440 1860
rect 9842 1828 11440 1858
rect 9842 1826 9858 1828
rect 9792 1810 9858 1826
rect 11424 1826 11440 1828
rect 11474 1858 11490 1860
rect 13056 1860 13122 1876
rect 13056 1858 13072 1860
rect 11474 1828 13072 1858
rect 11474 1826 11490 1828
rect 11424 1810 11490 1826
rect 13056 1826 13072 1828
rect 13106 1858 13122 1860
rect 14688 1860 14754 1876
rect 14688 1858 14704 1860
rect 13106 1828 14704 1858
rect 13106 1826 13122 1828
rect 13056 1810 13122 1826
rect 14688 1826 14704 1828
rect 14738 1858 14754 1860
rect 16320 1860 16386 1876
rect 16320 1858 16336 1860
rect 14738 1828 16336 1858
rect 14738 1826 14754 1828
rect 14688 1810 14754 1826
rect 16320 1826 16336 1828
rect 16370 1858 16386 1860
rect 17952 1860 18018 1876
rect 17952 1858 17968 1860
rect 16370 1828 17968 1858
rect 16370 1826 16386 1828
rect 16320 1810 16386 1826
rect 17952 1826 17968 1828
rect 18002 1858 18018 1860
rect 19584 1860 19650 1876
rect 19584 1858 19600 1860
rect 18002 1828 19600 1858
rect 18002 1826 18018 1828
rect 17952 1810 18018 1826
rect 19584 1826 19600 1828
rect 19634 1858 19650 1860
rect 21216 1860 21282 1876
rect 21216 1858 21232 1860
rect 19634 1828 21232 1858
rect 19634 1826 19650 1828
rect 19584 1810 19650 1826
rect 21216 1826 21232 1828
rect 21266 1858 21282 1860
rect 22848 1860 22914 1876
rect 22848 1858 22864 1860
rect 21266 1828 22864 1858
rect 21266 1826 21282 1828
rect 21216 1810 21282 1826
rect 22848 1826 22864 1828
rect 22898 1858 22914 1860
rect 24480 1860 24546 1876
rect 24480 1858 24496 1860
rect 22898 1828 24496 1858
rect 22898 1826 22914 1828
rect 22848 1810 22914 1826
rect 24480 1826 24496 1828
rect 24530 1858 24546 1860
rect 26112 1860 26178 1876
rect 26112 1858 26128 1860
rect 24530 1828 26128 1858
rect 24530 1826 24546 1828
rect 24480 1810 24546 1826
rect 26112 1826 26128 1828
rect 26162 1858 26178 1860
rect 27744 1860 27810 1876
rect 27744 1858 27760 1860
rect 26162 1828 27760 1858
rect 26162 1826 26178 1828
rect 26112 1810 26178 1826
rect 27744 1826 27760 1828
rect 27794 1858 27810 1860
rect 29376 1860 29442 1876
rect 29376 1858 29392 1860
rect 27794 1828 29392 1858
rect 27794 1826 27810 1828
rect 27744 1810 27810 1826
rect 29376 1826 29392 1828
rect 29426 1858 29442 1860
rect 31008 1860 31074 1876
rect 31008 1858 31024 1860
rect 29426 1828 31024 1858
rect 29426 1826 29442 1828
rect 29376 1810 29442 1826
rect 31008 1826 31024 1828
rect 31058 1858 31074 1860
rect 32640 1860 32706 1876
rect 32640 1858 32656 1860
rect 31058 1828 32656 1858
rect 31058 1826 31074 1828
rect 31008 1810 31074 1826
rect 32640 1826 32656 1828
rect 32690 1858 32706 1860
rect 34272 1860 34338 1876
rect 34272 1858 34288 1860
rect 32690 1828 34288 1858
rect 32690 1826 32706 1828
rect 32640 1810 32706 1826
rect 34272 1826 34288 1828
rect 34322 1858 34338 1860
rect 35904 1860 35970 1876
rect 35904 1858 35920 1860
rect 34322 1828 35920 1858
rect 34322 1826 34338 1828
rect 34272 1810 34338 1826
rect 35904 1826 35920 1828
rect 35954 1858 35970 1860
rect 37536 1860 37602 1876
rect 37536 1858 37552 1860
rect 35954 1828 37552 1858
rect 35954 1826 35970 1828
rect 35904 1810 35970 1826
rect 37536 1826 37552 1828
rect 37586 1858 37602 1860
rect 39168 1860 39234 1876
rect 39168 1858 39184 1860
rect 37586 1828 39184 1858
rect 37586 1826 37602 1828
rect 37536 1810 37602 1826
rect 39168 1826 39184 1828
rect 39218 1858 39234 1860
rect 40800 1860 40866 1876
rect 40800 1858 40816 1860
rect 39218 1828 40816 1858
rect 39218 1826 39234 1828
rect 39168 1810 39234 1826
rect 40800 1826 40816 1828
rect 40850 1858 40866 1860
rect 42432 1860 42498 1876
rect 42432 1858 42448 1860
rect 40850 1828 42448 1858
rect 40850 1826 40866 1828
rect 40800 1810 40866 1826
rect 42432 1826 42448 1828
rect 42482 1858 42498 1860
rect 44064 1860 44130 1876
rect 44064 1858 44080 1860
rect 42482 1828 44080 1858
rect 42482 1826 42498 1828
rect 42432 1810 42498 1826
rect 44064 1826 44080 1828
rect 44114 1858 44130 1860
rect 45696 1860 45762 1876
rect 45696 1858 45712 1860
rect 44114 1828 45712 1858
rect 44114 1826 44130 1828
rect 44064 1810 44130 1826
rect 45696 1826 45712 1828
rect 45746 1858 45762 1860
rect 47328 1860 47394 1876
rect 47328 1858 47344 1860
rect 45746 1828 47344 1858
rect 45746 1826 45762 1828
rect 45696 1810 45762 1826
rect 47328 1826 47344 1828
rect 47378 1858 47394 1860
rect 48960 1860 49026 1876
rect 48960 1858 48976 1860
rect 47378 1828 48976 1858
rect 47378 1826 47394 1828
rect 47328 1810 47394 1826
rect 48960 1826 48976 1828
rect 49010 1858 49026 1860
rect 50592 1860 50658 1876
rect 50592 1858 50608 1860
rect 49010 1828 50608 1858
rect 49010 1826 49026 1828
rect 48960 1810 49026 1826
rect 50592 1826 50608 1828
rect 50642 1858 50658 1860
rect 52224 1860 52290 1876
rect 52224 1858 52240 1860
rect 50642 1828 52240 1858
rect 50642 1826 50658 1828
rect 50592 1810 50658 1826
rect 52224 1826 52240 1828
rect 52274 1826 52290 1860
rect 52224 1810 52290 1826
rect 0 1656 66 1672
rect 0 1622 16 1656
rect 50 1654 66 1656
rect 1632 1656 1698 1672
rect 1632 1654 1648 1656
rect 50 1624 1648 1654
rect 50 1622 66 1624
rect 0 1606 66 1622
rect 1632 1622 1648 1624
rect 1682 1654 1698 1656
rect 3264 1656 3330 1672
rect 3264 1654 3280 1656
rect 1682 1624 3280 1654
rect 1682 1622 1698 1624
rect 1632 1606 1698 1622
rect 3264 1622 3280 1624
rect 3314 1654 3330 1656
rect 4896 1656 4962 1672
rect 4896 1654 4912 1656
rect 3314 1624 4912 1654
rect 3314 1622 3330 1624
rect 3264 1606 3330 1622
rect 4896 1622 4912 1624
rect 4946 1654 4962 1656
rect 6528 1656 6594 1672
rect 6528 1654 6544 1656
rect 4946 1624 6544 1654
rect 4946 1622 4962 1624
rect 4896 1606 4962 1622
rect 6528 1622 6544 1624
rect 6578 1654 6594 1656
rect 8160 1656 8226 1672
rect 8160 1654 8176 1656
rect 6578 1624 8176 1654
rect 6578 1622 6594 1624
rect 6528 1606 6594 1622
rect 8160 1622 8176 1624
rect 8210 1654 8226 1656
rect 9792 1656 9858 1672
rect 9792 1654 9808 1656
rect 8210 1624 9808 1654
rect 8210 1622 8226 1624
rect 8160 1606 8226 1622
rect 9792 1622 9808 1624
rect 9842 1654 9858 1656
rect 11424 1656 11490 1672
rect 11424 1654 11440 1656
rect 9842 1624 11440 1654
rect 9842 1622 9858 1624
rect 9792 1606 9858 1622
rect 11424 1622 11440 1624
rect 11474 1654 11490 1656
rect 13056 1656 13122 1672
rect 13056 1654 13072 1656
rect 11474 1624 13072 1654
rect 11474 1622 11490 1624
rect 11424 1606 11490 1622
rect 13056 1622 13072 1624
rect 13106 1654 13122 1656
rect 14688 1656 14754 1672
rect 14688 1654 14704 1656
rect 13106 1624 14704 1654
rect 13106 1622 13122 1624
rect 13056 1606 13122 1622
rect 14688 1622 14704 1624
rect 14738 1654 14754 1656
rect 16320 1656 16386 1672
rect 16320 1654 16336 1656
rect 14738 1624 16336 1654
rect 14738 1622 14754 1624
rect 14688 1606 14754 1622
rect 16320 1622 16336 1624
rect 16370 1654 16386 1656
rect 17952 1656 18018 1672
rect 17952 1654 17968 1656
rect 16370 1624 17968 1654
rect 16370 1622 16386 1624
rect 16320 1606 16386 1622
rect 17952 1622 17968 1624
rect 18002 1654 18018 1656
rect 19584 1656 19650 1672
rect 19584 1654 19600 1656
rect 18002 1624 19600 1654
rect 18002 1622 18018 1624
rect 17952 1606 18018 1622
rect 19584 1622 19600 1624
rect 19634 1654 19650 1656
rect 21216 1656 21282 1672
rect 21216 1654 21232 1656
rect 19634 1624 21232 1654
rect 19634 1622 19650 1624
rect 19584 1606 19650 1622
rect 21216 1622 21232 1624
rect 21266 1654 21282 1656
rect 22848 1656 22914 1672
rect 22848 1654 22864 1656
rect 21266 1624 22864 1654
rect 21266 1622 21282 1624
rect 21216 1606 21282 1622
rect 22848 1622 22864 1624
rect 22898 1654 22914 1656
rect 24480 1656 24546 1672
rect 24480 1654 24496 1656
rect 22898 1624 24496 1654
rect 22898 1622 22914 1624
rect 22848 1606 22914 1622
rect 24480 1622 24496 1624
rect 24530 1654 24546 1656
rect 26112 1656 26178 1672
rect 26112 1654 26128 1656
rect 24530 1624 26128 1654
rect 24530 1622 24546 1624
rect 24480 1606 24546 1622
rect 26112 1622 26128 1624
rect 26162 1654 26178 1656
rect 27744 1656 27810 1672
rect 27744 1654 27760 1656
rect 26162 1624 27760 1654
rect 26162 1622 26178 1624
rect 26112 1606 26178 1622
rect 27744 1622 27760 1624
rect 27794 1654 27810 1656
rect 29376 1656 29442 1672
rect 29376 1654 29392 1656
rect 27794 1624 29392 1654
rect 27794 1622 27810 1624
rect 27744 1606 27810 1622
rect 29376 1622 29392 1624
rect 29426 1654 29442 1656
rect 31008 1656 31074 1672
rect 31008 1654 31024 1656
rect 29426 1624 31024 1654
rect 29426 1622 29442 1624
rect 29376 1606 29442 1622
rect 31008 1622 31024 1624
rect 31058 1654 31074 1656
rect 32640 1656 32706 1672
rect 32640 1654 32656 1656
rect 31058 1624 32656 1654
rect 31058 1622 31074 1624
rect 31008 1606 31074 1622
rect 32640 1622 32656 1624
rect 32690 1654 32706 1656
rect 34272 1656 34338 1672
rect 34272 1654 34288 1656
rect 32690 1624 34288 1654
rect 32690 1622 32706 1624
rect 32640 1606 32706 1622
rect 34272 1622 34288 1624
rect 34322 1654 34338 1656
rect 35904 1656 35970 1672
rect 35904 1654 35920 1656
rect 34322 1624 35920 1654
rect 34322 1622 34338 1624
rect 34272 1606 34338 1622
rect 35904 1622 35920 1624
rect 35954 1654 35970 1656
rect 37536 1656 37602 1672
rect 37536 1654 37552 1656
rect 35954 1624 37552 1654
rect 35954 1622 35970 1624
rect 35904 1606 35970 1622
rect 37536 1622 37552 1624
rect 37586 1654 37602 1656
rect 39168 1656 39234 1672
rect 39168 1654 39184 1656
rect 37586 1624 39184 1654
rect 37586 1622 37602 1624
rect 37536 1606 37602 1622
rect 39168 1622 39184 1624
rect 39218 1654 39234 1656
rect 40800 1656 40866 1672
rect 40800 1654 40816 1656
rect 39218 1624 40816 1654
rect 39218 1622 39234 1624
rect 39168 1606 39234 1622
rect 40800 1622 40816 1624
rect 40850 1654 40866 1656
rect 42432 1656 42498 1672
rect 42432 1654 42448 1656
rect 40850 1624 42448 1654
rect 40850 1622 40866 1624
rect 40800 1606 40866 1622
rect 42432 1622 42448 1624
rect 42482 1654 42498 1656
rect 44064 1656 44130 1672
rect 44064 1654 44080 1656
rect 42482 1624 44080 1654
rect 42482 1622 42498 1624
rect 42432 1606 42498 1622
rect 44064 1622 44080 1624
rect 44114 1654 44130 1656
rect 45696 1656 45762 1672
rect 45696 1654 45712 1656
rect 44114 1624 45712 1654
rect 44114 1622 44130 1624
rect 44064 1606 44130 1622
rect 45696 1622 45712 1624
rect 45746 1654 45762 1656
rect 47328 1656 47394 1672
rect 47328 1654 47344 1656
rect 45746 1624 47344 1654
rect 45746 1622 45762 1624
rect 45696 1606 45762 1622
rect 47328 1622 47344 1624
rect 47378 1654 47394 1656
rect 48960 1656 49026 1672
rect 48960 1654 48976 1656
rect 47378 1624 48976 1654
rect 47378 1622 47394 1624
rect 47328 1606 47394 1622
rect 48960 1622 48976 1624
rect 49010 1654 49026 1656
rect 50592 1656 50658 1672
rect 50592 1654 50608 1656
rect 49010 1624 50608 1654
rect 49010 1622 49026 1624
rect 48960 1606 49026 1622
rect 50592 1622 50608 1624
rect 50642 1654 50658 1656
rect 52224 1656 52290 1672
rect 52224 1654 52240 1656
rect 50642 1624 52240 1654
rect 50642 1622 50658 1624
rect 50592 1606 50658 1622
rect 52224 1622 52240 1624
rect 52274 1622 52290 1656
rect 52224 1606 52290 1622
rect 0 1452 66 1468
rect 0 1418 16 1452
rect 50 1450 66 1452
rect 1632 1452 1698 1468
rect 1632 1450 1648 1452
rect 50 1420 1648 1450
rect 50 1418 66 1420
rect 0 1402 66 1418
rect 1632 1418 1648 1420
rect 1682 1450 1698 1452
rect 3264 1452 3330 1468
rect 3264 1450 3280 1452
rect 1682 1420 3280 1450
rect 1682 1418 1698 1420
rect 1632 1402 1698 1418
rect 3264 1418 3280 1420
rect 3314 1450 3330 1452
rect 4896 1452 4962 1468
rect 4896 1450 4912 1452
rect 3314 1420 4912 1450
rect 3314 1418 3330 1420
rect 3264 1402 3330 1418
rect 4896 1418 4912 1420
rect 4946 1450 4962 1452
rect 6528 1452 6594 1468
rect 6528 1450 6544 1452
rect 4946 1420 6544 1450
rect 4946 1418 4962 1420
rect 4896 1402 4962 1418
rect 6528 1418 6544 1420
rect 6578 1450 6594 1452
rect 8160 1452 8226 1468
rect 8160 1450 8176 1452
rect 6578 1420 8176 1450
rect 6578 1418 6594 1420
rect 6528 1402 6594 1418
rect 8160 1418 8176 1420
rect 8210 1450 8226 1452
rect 9792 1452 9858 1468
rect 9792 1450 9808 1452
rect 8210 1420 9808 1450
rect 8210 1418 8226 1420
rect 8160 1402 8226 1418
rect 9792 1418 9808 1420
rect 9842 1450 9858 1452
rect 11424 1452 11490 1468
rect 11424 1450 11440 1452
rect 9842 1420 11440 1450
rect 9842 1418 9858 1420
rect 9792 1402 9858 1418
rect 11424 1418 11440 1420
rect 11474 1450 11490 1452
rect 13056 1452 13122 1468
rect 13056 1450 13072 1452
rect 11474 1420 13072 1450
rect 11474 1418 11490 1420
rect 11424 1402 11490 1418
rect 13056 1418 13072 1420
rect 13106 1450 13122 1452
rect 14688 1452 14754 1468
rect 14688 1450 14704 1452
rect 13106 1420 14704 1450
rect 13106 1418 13122 1420
rect 13056 1402 13122 1418
rect 14688 1418 14704 1420
rect 14738 1450 14754 1452
rect 16320 1452 16386 1468
rect 16320 1450 16336 1452
rect 14738 1420 16336 1450
rect 14738 1418 14754 1420
rect 14688 1402 14754 1418
rect 16320 1418 16336 1420
rect 16370 1450 16386 1452
rect 17952 1452 18018 1468
rect 17952 1450 17968 1452
rect 16370 1420 17968 1450
rect 16370 1418 16386 1420
rect 16320 1402 16386 1418
rect 17952 1418 17968 1420
rect 18002 1450 18018 1452
rect 19584 1452 19650 1468
rect 19584 1450 19600 1452
rect 18002 1420 19600 1450
rect 18002 1418 18018 1420
rect 17952 1402 18018 1418
rect 19584 1418 19600 1420
rect 19634 1450 19650 1452
rect 21216 1452 21282 1468
rect 21216 1450 21232 1452
rect 19634 1420 21232 1450
rect 19634 1418 19650 1420
rect 19584 1402 19650 1418
rect 21216 1418 21232 1420
rect 21266 1450 21282 1452
rect 22848 1452 22914 1468
rect 22848 1450 22864 1452
rect 21266 1420 22864 1450
rect 21266 1418 21282 1420
rect 21216 1402 21282 1418
rect 22848 1418 22864 1420
rect 22898 1450 22914 1452
rect 24480 1452 24546 1468
rect 24480 1450 24496 1452
rect 22898 1420 24496 1450
rect 22898 1418 22914 1420
rect 22848 1402 22914 1418
rect 24480 1418 24496 1420
rect 24530 1450 24546 1452
rect 26112 1452 26178 1468
rect 26112 1450 26128 1452
rect 24530 1420 26128 1450
rect 24530 1418 24546 1420
rect 24480 1402 24546 1418
rect 26112 1418 26128 1420
rect 26162 1450 26178 1452
rect 27744 1452 27810 1468
rect 27744 1450 27760 1452
rect 26162 1420 27760 1450
rect 26162 1418 26178 1420
rect 26112 1402 26178 1418
rect 27744 1418 27760 1420
rect 27794 1450 27810 1452
rect 29376 1452 29442 1468
rect 29376 1450 29392 1452
rect 27794 1420 29392 1450
rect 27794 1418 27810 1420
rect 27744 1402 27810 1418
rect 29376 1418 29392 1420
rect 29426 1450 29442 1452
rect 31008 1452 31074 1468
rect 31008 1450 31024 1452
rect 29426 1420 31024 1450
rect 29426 1418 29442 1420
rect 29376 1402 29442 1418
rect 31008 1418 31024 1420
rect 31058 1450 31074 1452
rect 32640 1452 32706 1468
rect 32640 1450 32656 1452
rect 31058 1420 32656 1450
rect 31058 1418 31074 1420
rect 31008 1402 31074 1418
rect 32640 1418 32656 1420
rect 32690 1450 32706 1452
rect 34272 1452 34338 1468
rect 34272 1450 34288 1452
rect 32690 1420 34288 1450
rect 32690 1418 32706 1420
rect 32640 1402 32706 1418
rect 34272 1418 34288 1420
rect 34322 1450 34338 1452
rect 35904 1452 35970 1468
rect 35904 1450 35920 1452
rect 34322 1420 35920 1450
rect 34322 1418 34338 1420
rect 34272 1402 34338 1418
rect 35904 1418 35920 1420
rect 35954 1450 35970 1452
rect 37536 1452 37602 1468
rect 37536 1450 37552 1452
rect 35954 1420 37552 1450
rect 35954 1418 35970 1420
rect 35904 1402 35970 1418
rect 37536 1418 37552 1420
rect 37586 1450 37602 1452
rect 39168 1452 39234 1468
rect 39168 1450 39184 1452
rect 37586 1420 39184 1450
rect 37586 1418 37602 1420
rect 37536 1402 37602 1418
rect 39168 1418 39184 1420
rect 39218 1450 39234 1452
rect 40800 1452 40866 1468
rect 40800 1450 40816 1452
rect 39218 1420 40816 1450
rect 39218 1418 39234 1420
rect 39168 1402 39234 1418
rect 40800 1418 40816 1420
rect 40850 1450 40866 1452
rect 42432 1452 42498 1468
rect 42432 1450 42448 1452
rect 40850 1420 42448 1450
rect 40850 1418 40866 1420
rect 40800 1402 40866 1418
rect 42432 1418 42448 1420
rect 42482 1450 42498 1452
rect 44064 1452 44130 1468
rect 44064 1450 44080 1452
rect 42482 1420 44080 1450
rect 42482 1418 42498 1420
rect 42432 1402 42498 1418
rect 44064 1418 44080 1420
rect 44114 1450 44130 1452
rect 45696 1452 45762 1468
rect 45696 1450 45712 1452
rect 44114 1420 45712 1450
rect 44114 1418 44130 1420
rect 44064 1402 44130 1418
rect 45696 1418 45712 1420
rect 45746 1450 45762 1452
rect 47328 1452 47394 1468
rect 47328 1450 47344 1452
rect 45746 1420 47344 1450
rect 45746 1418 45762 1420
rect 45696 1402 45762 1418
rect 47328 1418 47344 1420
rect 47378 1450 47394 1452
rect 48960 1452 49026 1468
rect 48960 1450 48976 1452
rect 47378 1420 48976 1450
rect 47378 1418 47394 1420
rect 47328 1402 47394 1418
rect 48960 1418 48976 1420
rect 49010 1450 49026 1452
rect 50592 1452 50658 1468
rect 50592 1450 50608 1452
rect 49010 1420 50608 1450
rect 49010 1418 49026 1420
rect 48960 1402 49026 1418
rect 50592 1418 50608 1420
rect 50642 1450 50658 1452
rect 52224 1452 52290 1468
rect 52224 1450 52240 1452
rect 50642 1420 52240 1450
rect 50642 1418 50658 1420
rect 50592 1402 50658 1418
rect 52224 1418 52240 1420
rect 52274 1418 52290 1452
rect 52224 1402 52290 1418
rect 0 1248 66 1264
rect 0 1214 16 1248
rect 50 1246 66 1248
rect 1632 1248 1698 1264
rect 1632 1246 1648 1248
rect 50 1216 1648 1246
rect 50 1214 66 1216
rect 0 1198 66 1214
rect 1632 1214 1648 1216
rect 1682 1246 1698 1248
rect 3264 1248 3330 1264
rect 3264 1246 3280 1248
rect 1682 1216 3280 1246
rect 1682 1214 1698 1216
rect 1632 1198 1698 1214
rect 3264 1214 3280 1216
rect 3314 1246 3330 1248
rect 4896 1248 4962 1264
rect 4896 1246 4912 1248
rect 3314 1216 4912 1246
rect 3314 1214 3330 1216
rect 3264 1198 3330 1214
rect 4896 1214 4912 1216
rect 4946 1246 4962 1248
rect 6528 1248 6594 1264
rect 6528 1246 6544 1248
rect 4946 1216 6544 1246
rect 4946 1214 4962 1216
rect 4896 1198 4962 1214
rect 6528 1214 6544 1216
rect 6578 1246 6594 1248
rect 8160 1248 8226 1264
rect 8160 1246 8176 1248
rect 6578 1216 8176 1246
rect 6578 1214 6594 1216
rect 6528 1198 6594 1214
rect 8160 1214 8176 1216
rect 8210 1246 8226 1248
rect 9792 1248 9858 1264
rect 9792 1246 9808 1248
rect 8210 1216 9808 1246
rect 8210 1214 8226 1216
rect 8160 1198 8226 1214
rect 9792 1214 9808 1216
rect 9842 1246 9858 1248
rect 11424 1248 11490 1264
rect 11424 1246 11440 1248
rect 9842 1216 11440 1246
rect 9842 1214 9858 1216
rect 9792 1198 9858 1214
rect 11424 1214 11440 1216
rect 11474 1246 11490 1248
rect 13056 1248 13122 1264
rect 13056 1246 13072 1248
rect 11474 1216 13072 1246
rect 11474 1214 11490 1216
rect 11424 1198 11490 1214
rect 13056 1214 13072 1216
rect 13106 1246 13122 1248
rect 14688 1248 14754 1264
rect 14688 1246 14704 1248
rect 13106 1216 14704 1246
rect 13106 1214 13122 1216
rect 13056 1198 13122 1214
rect 14688 1214 14704 1216
rect 14738 1246 14754 1248
rect 16320 1248 16386 1264
rect 16320 1246 16336 1248
rect 14738 1216 16336 1246
rect 14738 1214 14754 1216
rect 14688 1198 14754 1214
rect 16320 1214 16336 1216
rect 16370 1246 16386 1248
rect 17952 1248 18018 1264
rect 17952 1246 17968 1248
rect 16370 1216 17968 1246
rect 16370 1214 16386 1216
rect 16320 1198 16386 1214
rect 17952 1214 17968 1216
rect 18002 1246 18018 1248
rect 19584 1248 19650 1264
rect 19584 1246 19600 1248
rect 18002 1216 19600 1246
rect 18002 1214 18018 1216
rect 17952 1198 18018 1214
rect 19584 1214 19600 1216
rect 19634 1246 19650 1248
rect 21216 1248 21282 1264
rect 21216 1246 21232 1248
rect 19634 1216 21232 1246
rect 19634 1214 19650 1216
rect 19584 1198 19650 1214
rect 21216 1214 21232 1216
rect 21266 1246 21282 1248
rect 22848 1248 22914 1264
rect 22848 1246 22864 1248
rect 21266 1216 22864 1246
rect 21266 1214 21282 1216
rect 21216 1198 21282 1214
rect 22848 1214 22864 1216
rect 22898 1246 22914 1248
rect 24480 1248 24546 1264
rect 24480 1246 24496 1248
rect 22898 1216 24496 1246
rect 22898 1214 22914 1216
rect 22848 1198 22914 1214
rect 24480 1214 24496 1216
rect 24530 1246 24546 1248
rect 26112 1248 26178 1264
rect 26112 1246 26128 1248
rect 24530 1216 26128 1246
rect 24530 1214 24546 1216
rect 24480 1198 24546 1214
rect 26112 1214 26128 1216
rect 26162 1246 26178 1248
rect 27744 1248 27810 1264
rect 27744 1246 27760 1248
rect 26162 1216 27760 1246
rect 26162 1214 26178 1216
rect 26112 1198 26178 1214
rect 27744 1214 27760 1216
rect 27794 1246 27810 1248
rect 29376 1248 29442 1264
rect 29376 1246 29392 1248
rect 27794 1216 29392 1246
rect 27794 1214 27810 1216
rect 27744 1198 27810 1214
rect 29376 1214 29392 1216
rect 29426 1246 29442 1248
rect 31008 1248 31074 1264
rect 31008 1246 31024 1248
rect 29426 1216 31024 1246
rect 29426 1214 29442 1216
rect 29376 1198 29442 1214
rect 31008 1214 31024 1216
rect 31058 1246 31074 1248
rect 32640 1248 32706 1264
rect 32640 1246 32656 1248
rect 31058 1216 32656 1246
rect 31058 1214 31074 1216
rect 31008 1198 31074 1214
rect 32640 1214 32656 1216
rect 32690 1246 32706 1248
rect 34272 1248 34338 1264
rect 34272 1246 34288 1248
rect 32690 1216 34288 1246
rect 32690 1214 32706 1216
rect 32640 1198 32706 1214
rect 34272 1214 34288 1216
rect 34322 1246 34338 1248
rect 35904 1248 35970 1264
rect 35904 1246 35920 1248
rect 34322 1216 35920 1246
rect 34322 1214 34338 1216
rect 34272 1198 34338 1214
rect 35904 1214 35920 1216
rect 35954 1246 35970 1248
rect 37536 1248 37602 1264
rect 37536 1246 37552 1248
rect 35954 1216 37552 1246
rect 35954 1214 35970 1216
rect 35904 1198 35970 1214
rect 37536 1214 37552 1216
rect 37586 1246 37602 1248
rect 39168 1248 39234 1264
rect 39168 1246 39184 1248
rect 37586 1216 39184 1246
rect 37586 1214 37602 1216
rect 37536 1198 37602 1214
rect 39168 1214 39184 1216
rect 39218 1246 39234 1248
rect 40800 1248 40866 1264
rect 40800 1246 40816 1248
rect 39218 1216 40816 1246
rect 39218 1214 39234 1216
rect 39168 1198 39234 1214
rect 40800 1214 40816 1216
rect 40850 1246 40866 1248
rect 42432 1248 42498 1264
rect 42432 1246 42448 1248
rect 40850 1216 42448 1246
rect 40850 1214 40866 1216
rect 40800 1198 40866 1214
rect 42432 1214 42448 1216
rect 42482 1246 42498 1248
rect 44064 1248 44130 1264
rect 44064 1246 44080 1248
rect 42482 1216 44080 1246
rect 42482 1214 42498 1216
rect 42432 1198 42498 1214
rect 44064 1214 44080 1216
rect 44114 1246 44130 1248
rect 45696 1248 45762 1264
rect 45696 1246 45712 1248
rect 44114 1216 45712 1246
rect 44114 1214 44130 1216
rect 44064 1198 44130 1214
rect 45696 1214 45712 1216
rect 45746 1246 45762 1248
rect 47328 1248 47394 1264
rect 47328 1246 47344 1248
rect 45746 1216 47344 1246
rect 45746 1214 45762 1216
rect 45696 1198 45762 1214
rect 47328 1214 47344 1216
rect 47378 1246 47394 1248
rect 48960 1248 49026 1264
rect 48960 1246 48976 1248
rect 47378 1216 48976 1246
rect 47378 1214 47394 1216
rect 47328 1198 47394 1214
rect 48960 1214 48976 1216
rect 49010 1246 49026 1248
rect 50592 1248 50658 1264
rect 50592 1246 50608 1248
rect 49010 1216 50608 1246
rect 49010 1214 49026 1216
rect 48960 1198 49026 1214
rect 50592 1214 50608 1216
rect 50642 1246 50658 1248
rect 52224 1248 52290 1264
rect 52224 1246 52240 1248
rect 50642 1216 52240 1246
rect 50642 1214 50658 1216
rect 50592 1198 50658 1214
rect 52224 1214 52240 1216
rect 52274 1214 52290 1248
rect 52224 1198 52290 1214
rect 0 1044 66 1060
rect 0 1010 16 1044
rect 50 1042 66 1044
rect 1632 1044 1698 1060
rect 1632 1042 1648 1044
rect 50 1012 1648 1042
rect 50 1010 66 1012
rect 0 994 66 1010
rect 1632 1010 1648 1012
rect 1682 1042 1698 1044
rect 3264 1044 3330 1060
rect 3264 1042 3280 1044
rect 1682 1012 3280 1042
rect 1682 1010 1698 1012
rect 1632 994 1698 1010
rect 3264 1010 3280 1012
rect 3314 1042 3330 1044
rect 4896 1044 4962 1060
rect 4896 1042 4912 1044
rect 3314 1012 4912 1042
rect 3314 1010 3330 1012
rect 3264 994 3330 1010
rect 4896 1010 4912 1012
rect 4946 1042 4962 1044
rect 6528 1044 6594 1060
rect 6528 1042 6544 1044
rect 4946 1012 6544 1042
rect 4946 1010 4962 1012
rect 4896 994 4962 1010
rect 6528 1010 6544 1012
rect 6578 1042 6594 1044
rect 8160 1044 8226 1060
rect 8160 1042 8176 1044
rect 6578 1012 8176 1042
rect 6578 1010 6594 1012
rect 6528 994 6594 1010
rect 8160 1010 8176 1012
rect 8210 1042 8226 1044
rect 9792 1044 9858 1060
rect 9792 1042 9808 1044
rect 8210 1012 9808 1042
rect 8210 1010 8226 1012
rect 8160 994 8226 1010
rect 9792 1010 9808 1012
rect 9842 1042 9858 1044
rect 11424 1044 11490 1060
rect 11424 1042 11440 1044
rect 9842 1012 11440 1042
rect 9842 1010 9858 1012
rect 9792 994 9858 1010
rect 11424 1010 11440 1012
rect 11474 1042 11490 1044
rect 13056 1044 13122 1060
rect 13056 1042 13072 1044
rect 11474 1012 13072 1042
rect 11474 1010 11490 1012
rect 11424 994 11490 1010
rect 13056 1010 13072 1012
rect 13106 1042 13122 1044
rect 14688 1044 14754 1060
rect 14688 1042 14704 1044
rect 13106 1012 14704 1042
rect 13106 1010 13122 1012
rect 13056 994 13122 1010
rect 14688 1010 14704 1012
rect 14738 1042 14754 1044
rect 16320 1044 16386 1060
rect 16320 1042 16336 1044
rect 14738 1012 16336 1042
rect 14738 1010 14754 1012
rect 14688 994 14754 1010
rect 16320 1010 16336 1012
rect 16370 1042 16386 1044
rect 17952 1044 18018 1060
rect 17952 1042 17968 1044
rect 16370 1012 17968 1042
rect 16370 1010 16386 1012
rect 16320 994 16386 1010
rect 17952 1010 17968 1012
rect 18002 1042 18018 1044
rect 19584 1044 19650 1060
rect 19584 1042 19600 1044
rect 18002 1012 19600 1042
rect 18002 1010 18018 1012
rect 17952 994 18018 1010
rect 19584 1010 19600 1012
rect 19634 1042 19650 1044
rect 21216 1044 21282 1060
rect 21216 1042 21232 1044
rect 19634 1012 21232 1042
rect 19634 1010 19650 1012
rect 19584 994 19650 1010
rect 21216 1010 21232 1012
rect 21266 1042 21282 1044
rect 22848 1044 22914 1060
rect 22848 1042 22864 1044
rect 21266 1012 22864 1042
rect 21266 1010 21282 1012
rect 21216 994 21282 1010
rect 22848 1010 22864 1012
rect 22898 1042 22914 1044
rect 24480 1044 24546 1060
rect 24480 1042 24496 1044
rect 22898 1012 24496 1042
rect 22898 1010 22914 1012
rect 22848 994 22914 1010
rect 24480 1010 24496 1012
rect 24530 1042 24546 1044
rect 26112 1044 26178 1060
rect 26112 1042 26128 1044
rect 24530 1012 26128 1042
rect 24530 1010 24546 1012
rect 24480 994 24546 1010
rect 26112 1010 26128 1012
rect 26162 1042 26178 1044
rect 27744 1044 27810 1060
rect 27744 1042 27760 1044
rect 26162 1012 27760 1042
rect 26162 1010 26178 1012
rect 26112 994 26178 1010
rect 27744 1010 27760 1012
rect 27794 1042 27810 1044
rect 29376 1044 29442 1060
rect 29376 1042 29392 1044
rect 27794 1012 29392 1042
rect 27794 1010 27810 1012
rect 27744 994 27810 1010
rect 29376 1010 29392 1012
rect 29426 1042 29442 1044
rect 31008 1044 31074 1060
rect 31008 1042 31024 1044
rect 29426 1012 31024 1042
rect 29426 1010 29442 1012
rect 29376 994 29442 1010
rect 31008 1010 31024 1012
rect 31058 1042 31074 1044
rect 32640 1044 32706 1060
rect 32640 1042 32656 1044
rect 31058 1012 32656 1042
rect 31058 1010 31074 1012
rect 31008 994 31074 1010
rect 32640 1010 32656 1012
rect 32690 1042 32706 1044
rect 34272 1044 34338 1060
rect 34272 1042 34288 1044
rect 32690 1012 34288 1042
rect 32690 1010 32706 1012
rect 32640 994 32706 1010
rect 34272 1010 34288 1012
rect 34322 1042 34338 1044
rect 35904 1044 35970 1060
rect 35904 1042 35920 1044
rect 34322 1012 35920 1042
rect 34322 1010 34338 1012
rect 34272 994 34338 1010
rect 35904 1010 35920 1012
rect 35954 1042 35970 1044
rect 37536 1044 37602 1060
rect 37536 1042 37552 1044
rect 35954 1012 37552 1042
rect 35954 1010 35970 1012
rect 35904 994 35970 1010
rect 37536 1010 37552 1012
rect 37586 1042 37602 1044
rect 39168 1044 39234 1060
rect 39168 1042 39184 1044
rect 37586 1012 39184 1042
rect 37586 1010 37602 1012
rect 37536 994 37602 1010
rect 39168 1010 39184 1012
rect 39218 1042 39234 1044
rect 40800 1044 40866 1060
rect 40800 1042 40816 1044
rect 39218 1012 40816 1042
rect 39218 1010 39234 1012
rect 39168 994 39234 1010
rect 40800 1010 40816 1012
rect 40850 1042 40866 1044
rect 42432 1044 42498 1060
rect 42432 1042 42448 1044
rect 40850 1012 42448 1042
rect 40850 1010 40866 1012
rect 40800 994 40866 1010
rect 42432 1010 42448 1012
rect 42482 1042 42498 1044
rect 44064 1044 44130 1060
rect 44064 1042 44080 1044
rect 42482 1012 44080 1042
rect 42482 1010 42498 1012
rect 42432 994 42498 1010
rect 44064 1010 44080 1012
rect 44114 1042 44130 1044
rect 45696 1044 45762 1060
rect 45696 1042 45712 1044
rect 44114 1012 45712 1042
rect 44114 1010 44130 1012
rect 44064 994 44130 1010
rect 45696 1010 45712 1012
rect 45746 1042 45762 1044
rect 47328 1044 47394 1060
rect 47328 1042 47344 1044
rect 45746 1012 47344 1042
rect 45746 1010 45762 1012
rect 45696 994 45762 1010
rect 47328 1010 47344 1012
rect 47378 1042 47394 1044
rect 48960 1044 49026 1060
rect 48960 1042 48976 1044
rect 47378 1012 48976 1042
rect 47378 1010 47394 1012
rect 47328 994 47394 1010
rect 48960 1010 48976 1012
rect 49010 1042 49026 1044
rect 50592 1044 50658 1060
rect 50592 1042 50608 1044
rect 49010 1012 50608 1042
rect 49010 1010 49026 1012
rect 48960 994 49026 1010
rect 50592 1010 50608 1012
rect 50642 1042 50658 1044
rect 52224 1044 52290 1060
rect 52224 1042 52240 1044
rect 50642 1012 52240 1042
rect 50642 1010 50658 1012
rect 50592 994 50658 1010
rect 52224 1010 52240 1012
rect 52274 1010 52290 1044
rect 52224 994 52290 1010
<< polycont >>
rect 16 2642 50 2676
rect 1648 2642 1682 2676
rect 3280 2642 3314 2676
rect 4912 2642 4946 2676
rect 6544 2642 6578 2676
rect 8176 2642 8210 2676
rect 9808 2642 9842 2676
rect 11440 2642 11474 2676
rect 13072 2642 13106 2676
rect 14704 2642 14738 2676
rect 16336 2642 16370 2676
rect 17968 2642 18002 2676
rect 19600 2642 19634 2676
rect 21232 2642 21266 2676
rect 22864 2642 22898 2676
rect 24496 2642 24530 2676
rect 26128 2642 26162 2676
rect 27760 2642 27794 2676
rect 29392 2642 29426 2676
rect 31024 2642 31058 2676
rect 32656 2642 32690 2676
rect 34288 2642 34322 2676
rect 35920 2642 35954 2676
rect 37552 2642 37586 2676
rect 39184 2642 39218 2676
rect 40816 2642 40850 2676
rect 42448 2642 42482 2676
rect 44080 2642 44114 2676
rect 45712 2642 45746 2676
rect 47344 2642 47378 2676
rect 48976 2642 49010 2676
rect 50608 2642 50642 2676
rect 52240 2642 52274 2676
rect 16 2438 50 2472
rect 1648 2438 1682 2472
rect 3280 2438 3314 2472
rect 4912 2438 4946 2472
rect 6544 2438 6578 2472
rect 8176 2438 8210 2472
rect 9808 2438 9842 2472
rect 11440 2438 11474 2472
rect 13072 2438 13106 2472
rect 14704 2438 14738 2472
rect 16336 2438 16370 2472
rect 17968 2438 18002 2472
rect 19600 2438 19634 2472
rect 21232 2438 21266 2472
rect 22864 2438 22898 2472
rect 24496 2438 24530 2472
rect 26128 2438 26162 2472
rect 27760 2438 27794 2472
rect 29392 2438 29426 2472
rect 31024 2438 31058 2472
rect 32656 2438 32690 2472
rect 34288 2438 34322 2472
rect 35920 2438 35954 2472
rect 37552 2438 37586 2472
rect 39184 2438 39218 2472
rect 40816 2438 40850 2472
rect 42448 2438 42482 2472
rect 44080 2438 44114 2472
rect 45712 2438 45746 2472
rect 47344 2438 47378 2472
rect 48976 2438 49010 2472
rect 50608 2438 50642 2472
rect 52240 2438 52274 2472
rect 16 2234 50 2268
rect 1648 2234 1682 2268
rect 3280 2234 3314 2268
rect 4912 2234 4946 2268
rect 6544 2234 6578 2268
rect 8176 2234 8210 2268
rect 9808 2234 9842 2268
rect 11440 2234 11474 2268
rect 13072 2234 13106 2268
rect 14704 2234 14738 2268
rect 16336 2234 16370 2268
rect 17968 2234 18002 2268
rect 19600 2234 19634 2268
rect 21232 2234 21266 2268
rect 22864 2234 22898 2268
rect 24496 2234 24530 2268
rect 26128 2234 26162 2268
rect 27760 2234 27794 2268
rect 29392 2234 29426 2268
rect 31024 2234 31058 2268
rect 32656 2234 32690 2268
rect 34288 2234 34322 2268
rect 35920 2234 35954 2268
rect 37552 2234 37586 2268
rect 39184 2234 39218 2268
rect 40816 2234 40850 2268
rect 42448 2234 42482 2268
rect 44080 2234 44114 2268
rect 45712 2234 45746 2268
rect 47344 2234 47378 2268
rect 48976 2234 49010 2268
rect 50608 2234 50642 2268
rect 52240 2234 52274 2268
rect 16 2030 50 2064
rect 1648 2030 1682 2064
rect 3280 2030 3314 2064
rect 4912 2030 4946 2064
rect 6544 2030 6578 2064
rect 8176 2030 8210 2064
rect 9808 2030 9842 2064
rect 11440 2030 11474 2064
rect 13072 2030 13106 2064
rect 14704 2030 14738 2064
rect 16336 2030 16370 2064
rect 17968 2030 18002 2064
rect 19600 2030 19634 2064
rect 21232 2030 21266 2064
rect 22864 2030 22898 2064
rect 24496 2030 24530 2064
rect 26128 2030 26162 2064
rect 27760 2030 27794 2064
rect 29392 2030 29426 2064
rect 31024 2030 31058 2064
rect 32656 2030 32690 2064
rect 34288 2030 34322 2064
rect 35920 2030 35954 2064
rect 37552 2030 37586 2064
rect 39184 2030 39218 2064
rect 40816 2030 40850 2064
rect 42448 2030 42482 2064
rect 44080 2030 44114 2064
rect 45712 2030 45746 2064
rect 47344 2030 47378 2064
rect 48976 2030 49010 2064
rect 50608 2030 50642 2064
rect 52240 2030 52274 2064
rect 16 1826 50 1860
rect 1648 1826 1682 1860
rect 3280 1826 3314 1860
rect 4912 1826 4946 1860
rect 6544 1826 6578 1860
rect 8176 1826 8210 1860
rect 9808 1826 9842 1860
rect 11440 1826 11474 1860
rect 13072 1826 13106 1860
rect 14704 1826 14738 1860
rect 16336 1826 16370 1860
rect 17968 1826 18002 1860
rect 19600 1826 19634 1860
rect 21232 1826 21266 1860
rect 22864 1826 22898 1860
rect 24496 1826 24530 1860
rect 26128 1826 26162 1860
rect 27760 1826 27794 1860
rect 29392 1826 29426 1860
rect 31024 1826 31058 1860
rect 32656 1826 32690 1860
rect 34288 1826 34322 1860
rect 35920 1826 35954 1860
rect 37552 1826 37586 1860
rect 39184 1826 39218 1860
rect 40816 1826 40850 1860
rect 42448 1826 42482 1860
rect 44080 1826 44114 1860
rect 45712 1826 45746 1860
rect 47344 1826 47378 1860
rect 48976 1826 49010 1860
rect 50608 1826 50642 1860
rect 52240 1826 52274 1860
rect 16 1622 50 1656
rect 1648 1622 1682 1656
rect 3280 1622 3314 1656
rect 4912 1622 4946 1656
rect 6544 1622 6578 1656
rect 8176 1622 8210 1656
rect 9808 1622 9842 1656
rect 11440 1622 11474 1656
rect 13072 1622 13106 1656
rect 14704 1622 14738 1656
rect 16336 1622 16370 1656
rect 17968 1622 18002 1656
rect 19600 1622 19634 1656
rect 21232 1622 21266 1656
rect 22864 1622 22898 1656
rect 24496 1622 24530 1656
rect 26128 1622 26162 1656
rect 27760 1622 27794 1656
rect 29392 1622 29426 1656
rect 31024 1622 31058 1656
rect 32656 1622 32690 1656
rect 34288 1622 34322 1656
rect 35920 1622 35954 1656
rect 37552 1622 37586 1656
rect 39184 1622 39218 1656
rect 40816 1622 40850 1656
rect 42448 1622 42482 1656
rect 44080 1622 44114 1656
rect 45712 1622 45746 1656
rect 47344 1622 47378 1656
rect 48976 1622 49010 1656
rect 50608 1622 50642 1656
rect 52240 1622 52274 1656
rect 16 1418 50 1452
rect 1648 1418 1682 1452
rect 3280 1418 3314 1452
rect 4912 1418 4946 1452
rect 6544 1418 6578 1452
rect 8176 1418 8210 1452
rect 9808 1418 9842 1452
rect 11440 1418 11474 1452
rect 13072 1418 13106 1452
rect 14704 1418 14738 1452
rect 16336 1418 16370 1452
rect 17968 1418 18002 1452
rect 19600 1418 19634 1452
rect 21232 1418 21266 1452
rect 22864 1418 22898 1452
rect 24496 1418 24530 1452
rect 26128 1418 26162 1452
rect 27760 1418 27794 1452
rect 29392 1418 29426 1452
rect 31024 1418 31058 1452
rect 32656 1418 32690 1452
rect 34288 1418 34322 1452
rect 35920 1418 35954 1452
rect 37552 1418 37586 1452
rect 39184 1418 39218 1452
rect 40816 1418 40850 1452
rect 42448 1418 42482 1452
rect 44080 1418 44114 1452
rect 45712 1418 45746 1452
rect 47344 1418 47378 1452
rect 48976 1418 49010 1452
rect 50608 1418 50642 1452
rect 52240 1418 52274 1452
rect 16 1214 50 1248
rect 1648 1214 1682 1248
rect 3280 1214 3314 1248
rect 4912 1214 4946 1248
rect 6544 1214 6578 1248
rect 8176 1214 8210 1248
rect 9808 1214 9842 1248
rect 11440 1214 11474 1248
rect 13072 1214 13106 1248
rect 14704 1214 14738 1248
rect 16336 1214 16370 1248
rect 17968 1214 18002 1248
rect 19600 1214 19634 1248
rect 21232 1214 21266 1248
rect 22864 1214 22898 1248
rect 24496 1214 24530 1248
rect 26128 1214 26162 1248
rect 27760 1214 27794 1248
rect 29392 1214 29426 1248
rect 31024 1214 31058 1248
rect 32656 1214 32690 1248
rect 34288 1214 34322 1248
rect 35920 1214 35954 1248
rect 37552 1214 37586 1248
rect 39184 1214 39218 1248
rect 40816 1214 40850 1248
rect 42448 1214 42482 1248
rect 44080 1214 44114 1248
rect 45712 1214 45746 1248
rect 47344 1214 47378 1248
rect 48976 1214 49010 1248
rect 50608 1214 50642 1248
rect 52240 1214 52274 1248
rect 16 1010 50 1044
rect 1648 1010 1682 1044
rect 3280 1010 3314 1044
rect 4912 1010 4946 1044
rect 6544 1010 6578 1044
rect 8176 1010 8210 1044
rect 9808 1010 9842 1044
rect 11440 1010 11474 1044
rect 13072 1010 13106 1044
rect 14704 1010 14738 1044
rect 16336 1010 16370 1044
rect 17968 1010 18002 1044
rect 19600 1010 19634 1044
rect 21232 1010 21266 1044
rect 22864 1010 22898 1044
rect 24496 1010 24530 1044
rect 26128 1010 26162 1044
rect 27760 1010 27794 1044
rect 29392 1010 29426 1044
rect 31024 1010 31058 1044
rect 32656 1010 32690 1044
rect 34288 1010 34322 1044
rect 35920 1010 35954 1044
rect 37552 1010 37586 1044
rect 39184 1010 39218 1044
rect 40816 1010 40850 1044
rect 42448 1010 42482 1044
rect 44080 1010 44114 1044
rect 45712 1010 45746 1044
rect 47344 1010 47378 1044
rect 48976 1010 49010 1044
rect 50608 1010 50642 1044
rect 52240 1010 52274 1044
<< locali >>
rect 16 2676 50 2692
rect 16 2626 50 2642
rect 1648 2676 1682 2692
rect 1648 2626 1682 2642
rect 3280 2676 3314 2692
rect 3280 2626 3314 2642
rect 4912 2676 4946 2692
rect 4912 2626 4946 2642
rect 6544 2676 6578 2692
rect 6544 2626 6578 2642
rect 8176 2676 8210 2692
rect 8176 2626 8210 2642
rect 9808 2676 9842 2692
rect 9808 2626 9842 2642
rect 11440 2676 11474 2692
rect 11440 2626 11474 2642
rect 13072 2676 13106 2692
rect 13072 2626 13106 2642
rect 14704 2676 14738 2692
rect 14704 2626 14738 2642
rect 16336 2676 16370 2692
rect 16336 2626 16370 2642
rect 17968 2676 18002 2692
rect 17968 2626 18002 2642
rect 19600 2676 19634 2692
rect 19600 2626 19634 2642
rect 21232 2676 21266 2692
rect 21232 2626 21266 2642
rect 22864 2676 22898 2692
rect 22864 2626 22898 2642
rect 24496 2676 24530 2692
rect 24496 2626 24530 2642
rect 26128 2676 26162 2692
rect 26128 2626 26162 2642
rect 27760 2676 27794 2692
rect 27760 2626 27794 2642
rect 29392 2676 29426 2692
rect 29392 2626 29426 2642
rect 31024 2676 31058 2692
rect 31024 2626 31058 2642
rect 32656 2676 32690 2692
rect 32656 2626 32690 2642
rect 34288 2676 34322 2692
rect 34288 2626 34322 2642
rect 35920 2676 35954 2692
rect 35920 2626 35954 2642
rect 37552 2676 37586 2692
rect 37552 2626 37586 2642
rect 39184 2676 39218 2692
rect 39184 2626 39218 2642
rect 40816 2676 40850 2692
rect 40816 2626 40850 2642
rect 42448 2676 42482 2692
rect 42448 2626 42482 2642
rect 44080 2676 44114 2692
rect 44080 2626 44114 2642
rect 45712 2676 45746 2692
rect 45712 2626 45746 2642
rect 47344 2676 47378 2692
rect 47344 2626 47378 2642
rect 48976 2676 49010 2692
rect 48976 2626 49010 2642
rect 50608 2676 50642 2692
rect 50608 2626 50642 2642
rect 52240 2676 52274 2692
rect 52240 2626 52274 2642
rect 16 2472 50 2488
rect 16 2422 50 2438
rect 1648 2472 1682 2488
rect 1648 2422 1682 2438
rect 3280 2472 3314 2488
rect 3280 2422 3314 2438
rect 4912 2472 4946 2488
rect 4912 2422 4946 2438
rect 6544 2472 6578 2488
rect 6544 2422 6578 2438
rect 8176 2472 8210 2488
rect 8176 2422 8210 2438
rect 9808 2472 9842 2488
rect 9808 2422 9842 2438
rect 11440 2472 11474 2488
rect 11440 2422 11474 2438
rect 13072 2472 13106 2488
rect 13072 2422 13106 2438
rect 14704 2472 14738 2488
rect 14704 2422 14738 2438
rect 16336 2472 16370 2488
rect 16336 2422 16370 2438
rect 17968 2472 18002 2488
rect 17968 2422 18002 2438
rect 19600 2472 19634 2488
rect 19600 2422 19634 2438
rect 21232 2472 21266 2488
rect 21232 2422 21266 2438
rect 22864 2472 22898 2488
rect 22864 2422 22898 2438
rect 24496 2472 24530 2488
rect 24496 2422 24530 2438
rect 26128 2472 26162 2488
rect 26128 2422 26162 2438
rect 27760 2472 27794 2488
rect 27760 2422 27794 2438
rect 29392 2472 29426 2488
rect 29392 2422 29426 2438
rect 31024 2472 31058 2488
rect 31024 2422 31058 2438
rect 32656 2472 32690 2488
rect 32656 2422 32690 2438
rect 34288 2472 34322 2488
rect 34288 2422 34322 2438
rect 35920 2472 35954 2488
rect 35920 2422 35954 2438
rect 37552 2472 37586 2488
rect 37552 2422 37586 2438
rect 39184 2472 39218 2488
rect 39184 2422 39218 2438
rect 40816 2472 40850 2488
rect 40816 2422 40850 2438
rect 42448 2472 42482 2488
rect 42448 2422 42482 2438
rect 44080 2472 44114 2488
rect 44080 2422 44114 2438
rect 45712 2472 45746 2488
rect 45712 2422 45746 2438
rect 47344 2472 47378 2488
rect 47344 2422 47378 2438
rect 48976 2472 49010 2488
rect 48976 2422 49010 2438
rect 50608 2472 50642 2488
rect 50608 2422 50642 2438
rect 52240 2472 52274 2488
rect 52240 2422 52274 2438
rect 16 2268 50 2284
rect 16 2218 50 2234
rect 1648 2268 1682 2284
rect 1648 2218 1682 2234
rect 3280 2268 3314 2284
rect 3280 2218 3314 2234
rect 4912 2268 4946 2284
rect 4912 2218 4946 2234
rect 6544 2268 6578 2284
rect 6544 2218 6578 2234
rect 8176 2268 8210 2284
rect 8176 2218 8210 2234
rect 9808 2268 9842 2284
rect 9808 2218 9842 2234
rect 11440 2268 11474 2284
rect 11440 2218 11474 2234
rect 13072 2268 13106 2284
rect 13072 2218 13106 2234
rect 14704 2268 14738 2284
rect 14704 2218 14738 2234
rect 16336 2268 16370 2284
rect 16336 2218 16370 2234
rect 17968 2268 18002 2284
rect 17968 2218 18002 2234
rect 19600 2268 19634 2284
rect 19600 2218 19634 2234
rect 21232 2268 21266 2284
rect 21232 2218 21266 2234
rect 22864 2268 22898 2284
rect 22864 2218 22898 2234
rect 24496 2268 24530 2284
rect 24496 2218 24530 2234
rect 26128 2268 26162 2284
rect 26128 2218 26162 2234
rect 27760 2268 27794 2284
rect 27760 2218 27794 2234
rect 29392 2268 29426 2284
rect 29392 2218 29426 2234
rect 31024 2268 31058 2284
rect 31024 2218 31058 2234
rect 32656 2268 32690 2284
rect 32656 2218 32690 2234
rect 34288 2268 34322 2284
rect 34288 2218 34322 2234
rect 35920 2268 35954 2284
rect 35920 2218 35954 2234
rect 37552 2268 37586 2284
rect 37552 2218 37586 2234
rect 39184 2268 39218 2284
rect 39184 2218 39218 2234
rect 40816 2268 40850 2284
rect 40816 2218 40850 2234
rect 42448 2268 42482 2284
rect 42448 2218 42482 2234
rect 44080 2268 44114 2284
rect 44080 2218 44114 2234
rect 45712 2268 45746 2284
rect 45712 2218 45746 2234
rect 47344 2268 47378 2284
rect 47344 2218 47378 2234
rect 48976 2268 49010 2284
rect 48976 2218 49010 2234
rect 50608 2268 50642 2284
rect 50608 2218 50642 2234
rect 52240 2268 52274 2284
rect 52240 2218 52274 2234
rect 16 2064 50 2080
rect 16 2014 50 2030
rect 1648 2064 1682 2080
rect 1648 2014 1682 2030
rect 3280 2064 3314 2080
rect 3280 2014 3314 2030
rect 4912 2064 4946 2080
rect 4912 2014 4946 2030
rect 6544 2064 6578 2080
rect 6544 2014 6578 2030
rect 8176 2064 8210 2080
rect 8176 2014 8210 2030
rect 9808 2064 9842 2080
rect 9808 2014 9842 2030
rect 11440 2064 11474 2080
rect 11440 2014 11474 2030
rect 13072 2064 13106 2080
rect 13072 2014 13106 2030
rect 14704 2064 14738 2080
rect 14704 2014 14738 2030
rect 16336 2064 16370 2080
rect 16336 2014 16370 2030
rect 17968 2064 18002 2080
rect 17968 2014 18002 2030
rect 19600 2064 19634 2080
rect 19600 2014 19634 2030
rect 21232 2064 21266 2080
rect 21232 2014 21266 2030
rect 22864 2064 22898 2080
rect 22864 2014 22898 2030
rect 24496 2064 24530 2080
rect 24496 2014 24530 2030
rect 26128 2064 26162 2080
rect 26128 2014 26162 2030
rect 27760 2064 27794 2080
rect 27760 2014 27794 2030
rect 29392 2064 29426 2080
rect 29392 2014 29426 2030
rect 31024 2064 31058 2080
rect 31024 2014 31058 2030
rect 32656 2064 32690 2080
rect 32656 2014 32690 2030
rect 34288 2064 34322 2080
rect 34288 2014 34322 2030
rect 35920 2064 35954 2080
rect 35920 2014 35954 2030
rect 37552 2064 37586 2080
rect 37552 2014 37586 2030
rect 39184 2064 39218 2080
rect 39184 2014 39218 2030
rect 40816 2064 40850 2080
rect 40816 2014 40850 2030
rect 42448 2064 42482 2080
rect 42448 2014 42482 2030
rect 44080 2064 44114 2080
rect 44080 2014 44114 2030
rect 45712 2064 45746 2080
rect 45712 2014 45746 2030
rect 47344 2064 47378 2080
rect 47344 2014 47378 2030
rect 48976 2064 49010 2080
rect 48976 2014 49010 2030
rect 50608 2064 50642 2080
rect 50608 2014 50642 2030
rect 52240 2064 52274 2080
rect 52240 2014 52274 2030
rect 16 1860 50 1876
rect 16 1810 50 1826
rect 1648 1860 1682 1876
rect 1648 1810 1682 1826
rect 3280 1860 3314 1876
rect 3280 1810 3314 1826
rect 4912 1860 4946 1876
rect 4912 1810 4946 1826
rect 6544 1860 6578 1876
rect 6544 1810 6578 1826
rect 8176 1860 8210 1876
rect 8176 1810 8210 1826
rect 9808 1860 9842 1876
rect 9808 1810 9842 1826
rect 11440 1860 11474 1876
rect 11440 1810 11474 1826
rect 13072 1860 13106 1876
rect 13072 1810 13106 1826
rect 14704 1860 14738 1876
rect 14704 1810 14738 1826
rect 16336 1860 16370 1876
rect 16336 1810 16370 1826
rect 17968 1860 18002 1876
rect 17968 1810 18002 1826
rect 19600 1860 19634 1876
rect 19600 1810 19634 1826
rect 21232 1860 21266 1876
rect 21232 1810 21266 1826
rect 22864 1860 22898 1876
rect 22864 1810 22898 1826
rect 24496 1860 24530 1876
rect 24496 1810 24530 1826
rect 26128 1860 26162 1876
rect 26128 1810 26162 1826
rect 27760 1860 27794 1876
rect 27760 1810 27794 1826
rect 29392 1860 29426 1876
rect 29392 1810 29426 1826
rect 31024 1860 31058 1876
rect 31024 1810 31058 1826
rect 32656 1860 32690 1876
rect 32656 1810 32690 1826
rect 34288 1860 34322 1876
rect 34288 1810 34322 1826
rect 35920 1860 35954 1876
rect 35920 1810 35954 1826
rect 37552 1860 37586 1876
rect 37552 1810 37586 1826
rect 39184 1860 39218 1876
rect 39184 1810 39218 1826
rect 40816 1860 40850 1876
rect 40816 1810 40850 1826
rect 42448 1860 42482 1876
rect 42448 1810 42482 1826
rect 44080 1860 44114 1876
rect 44080 1810 44114 1826
rect 45712 1860 45746 1876
rect 45712 1810 45746 1826
rect 47344 1860 47378 1876
rect 47344 1810 47378 1826
rect 48976 1860 49010 1876
rect 48976 1810 49010 1826
rect 50608 1860 50642 1876
rect 50608 1810 50642 1826
rect 52240 1860 52274 1876
rect 52240 1810 52274 1826
rect 16 1656 50 1672
rect 16 1606 50 1622
rect 1648 1656 1682 1672
rect 1648 1606 1682 1622
rect 3280 1656 3314 1672
rect 3280 1606 3314 1622
rect 4912 1656 4946 1672
rect 4912 1606 4946 1622
rect 6544 1656 6578 1672
rect 6544 1606 6578 1622
rect 8176 1656 8210 1672
rect 8176 1606 8210 1622
rect 9808 1656 9842 1672
rect 9808 1606 9842 1622
rect 11440 1656 11474 1672
rect 11440 1606 11474 1622
rect 13072 1656 13106 1672
rect 13072 1606 13106 1622
rect 14704 1656 14738 1672
rect 14704 1606 14738 1622
rect 16336 1656 16370 1672
rect 16336 1606 16370 1622
rect 17968 1656 18002 1672
rect 17968 1606 18002 1622
rect 19600 1656 19634 1672
rect 19600 1606 19634 1622
rect 21232 1656 21266 1672
rect 21232 1606 21266 1622
rect 22864 1656 22898 1672
rect 22864 1606 22898 1622
rect 24496 1656 24530 1672
rect 24496 1606 24530 1622
rect 26128 1656 26162 1672
rect 26128 1606 26162 1622
rect 27760 1656 27794 1672
rect 27760 1606 27794 1622
rect 29392 1656 29426 1672
rect 29392 1606 29426 1622
rect 31024 1656 31058 1672
rect 31024 1606 31058 1622
rect 32656 1656 32690 1672
rect 32656 1606 32690 1622
rect 34288 1656 34322 1672
rect 34288 1606 34322 1622
rect 35920 1656 35954 1672
rect 35920 1606 35954 1622
rect 37552 1656 37586 1672
rect 37552 1606 37586 1622
rect 39184 1656 39218 1672
rect 39184 1606 39218 1622
rect 40816 1656 40850 1672
rect 40816 1606 40850 1622
rect 42448 1656 42482 1672
rect 42448 1606 42482 1622
rect 44080 1656 44114 1672
rect 44080 1606 44114 1622
rect 45712 1656 45746 1672
rect 45712 1606 45746 1622
rect 47344 1656 47378 1672
rect 47344 1606 47378 1622
rect 48976 1656 49010 1672
rect 48976 1606 49010 1622
rect 50608 1656 50642 1672
rect 50608 1606 50642 1622
rect 52240 1656 52274 1672
rect 52240 1606 52274 1622
rect 16 1452 50 1468
rect 16 1402 50 1418
rect 1648 1452 1682 1468
rect 1648 1402 1682 1418
rect 3280 1452 3314 1468
rect 3280 1402 3314 1418
rect 4912 1452 4946 1468
rect 4912 1402 4946 1418
rect 6544 1452 6578 1468
rect 6544 1402 6578 1418
rect 8176 1452 8210 1468
rect 8176 1402 8210 1418
rect 9808 1452 9842 1468
rect 9808 1402 9842 1418
rect 11440 1452 11474 1468
rect 11440 1402 11474 1418
rect 13072 1452 13106 1468
rect 13072 1402 13106 1418
rect 14704 1452 14738 1468
rect 14704 1402 14738 1418
rect 16336 1452 16370 1468
rect 16336 1402 16370 1418
rect 17968 1452 18002 1468
rect 17968 1402 18002 1418
rect 19600 1452 19634 1468
rect 19600 1402 19634 1418
rect 21232 1452 21266 1468
rect 21232 1402 21266 1418
rect 22864 1452 22898 1468
rect 22864 1402 22898 1418
rect 24496 1452 24530 1468
rect 24496 1402 24530 1418
rect 26128 1452 26162 1468
rect 26128 1402 26162 1418
rect 27760 1452 27794 1468
rect 27760 1402 27794 1418
rect 29392 1452 29426 1468
rect 29392 1402 29426 1418
rect 31024 1452 31058 1468
rect 31024 1402 31058 1418
rect 32656 1452 32690 1468
rect 32656 1402 32690 1418
rect 34288 1452 34322 1468
rect 34288 1402 34322 1418
rect 35920 1452 35954 1468
rect 35920 1402 35954 1418
rect 37552 1452 37586 1468
rect 37552 1402 37586 1418
rect 39184 1452 39218 1468
rect 39184 1402 39218 1418
rect 40816 1452 40850 1468
rect 40816 1402 40850 1418
rect 42448 1452 42482 1468
rect 42448 1402 42482 1418
rect 44080 1452 44114 1468
rect 44080 1402 44114 1418
rect 45712 1452 45746 1468
rect 45712 1402 45746 1418
rect 47344 1452 47378 1468
rect 47344 1402 47378 1418
rect 48976 1452 49010 1468
rect 48976 1402 49010 1418
rect 50608 1452 50642 1468
rect 50608 1402 50642 1418
rect 52240 1452 52274 1468
rect 52240 1402 52274 1418
rect 16 1248 50 1264
rect 16 1198 50 1214
rect 1648 1248 1682 1264
rect 1648 1198 1682 1214
rect 3280 1248 3314 1264
rect 3280 1198 3314 1214
rect 4912 1248 4946 1264
rect 4912 1198 4946 1214
rect 6544 1248 6578 1264
rect 6544 1198 6578 1214
rect 8176 1248 8210 1264
rect 8176 1198 8210 1214
rect 9808 1248 9842 1264
rect 9808 1198 9842 1214
rect 11440 1248 11474 1264
rect 11440 1198 11474 1214
rect 13072 1248 13106 1264
rect 13072 1198 13106 1214
rect 14704 1248 14738 1264
rect 14704 1198 14738 1214
rect 16336 1248 16370 1264
rect 16336 1198 16370 1214
rect 17968 1248 18002 1264
rect 17968 1198 18002 1214
rect 19600 1248 19634 1264
rect 19600 1198 19634 1214
rect 21232 1248 21266 1264
rect 21232 1198 21266 1214
rect 22864 1248 22898 1264
rect 22864 1198 22898 1214
rect 24496 1248 24530 1264
rect 24496 1198 24530 1214
rect 26128 1248 26162 1264
rect 26128 1198 26162 1214
rect 27760 1248 27794 1264
rect 27760 1198 27794 1214
rect 29392 1248 29426 1264
rect 29392 1198 29426 1214
rect 31024 1248 31058 1264
rect 31024 1198 31058 1214
rect 32656 1248 32690 1264
rect 32656 1198 32690 1214
rect 34288 1248 34322 1264
rect 34288 1198 34322 1214
rect 35920 1248 35954 1264
rect 35920 1198 35954 1214
rect 37552 1248 37586 1264
rect 37552 1198 37586 1214
rect 39184 1248 39218 1264
rect 39184 1198 39218 1214
rect 40816 1248 40850 1264
rect 40816 1198 40850 1214
rect 42448 1248 42482 1264
rect 42448 1198 42482 1214
rect 44080 1248 44114 1264
rect 44080 1198 44114 1214
rect 45712 1248 45746 1264
rect 45712 1198 45746 1214
rect 47344 1248 47378 1264
rect 47344 1198 47378 1214
rect 48976 1248 49010 1264
rect 48976 1198 49010 1214
rect 50608 1248 50642 1264
rect 50608 1198 50642 1214
rect 52240 1248 52274 1264
rect 52240 1198 52274 1214
rect 16 1044 50 1060
rect 16 994 50 1010
rect 1648 1044 1682 1060
rect 1648 994 1682 1010
rect 3280 1044 3314 1060
rect 3280 994 3314 1010
rect 4912 1044 4946 1060
rect 4912 994 4946 1010
rect 6544 1044 6578 1060
rect 6544 994 6578 1010
rect 8176 1044 8210 1060
rect 8176 994 8210 1010
rect 9808 1044 9842 1060
rect 9808 994 9842 1010
rect 11440 1044 11474 1060
rect 11440 994 11474 1010
rect 13072 1044 13106 1060
rect 13072 994 13106 1010
rect 14704 1044 14738 1060
rect 14704 994 14738 1010
rect 16336 1044 16370 1060
rect 16336 994 16370 1010
rect 17968 1044 18002 1060
rect 17968 994 18002 1010
rect 19600 1044 19634 1060
rect 19600 994 19634 1010
rect 21232 1044 21266 1060
rect 21232 994 21266 1010
rect 22864 1044 22898 1060
rect 22864 994 22898 1010
rect 24496 1044 24530 1060
rect 24496 994 24530 1010
rect 26128 1044 26162 1060
rect 26128 994 26162 1010
rect 27760 1044 27794 1060
rect 27760 994 27794 1010
rect 29392 1044 29426 1060
rect 29392 994 29426 1010
rect 31024 1044 31058 1060
rect 31024 994 31058 1010
rect 32656 1044 32690 1060
rect 32656 994 32690 1010
rect 34288 1044 34322 1060
rect 34288 994 34322 1010
rect 35920 1044 35954 1060
rect 35920 994 35954 1010
rect 37552 1044 37586 1060
rect 37552 994 37586 1010
rect 39184 1044 39218 1060
rect 39184 994 39218 1010
rect 40816 1044 40850 1060
rect 40816 994 40850 1010
rect 42448 1044 42482 1060
rect 42448 994 42482 1010
rect 44080 1044 44114 1060
rect 44080 994 44114 1010
rect 45712 1044 45746 1060
rect 45712 994 45746 1010
rect 47344 1044 47378 1060
rect 47344 994 47378 1010
rect 48976 1044 49010 1060
rect 48976 994 49010 1010
rect 50608 1044 50642 1060
rect 50608 994 50642 1010
rect 52240 1044 52274 1060
rect 52240 994 52274 1010
rect 211 856 227 890
rect 261 856 277 890
rect 415 856 431 890
rect 465 856 481 890
rect 619 856 635 890
rect 669 856 685 890
rect 823 856 839 890
rect 873 856 889 890
rect 1027 856 1043 890
rect 1077 856 1093 890
rect 1231 856 1247 890
rect 1281 856 1297 890
rect 1435 856 1451 890
rect 1485 856 1501 890
rect 1639 856 1655 890
rect 1689 856 1705 890
rect 1843 856 1859 890
rect 1893 856 1909 890
rect 2047 856 2063 890
rect 2097 856 2113 890
rect 2251 856 2267 890
rect 2301 856 2317 890
rect 2455 856 2471 890
rect 2505 856 2521 890
rect 2659 856 2675 890
rect 2709 856 2725 890
rect 2863 856 2879 890
rect 2913 856 2929 890
rect 3067 856 3083 890
rect 3117 856 3133 890
rect 3271 856 3287 890
rect 3321 856 3337 890
rect 3475 856 3491 890
rect 3525 856 3541 890
rect 3679 856 3695 890
rect 3729 856 3745 890
rect 3883 856 3899 890
rect 3933 856 3949 890
rect 4087 856 4103 890
rect 4137 856 4153 890
rect 4291 856 4307 890
rect 4341 856 4357 890
rect 4495 856 4511 890
rect 4545 856 4561 890
rect 4699 856 4715 890
rect 4749 856 4765 890
rect 4903 856 4919 890
rect 4953 856 4969 890
rect 5107 856 5123 890
rect 5157 856 5173 890
rect 5311 856 5327 890
rect 5361 856 5377 890
rect 5515 856 5531 890
rect 5565 856 5581 890
rect 5719 856 5735 890
rect 5769 856 5785 890
rect 5923 856 5939 890
rect 5973 856 5989 890
rect 6127 856 6143 890
rect 6177 856 6193 890
rect 6331 856 6347 890
rect 6381 856 6397 890
rect 6535 856 6551 890
rect 6585 856 6601 890
rect 6739 856 6755 890
rect 6789 856 6805 890
rect 6943 856 6959 890
rect 6993 856 7009 890
rect 7147 856 7163 890
rect 7197 856 7213 890
rect 7351 856 7367 890
rect 7401 856 7417 890
rect 7555 856 7571 890
rect 7605 856 7621 890
rect 7759 856 7775 890
rect 7809 856 7825 890
rect 7963 856 7979 890
rect 8013 856 8029 890
rect 8167 856 8183 890
rect 8217 856 8233 890
rect 8371 856 8387 890
rect 8421 856 8437 890
rect 8575 856 8591 890
rect 8625 856 8641 890
rect 8779 856 8795 890
rect 8829 856 8845 890
rect 8983 856 8999 890
rect 9033 856 9049 890
rect 9187 856 9203 890
rect 9237 856 9253 890
rect 9391 856 9407 890
rect 9441 856 9457 890
rect 9595 856 9611 890
rect 9645 856 9661 890
rect 9799 856 9815 890
rect 9849 856 9865 890
rect 10003 856 10019 890
rect 10053 856 10069 890
rect 10207 856 10223 890
rect 10257 856 10273 890
rect 10411 856 10427 890
rect 10461 856 10477 890
rect 10615 856 10631 890
rect 10665 856 10681 890
rect 10819 856 10835 890
rect 10869 856 10885 890
rect 11023 856 11039 890
rect 11073 856 11089 890
rect 11227 856 11243 890
rect 11277 856 11293 890
rect 11431 856 11447 890
rect 11481 856 11497 890
rect 11635 856 11651 890
rect 11685 856 11701 890
rect 11839 856 11855 890
rect 11889 856 11905 890
rect 12043 856 12059 890
rect 12093 856 12109 890
rect 12247 856 12263 890
rect 12297 856 12313 890
rect 12451 856 12467 890
rect 12501 856 12517 890
rect 12655 856 12671 890
rect 12705 856 12721 890
rect 12859 856 12875 890
rect 12909 856 12925 890
rect 13063 856 13079 890
rect 13113 856 13129 890
rect 13267 856 13283 890
rect 13317 856 13333 890
rect 13471 856 13487 890
rect 13521 856 13537 890
rect 13675 856 13691 890
rect 13725 856 13741 890
rect 13879 856 13895 890
rect 13929 856 13945 890
rect 14083 856 14099 890
rect 14133 856 14149 890
rect 14287 856 14303 890
rect 14337 856 14353 890
rect 14491 856 14507 890
rect 14541 856 14557 890
rect 14695 856 14711 890
rect 14745 856 14761 890
rect 14899 856 14915 890
rect 14949 856 14965 890
rect 15103 856 15119 890
rect 15153 856 15169 890
rect 15307 856 15323 890
rect 15357 856 15373 890
rect 15511 856 15527 890
rect 15561 856 15577 890
rect 15715 856 15731 890
rect 15765 856 15781 890
rect 15919 856 15935 890
rect 15969 856 15985 890
rect 16123 856 16139 890
rect 16173 856 16189 890
rect 16327 856 16343 890
rect 16377 856 16393 890
rect 16531 856 16547 890
rect 16581 856 16597 890
rect 16735 856 16751 890
rect 16785 856 16801 890
rect 16939 856 16955 890
rect 16989 856 17005 890
rect 17143 856 17159 890
rect 17193 856 17209 890
rect 17347 856 17363 890
rect 17397 856 17413 890
rect 17551 856 17567 890
rect 17601 856 17617 890
rect 17755 856 17771 890
rect 17805 856 17821 890
rect 17959 856 17975 890
rect 18009 856 18025 890
rect 18163 856 18179 890
rect 18213 856 18229 890
rect 18367 856 18383 890
rect 18417 856 18433 890
rect 18571 856 18587 890
rect 18621 856 18637 890
rect 18775 856 18791 890
rect 18825 856 18841 890
rect 18979 856 18995 890
rect 19029 856 19045 890
rect 19183 856 19199 890
rect 19233 856 19249 890
rect 19387 856 19403 890
rect 19437 856 19453 890
rect 19591 856 19607 890
rect 19641 856 19657 890
rect 19795 856 19811 890
rect 19845 856 19861 890
rect 19999 856 20015 890
rect 20049 856 20065 890
rect 20203 856 20219 890
rect 20253 856 20269 890
rect 20407 856 20423 890
rect 20457 856 20473 890
rect 20611 856 20627 890
rect 20661 856 20677 890
rect 20815 856 20831 890
rect 20865 856 20881 890
rect 21019 856 21035 890
rect 21069 856 21085 890
rect 21223 856 21239 890
rect 21273 856 21289 890
rect 21427 856 21443 890
rect 21477 856 21493 890
rect 21631 856 21647 890
rect 21681 856 21697 890
rect 21835 856 21851 890
rect 21885 856 21901 890
rect 22039 856 22055 890
rect 22089 856 22105 890
rect 22243 856 22259 890
rect 22293 856 22309 890
rect 22447 856 22463 890
rect 22497 856 22513 890
rect 22651 856 22667 890
rect 22701 856 22717 890
rect 22855 856 22871 890
rect 22905 856 22921 890
rect 23059 856 23075 890
rect 23109 856 23125 890
rect 23263 856 23279 890
rect 23313 856 23329 890
rect 23467 856 23483 890
rect 23517 856 23533 890
rect 23671 856 23687 890
rect 23721 856 23737 890
rect 23875 856 23891 890
rect 23925 856 23941 890
rect 24079 856 24095 890
rect 24129 856 24145 890
rect 24283 856 24299 890
rect 24333 856 24349 890
rect 24487 856 24503 890
rect 24537 856 24553 890
rect 24691 856 24707 890
rect 24741 856 24757 890
rect 24895 856 24911 890
rect 24945 856 24961 890
rect 25099 856 25115 890
rect 25149 856 25165 890
rect 25303 856 25319 890
rect 25353 856 25369 890
rect 25507 856 25523 890
rect 25557 856 25573 890
rect 25711 856 25727 890
rect 25761 856 25777 890
rect 25915 856 25931 890
rect 25965 856 25981 890
rect 26119 856 26135 890
rect 26169 856 26185 890
rect 26323 856 26339 890
rect 26373 856 26389 890
rect 26527 856 26543 890
rect 26577 856 26593 890
rect 26731 856 26747 890
rect 26781 856 26797 890
rect 26935 856 26951 890
rect 26985 856 27001 890
rect 27139 856 27155 890
rect 27189 856 27205 890
rect 27343 856 27359 890
rect 27393 856 27409 890
rect 27547 856 27563 890
rect 27597 856 27613 890
rect 27751 856 27767 890
rect 27801 856 27817 890
rect 27955 856 27971 890
rect 28005 856 28021 890
rect 28159 856 28175 890
rect 28209 856 28225 890
rect 28363 856 28379 890
rect 28413 856 28429 890
rect 28567 856 28583 890
rect 28617 856 28633 890
rect 28771 856 28787 890
rect 28821 856 28837 890
rect 28975 856 28991 890
rect 29025 856 29041 890
rect 29179 856 29195 890
rect 29229 856 29245 890
rect 29383 856 29399 890
rect 29433 856 29449 890
rect 29587 856 29603 890
rect 29637 856 29653 890
rect 29791 856 29807 890
rect 29841 856 29857 890
rect 29995 856 30011 890
rect 30045 856 30061 890
rect 30199 856 30215 890
rect 30249 856 30265 890
rect 30403 856 30419 890
rect 30453 856 30469 890
rect 30607 856 30623 890
rect 30657 856 30673 890
rect 30811 856 30827 890
rect 30861 856 30877 890
rect 31015 856 31031 890
rect 31065 856 31081 890
rect 31219 856 31235 890
rect 31269 856 31285 890
rect 31423 856 31439 890
rect 31473 856 31489 890
rect 31627 856 31643 890
rect 31677 856 31693 890
rect 31831 856 31847 890
rect 31881 856 31897 890
rect 32035 856 32051 890
rect 32085 856 32101 890
rect 32239 856 32255 890
rect 32289 856 32305 890
rect 32443 856 32459 890
rect 32493 856 32509 890
rect 32647 856 32663 890
rect 32697 856 32713 890
rect 32851 856 32867 890
rect 32901 856 32917 890
rect 33055 856 33071 890
rect 33105 856 33121 890
rect 33259 856 33275 890
rect 33309 856 33325 890
rect 33463 856 33479 890
rect 33513 856 33529 890
rect 33667 856 33683 890
rect 33717 856 33733 890
rect 33871 856 33887 890
rect 33921 856 33937 890
rect 34075 856 34091 890
rect 34125 856 34141 890
rect 34279 856 34295 890
rect 34329 856 34345 890
rect 34483 856 34499 890
rect 34533 856 34549 890
rect 34687 856 34703 890
rect 34737 856 34753 890
rect 34891 856 34907 890
rect 34941 856 34957 890
rect 35095 856 35111 890
rect 35145 856 35161 890
rect 35299 856 35315 890
rect 35349 856 35365 890
rect 35503 856 35519 890
rect 35553 856 35569 890
rect 35707 856 35723 890
rect 35757 856 35773 890
rect 35911 856 35927 890
rect 35961 856 35977 890
rect 36115 856 36131 890
rect 36165 856 36181 890
rect 36319 856 36335 890
rect 36369 856 36385 890
rect 36523 856 36539 890
rect 36573 856 36589 890
rect 36727 856 36743 890
rect 36777 856 36793 890
rect 36931 856 36947 890
rect 36981 856 36997 890
rect 37135 856 37151 890
rect 37185 856 37201 890
rect 37339 856 37355 890
rect 37389 856 37405 890
rect 37543 856 37559 890
rect 37593 856 37609 890
rect 37747 856 37763 890
rect 37797 856 37813 890
rect 37951 856 37967 890
rect 38001 856 38017 890
rect 38155 856 38171 890
rect 38205 856 38221 890
rect 38359 856 38375 890
rect 38409 856 38425 890
rect 38563 856 38579 890
rect 38613 856 38629 890
rect 38767 856 38783 890
rect 38817 856 38833 890
rect 38971 856 38987 890
rect 39021 856 39037 890
rect 39175 856 39191 890
rect 39225 856 39241 890
rect 39379 856 39395 890
rect 39429 856 39445 890
rect 39583 856 39599 890
rect 39633 856 39649 890
rect 39787 856 39803 890
rect 39837 856 39853 890
rect 39991 856 40007 890
rect 40041 856 40057 890
rect 40195 856 40211 890
rect 40245 856 40261 890
rect 40399 856 40415 890
rect 40449 856 40465 890
rect 40603 856 40619 890
rect 40653 856 40669 890
rect 40807 856 40823 890
rect 40857 856 40873 890
rect 41011 856 41027 890
rect 41061 856 41077 890
rect 41215 856 41231 890
rect 41265 856 41281 890
rect 41419 856 41435 890
rect 41469 856 41485 890
rect 41623 856 41639 890
rect 41673 856 41689 890
rect 41827 856 41843 890
rect 41877 856 41893 890
rect 42031 856 42047 890
rect 42081 856 42097 890
rect 42235 856 42251 890
rect 42285 856 42301 890
rect 42439 856 42455 890
rect 42489 856 42505 890
rect 42643 856 42659 890
rect 42693 856 42709 890
rect 42847 856 42863 890
rect 42897 856 42913 890
rect 43051 856 43067 890
rect 43101 856 43117 890
rect 43255 856 43271 890
rect 43305 856 43321 890
rect 43459 856 43475 890
rect 43509 856 43525 890
rect 43663 856 43679 890
rect 43713 856 43729 890
rect 43867 856 43883 890
rect 43917 856 43933 890
rect 44071 856 44087 890
rect 44121 856 44137 890
rect 44275 856 44291 890
rect 44325 856 44341 890
rect 44479 856 44495 890
rect 44529 856 44545 890
rect 44683 856 44699 890
rect 44733 856 44749 890
rect 44887 856 44903 890
rect 44937 856 44953 890
rect 45091 856 45107 890
rect 45141 856 45157 890
rect 45295 856 45311 890
rect 45345 856 45361 890
rect 45499 856 45515 890
rect 45549 856 45565 890
rect 45703 856 45719 890
rect 45753 856 45769 890
rect 45907 856 45923 890
rect 45957 856 45973 890
rect 46111 856 46127 890
rect 46161 856 46177 890
rect 46315 856 46331 890
rect 46365 856 46381 890
rect 46519 856 46535 890
rect 46569 856 46585 890
rect 46723 856 46739 890
rect 46773 856 46789 890
rect 46927 856 46943 890
rect 46977 856 46993 890
rect 47131 856 47147 890
rect 47181 856 47197 890
rect 47335 856 47351 890
rect 47385 856 47401 890
rect 47539 856 47555 890
rect 47589 856 47605 890
rect 47743 856 47759 890
rect 47793 856 47809 890
rect 47947 856 47963 890
rect 47997 856 48013 890
rect 48151 856 48167 890
rect 48201 856 48217 890
rect 48355 856 48371 890
rect 48405 856 48421 890
rect 48559 856 48575 890
rect 48609 856 48625 890
rect 48763 856 48779 890
rect 48813 856 48829 890
rect 48967 856 48983 890
rect 49017 856 49033 890
rect 49171 856 49187 890
rect 49221 856 49237 890
rect 49375 856 49391 890
rect 49425 856 49441 890
rect 49579 856 49595 890
rect 49629 856 49645 890
rect 49783 856 49799 890
rect 49833 856 49849 890
rect 49987 856 50003 890
rect 50037 856 50053 890
rect 50191 856 50207 890
rect 50241 856 50257 890
rect 50395 856 50411 890
rect 50445 856 50461 890
rect 50599 856 50615 890
rect 50649 856 50665 890
rect 50803 856 50819 890
rect 50853 856 50869 890
rect 51007 856 51023 890
rect 51057 856 51073 890
rect 51211 856 51227 890
rect 51261 856 51277 890
rect 51415 856 51431 890
rect 51465 856 51481 890
rect 51619 856 51635 890
rect 51669 856 51685 890
rect 51823 856 51839 890
rect 51873 856 51889 890
rect 52027 856 52043 890
rect 52077 856 52093 890
rect 52245 856 52261 890
rect 52295 856 52311 890
<< viali >>
rect 16 2642 50 2676
rect 1648 2642 1682 2676
rect 3280 2642 3314 2676
rect 4912 2642 4946 2676
rect 6544 2642 6578 2676
rect 8176 2642 8210 2676
rect 9808 2642 9842 2676
rect 11440 2642 11474 2676
rect 13072 2642 13106 2676
rect 14704 2642 14738 2676
rect 16336 2642 16370 2676
rect 17968 2642 18002 2676
rect 19600 2642 19634 2676
rect 21232 2642 21266 2676
rect 22864 2642 22898 2676
rect 24496 2642 24530 2676
rect 26128 2642 26162 2676
rect 27760 2642 27794 2676
rect 29392 2642 29426 2676
rect 31024 2642 31058 2676
rect 32656 2642 32690 2676
rect 34288 2642 34322 2676
rect 35920 2642 35954 2676
rect 37552 2642 37586 2676
rect 39184 2642 39218 2676
rect 40816 2642 40850 2676
rect 42448 2642 42482 2676
rect 44080 2642 44114 2676
rect 45712 2642 45746 2676
rect 47344 2642 47378 2676
rect 48976 2642 49010 2676
rect 50608 2642 50642 2676
rect 52240 2642 52274 2676
rect 16 2438 50 2472
rect 1648 2438 1682 2472
rect 3280 2438 3314 2472
rect 4912 2438 4946 2472
rect 6544 2438 6578 2472
rect 8176 2438 8210 2472
rect 9808 2438 9842 2472
rect 11440 2438 11474 2472
rect 13072 2438 13106 2472
rect 14704 2438 14738 2472
rect 16336 2438 16370 2472
rect 17968 2438 18002 2472
rect 19600 2438 19634 2472
rect 21232 2438 21266 2472
rect 22864 2438 22898 2472
rect 24496 2438 24530 2472
rect 26128 2438 26162 2472
rect 27760 2438 27794 2472
rect 29392 2438 29426 2472
rect 31024 2438 31058 2472
rect 32656 2438 32690 2472
rect 34288 2438 34322 2472
rect 35920 2438 35954 2472
rect 37552 2438 37586 2472
rect 39184 2438 39218 2472
rect 40816 2438 40850 2472
rect 42448 2438 42482 2472
rect 44080 2438 44114 2472
rect 45712 2438 45746 2472
rect 47344 2438 47378 2472
rect 48976 2438 49010 2472
rect 50608 2438 50642 2472
rect 52240 2438 52274 2472
rect 16 2234 50 2268
rect 1648 2234 1682 2268
rect 3280 2234 3314 2268
rect 4912 2234 4946 2268
rect 6544 2234 6578 2268
rect 8176 2234 8210 2268
rect 9808 2234 9842 2268
rect 11440 2234 11474 2268
rect 13072 2234 13106 2268
rect 14704 2234 14738 2268
rect 16336 2234 16370 2268
rect 17968 2234 18002 2268
rect 19600 2234 19634 2268
rect 21232 2234 21266 2268
rect 22864 2234 22898 2268
rect 24496 2234 24530 2268
rect 26128 2234 26162 2268
rect 27760 2234 27794 2268
rect 29392 2234 29426 2268
rect 31024 2234 31058 2268
rect 32656 2234 32690 2268
rect 34288 2234 34322 2268
rect 35920 2234 35954 2268
rect 37552 2234 37586 2268
rect 39184 2234 39218 2268
rect 40816 2234 40850 2268
rect 42448 2234 42482 2268
rect 44080 2234 44114 2268
rect 45712 2234 45746 2268
rect 47344 2234 47378 2268
rect 48976 2234 49010 2268
rect 50608 2234 50642 2268
rect 52240 2234 52274 2268
rect 16 2030 50 2064
rect 1648 2030 1682 2064
rect 3280 2030 3314 2064
rect 4912 2030 4946 2064
rect 6544 2030 6578 2064
rect 8176 2030 8210 2064
rect 9808 2030 9842 2064
rect 11440 2030 11474 2064
rect 13072 2030 13106 2064
rect 14704 2030 14738 2064
rect 16336 2030 16370 2064
rect 17968 2030 18002 2064
rect 19600 2030 19634 2064
rect 21232 2030 21266 2064
rect 22864 2030 22898 2064
rect 24496 2030 24530 2064
rect 26128 2030 26162 2064
rect 27760 2030 27794 2064
rect 29392 2030 29426 2064
rect 31024 2030 31058 2064
rect 32656 2030 32690 2064
rect 34288 2030 34322 2064
rect 35920 2030 35954 2064
rect 37552 2030 37586 2064
rect 39184 2030 39218 2064
rect 40816 2030 40850 2064
rect 42448 2030 42482 2064
rect 44080 2030 44114 2064
rect 45712 2030 45746 2064
rect 47344 2030 47378 2064
rect 48976 2030 49010 2064
rect 50608 2030 50642 2064
rect 52240 2030 52274 2064
rect 16 1826 50 1860
rect 1648 1826 1682 1860
rect 3280 1826 3314 1860
rect 4912 1826 4946 1860
rect 6544 1826 6578 1860
rect 8176 1826 8210 1860
rect 9808 1826 9842 1860
rect 11440 1826 11474 1860
rect 13072 1826 13106 1860
rect 14704 1826 14738 1860
rect 16336 1826 16370 1860
rect 17968 1826 18002 1860
rect 19600 1826 19634 1860
rect 21232 1826 21266 1860
rect 22864 1826 22898 1860
rect 24496 1826 24530 1860
rect 26128 1826 26162 1860
rect 27760 1826 27794 1860
rect 29392 1826 29426 1860
rect 31024 1826 31058 1860
rect 32656 1826 32690 1860
rect 34288 1826 34322 1860
rect 35920 1826 35954 1860
rect 37552 1826 37586 1860
rect 39184 1826 39218 1860
rect 40816 1826 40850 1860
rect 42448 1826 42482 1860
rect 44080 1826 44114 1860
rect 45712 1826 45746 1860
rect 47344 1826 47378 1860
rect 48976 1826 49010 1860
rect 50608 1826 50642 1860
rect 52240 1826 52274 1860
rect 16 1622 50 1656
rect 1648 1622 1682 1656
rect 3280 1622 3314 1656
rect 4912 1622 4946 1656
rect 6544 1622 6578 1656
rect 8176 1622 8210 1656
rect 9808 1622 9842 1656
rect 11440 1622 11474 1656
rect 13072 1622 13106 1656
rect 14704 1622 14738 1656
rect 16336 1622 16370 1656
rect 17968 1622 18002 1656
rect 19600 1622 19634 1656
rect 21232 1622 21266 1656
rect 22864 1622 22898 1656
rect 24496 1622 24530 1656
rect 26128 1622 26162 1656
rect 27760 1622 27794 1656
rect 29392 1622 29426 1656
rect 31024 1622 31058 1656
rect 32656 1622 32690 1656
rect 34288 1622 34322 1656
rect 35920 1622 35954 1656
rect 37552 1622 37586 1656
rect 39184 1622 39218 1656
rect 40816 1622 40850 1656
rect 42448 1622 42482 1656
rect 44080 1622 44114 1656
rect 45712 1622 45746 1656
rect 47344 1622 47378 1656
rect 48976 1622 49010 1656
rect 50608 1622 50642 1656
rect 52240 1622 52274 1656
rect 16 1418 50 1452
rect 1648 1418 1682 1452
rect 3280 1418 3314 1452
rect 4912 1418 4946 1452
rect 6544 1418 6578 1452
rect 8176 1418 8210 1452
rect 9808 1418 9842 1452
rect 11440 1418 11474 1452
rect 13072 1418 13106 1452
rect 14704 1418 14738 1452
rect 16336 1418 16370 1452
rect 17968 1418 18002 1452
rect 19600 1418 19634 1452
rect 21232 1418 21266 1452
rect 22864 1418 22898 1452
rect 24496 1418 24530 1452
rect 26128 1418 26162 1452
rect 27760 1418 27794 1452
rect 29392 1418 29426 1452
rect 31024 1418 31058 1452
rect 32656 1418 32690 1452
rect 34288 1418 34322 1452
rect 35920 1418 35954 1452
rect 37552 1418 37586 1452
rect 39184 1418 39218 1452
rect 40816 1418 40850 1452
rect 42448 1418 42482 1452
rect 44080 1418 44114 1452
rect 45712 1418 45746 1452
rect 47344 1418 47378 1452
rect 48976 1418 49010 1452
rect 50608 1418 50642 1452
rect 52240 1418 52274 1452
rect 16 1214 50 1248
rect 1648 1214 1682 1248
rect 3280 1214 3314 1248
rect 4912 1214 4946 1248
rect 6544 1214 6578 1248
rect 8176 1214 8210 1248
rect 9808 1214 9842 1248
rect 11440 1214 11474 1248
rect 13072 1214 13106 1248
rect 14704 1214 14738 1248
rect 16336 1214 16370 1248
rect 17968 1214 18002 1248
rect 19600 1214 19634 1248
rect 21232 1214 21266 1248
rect 22864 1214 22898 1248
rect 24496 1214 24530 1248
rect 26128 1214 26162 1248
rect 27760 1214 27794 1248
rect 29392 1214 29426 1248
rect 31024 1214 31058 1248
rect 32656 1214 32690 1248
rect 34288 1214 34322 1248
rect 35920 1214 35954 1248
rect 37552 1214 37586 1248
rect 39184 1214 39218 1248
rect 40816 1214 40850 1248
rect 42448 1214 42482 1248
rect 44080 1214 44114 1248
rect 45712 1214 45746 1248
rect 47344 1214 47378 1248
rect 48976 1214 49010 1248
rect 50608 1214 50642 1248
rect 52240 1214 52274 1248
rect 16 1010 50 1044
rect 1648 1010 1682 1044
rect 3280 1010 3314 1044
rect 4912 1010 4946 1044
rect 6544 1010 6578 1044
rect 8176 1010 8210 1044
rect 9808 1010 9842 1044
rect 11440 1010 11474 1044
rect 13072 1010 13106 1044
rect 14704 1010 14738 1044
rect 16336 1010 16370 1044
rect 17968 1010 18002 1044
rect 19600 1010 19634 1044
rect 21232 1010 21266 1044
rect 22864 1010 22898 1044
rect 24496 1010 24530 1044
rect 26128 1010 26162 1044
rect 27760 1010 27794 1044
rect 29392 1010 29426 1044
rect 31024 1010 31058 1044
rect 32656 1010 32690 1044
rect 34288 1010 34322 1044
rect 35920 1010 35954 1044
rect 37552 1010 37586 1044
rect 39184 1010 39218 1044
rect 40816 1010 40850 1044
rect 42448 1010 42482 1044
rect 44080 1010 44114 1044
rect 45712 1010 45746 1044
rect 47344 1010 47378 1044
rect 48976 1010 49010 1044
rect 50608 1010 50642 1044
rect 52240 1010 52274 1044
rect 227 856 261 890
rect 431 856 465 890
rect 635 856 669 890
rect 839 856 873 890
rect 1043 856 1077 890
rect 1247 856 1281 890
rect 1451 856 1485 890
rect 1655 856 1689 890
rect 1859 856 1893 890
rect 2063 856 2097 890
rect 2267 856 2301 890
rect 2471 856 2505 890
rect 2675 856 2709 890
rect 2879 856 2913 890
rect 3083 856 3117 890
rect 3287 856 3321 890
rect 3491 856 3525 890
rect 3695 856 3729 890
rect 3899 856 3933 890
rect 4103 856 4137 890
rect 4307 856 4341 890
rect 4511 856 4545 890
rect 4715 856 4749 890
rect 4919 856 4953 890
rect 5123 856 5157 890
rect 5327 856 5361 890
rect 5531 856 5565 890
rect 5735 856 5769 890
rect 5939 856 5973 890
rect 6143 856 6177 890
rect 6347 856 6381 890
rect 6551 856 6585 890
rect 6755 856 6789 890
rect 6959 856 6993 890
rect 7163 856 7197 890
rect 7367 856 7401 890
rect 7571 856 7605 890
rect 7775 856 7809 890
rect 7979 856 8013 890
rect 8183 856 8217 890
rect 8387 856 8421 890
rect 8591 856 8625 890
rect 8795 856 8829 890
rect 8999 856 9033 890
rect 9203 856 9237 890
rect 9407 856 9441 890
rect 9611 856 9645 890
rect 9815 856 9849 890
rect 10019 856 10053 890
rect 10223 856 10257 890
rect 10427 856 10461 890
rect 10631 856 10665 890
rect 10835 856 10869 890
rect 11039 856 11073 890
rect 11243 856 11277 890
rect 11447 856 11481 890
rect 11651 856 11685 890
rect 11855 856 11889 890
rect 12059 856 12093 890
rect 12263 856 12297 890
rect 12467 856 12501 890
rect 12671 856 12705 890
rect 12875 856 12909 890
rect 13079 856 13113 890
rect 13283 856 13317 890
rect 13487 856 13521 890
rect 13691 856 13725 890
rect 13895 856 13929 890
rect 14099 856 14133 890
rect 14303 856 14337 890
rect 14507 856 14541 890
rect 14711 856 14745 890
rect 14915 856 14949 890
rect 15119 856 15153 890
rect 15323 856 15357 890
rect 15527 856 15561 890
rect 15731 856 15765 890
rect 15935 856 15969 890
rect 16139 856 16173 890
rect 16343 856 16377 890
rect 16547 856 16581 890
rect 16751 856 16785 890
rect 16955 856 16989 890
rect 17159 856 17193 890
rect 17363 856 17397 890
rect 17567 856 17601 890
rect 17771 856 17805 890
rect 17975 856 18009 890
rect 18179 856 18213 890
rect 18383 856 18417 890
rect 18587 856 18621 890
rect 18791 856 18825 890
rect 18995 856 19029 890
rect 19199 856 19233 890
rect 19403 856 19437 890
rect 19607 856 19641 890
rect 19811 856 19845 890
rect 20015 856 20049 890
rect 20219 856 20253 890
rect 20423 856 20457 890
rect 20627 856 20661 890
rect 20831 856 20865 890
rect 21035 856 21069 890
rect 21239 856 21273 890
rect 21443 856 21477 890
rect 21647 856 21681 890
rect 21851 856 21885 890
rect 22055 856 22089 890
rect 22259 856 22293 890
rect 22463 856 22497 890
rect 22667 856 22701 890
rect 22871 856 22905 890
rect 23075 856 23109 890
rect 23279 856 23313 890
rect 23483 856 23517 890
rect 23687 856 23721 890
rect 23891 856 23925 890
rect 24095 856 24129 890
rect 24299 856 24333 890
rect 24503 856 24537 890
rect 24707 856 24741 890
rect 24911 856 24945 890
rect 25115 856 25149 890
rect 25319 856 25353 890
rect 25523 856 25557 890
rect 25727 856 25761 890
rect 25931 856 25965 890
rect 26135 856 26169 890
rect 26339 856 26373 890
rect 26543 856 26577 890
rect 26747 856 26781 890
rect 26951 856 26985 890
rect 27155 856 27189 890
rect 27359 856 27393 890
rect 27563 856 27597 890
rect 27767 856 27801 890
rect 27971 856 28005 890
rect 28175 856 28209 890
rect 28379 856 28413 890
rect 28583 856 28617 890
rect 28787 856 28821 890
rect 28991 856 29025 890
rect 29195 856 29229 890
rect 29399 856 29433 890
rect 29603 856 29637 890
rect 29807 856 29841 890
rect 30011 856 30045 890
rect 30215 856 30249 890
rect 30419 856 30453 890
rect 30623 856 30657 890
rect 30827 856 30861 890
rect 31031 856 31065 890
rect 31235 856 31269 890
rect 31439 856 31473 890
rect 31643 856 31677 890
rect 31847 856 31881 890
rect 32051 856 32085 890
rect 32255 856 32289 890
rect 32459 856 32493 890
rect 32663 856 32697 890
rect 32867 856 32901 890
rect 33071 856 33105 890
rect 33275 856 33309 890
rect 33479 856 33513 890
rect 33683 856 33717 890
rect 33887 856 33921 890
rect 34091 856 34125 890
rect 34295 856 34329 890
rect 34499 856 34533 890
rect 34703 856 34737 890
rect 34907 856 34941 890
rect 35111 856 35145 890
rect 35315 856 35349 890
rect 35519 856 35553 890
rect 35723 856 35757 890
rect 35927 856 35961 890
rect 36131 856 36165 890
rect 36335 856 36369 890
rect 36539 856 36573 890
rect 36743 856 36777 890
rect 36947 856 36981 890
rect 37151 856 37185 890
rect 37355 856 37389 890
rect 37559 856 37593 890
rect 37763 856 37797 890
rect 37967 856 38001 890
rect 38171 856 38205 890
rect 38375 856 38409 890
rect 38579 856 38613 890
rect 38783 856 38817 890
rect 38987 856 39021 890
rect 39191 856 39225 890
rect 39395 856 39429 890
rect 39599 856 39633 890
rect 39803 856 39837 890
rect 40007 856 40041 890
rect 40211 856 40245 890
rect 40415 856 40449 890
rect 40619 856 40653 890
rect 40823 856 40857 890
rect 41027 856 41061 890
rect 41231 856 41265 890
rect 41435 856 41469 890
rect 41639 856 41673 890
rect 41843 856 41877 890
rect 42047 856 42081 890
rect 42251 856 42285 890
rect 42455 856 42489 890
rect 42659 856 42693 890
rect 42863 856 42897 890
rect 43067 856 43101 890
rect 43271 856 43305 890
rect 43475 856 43509 890
rect 43679 856 43713 890
rect 43883 856 43917 890
rect 44087 856 44121 890
rect 44291 856 44325 890
rect 44495 856 44529 890
rect 44699 856 44733 890
rect 44903 856 44937 890
rect 45107 856 45141 890
rect 45311 856 45345 890
rect 45515 856 45549 890
rect 45719 856 45753 890
rect 45923 856 45957 890
rect 46127 856 46161 890
rect 46331 856 46365 890
rect 46535 856 46569 890
rect 46739 856 46773 890
rect 46943 856 46977 890
rect 47147 856 47181 890
rect 47351 856 47385 890
rect 47555 856 47589 890
rect 47759 856 47793 890
rect 47963 856 47997 890
rect 48167 856 48201 890
rect 48371 856 48405 890
rect 48575 856 48609 890
rect 48779 856 48813 890
rect 48983 856 49017 890
rect 49187 856 49221 890
rect 49391 856 49425 890
rect 49595 856 49629 890
rect 49799 856 49833 890
rect 50003 856 50037 890
rect 50207 856 50241 890
rect 50411 856 50445 890
rect 50615 856 50649 890
rect 50819 856 50853 890
rect 51023 856 51057 890
rect 51227 856 51261 890
rect 51431 856 51465 890
rect 51635 856 51669 890
rect 51839 856 51873 890
rect 52043 856 52077 890
rect 52261 856 52295 890
<< metal1 >>
rect 114 2772 52190 2800
rect 8 2685 59 2692
rect 1640 2685 1691 2692
rect 3272 2685 3323 2692
rect 4904 2685 4955 2692
rect 6536 2685 6587 2692
rect 8168 2685 8219 2692
rect 9800 2685 9851 2692
rect 11432 2685 11483 2692
rect 13064 2685 13115 2692
rect 14696 2685 14747 2692
rect 16328 2685 16379 2692
rect 17960 2685 18011 2692
rect 19592 2685 19643 2692
rect 21224 2685 21275 2692
rect 22856 2685 22907 2692
rect 24488 2685 24539 2692
rect 26120 2685 26171 2692
rect 27752 2685 27803 2692
rect 29384 2685 29435 2692
rect 31016 2685 31067 2692
rect 32648 2685 32699 2692
rect 34280 2685 34331 2692
rect 35912 2685 35963 2692
rect 37544 2685 37595 2692
rect 39176 2685 39227 2692
rect 40808 2685 40859 2692
rect 42440 2685 42491 2692
rect 44072 2685 44123 2692
rect 45704 2685 45755 2692
rect 47336 2685 47387 2692
rect 48968 2685 49019 2692
rect 50600 2685 50651 2692
rect 52232 2685 52283 2692
rect 1 2633 7 2685
rect 59 2633 65 2685
rect 1633 2633 1639 2685
rect 1691 2633 1697 2685
rect 3265 2633 3271 2685
rect 3323 2633 3329 2685
rect 4897 2633 4903 2685
rect 4955 2633 4961 2685
rect 6529 2633 6535 2685
rect 6587 2633 6593 2685
rect 8161 2633 8167 2685
rect 8219 2633 8225 2685
rect 9793 2633 9799 2685
rect 9851 2633 9857 2685
rect 11425 2633 11431 2685
rect 11483 2633 11489 2685
rect 13057 2633 13063 2685
rect 13115 2633 13121 2685
rect 14689 2633 14695 2685
rect 14747 2633 14753 2685
rect 16321 2633 16327 2685
rect 16379 2633 16385 2685
rect 17953 2633 17959 2685
rect 18011 2633 18017 2685
rect 19585 2633 19591 2685
rect 19643 2633 19649 2685
rect 21217 2633 21223 2685
rect 21275 2633 21281 2685
rect 22849 2633 22855 2685
rect 22907 2633 22913 2685
rect 24481 2633 24487 2685
rect 24539 2633 24545 2685
rect 26113 2633 26119 2685
rect 26171 2633 26177 2685
rect 27745 2633 27751 2685
rect 27803 2633 27809 2685
rect 29377 2633 29383 2685
rect 29435 2633 29441 2685
rect 31009 2633 31015 2685
rect 31067 2633 31073 2685
rect 32641 2633 32647 2685
rect 32699 2633 32705 2685
rect 34273 2633 34279 2685
rect 34331 2633 34337 2685
rect 35905 2633 35911 2685
rect 35963 2633 35969 2685
rect 37537 2633 37543 2685
rect 37595 2633 37601 2685
rect 39169 2633 39175 2685
rect 39227 2633 39233 2685
rect 40801 2633 40807 2685
rect 40859 2633 40865 2685
rect 42433 2633 42439 2685
rect 42491 2633 42497 2685
rect 44065 2633 44071 2685
rect 44123 2633 44129 2685
rect 45697 2633 45703 2685
rect 45755 2633 45761 2685
rect 47329 2633 47335 2685
rect 47387 2633 47393 2685
rect 48961 2633 48967 2685
rect 49019 2633 49025 2685
rect 50593 2633 50599 2685
rect 50651 2633 50657 2685
rect 52225 2633 52231 2685
rect 52283 2673 52289 2685
rect 52283 2645 52473 2673
rect 52283 2633 52289 2645
rect 8 2626 59 2633
rect 1640 2626 1691 2633
rect 3272 2626 3323 2633
rect 4904 2626 4955 2633
rect 6536 2626 6587 2633
rect 8168 2626 8219 2633
rect 9800 2626 9851 2633
rect 11432 2626 11483 2633
rect 13064 2626 13115 2633
rect 14696 2626 14747 2633
rect 16328 2626 16379 2633
rect 17960 2626 18011 2633
rect 19592 2626 19643 2633
rect 21224 2626 21275 2633
rect 22856 2626 22907 2633
rect 24488 2626 24539 2633
rect 26120 2626 26171 2633
rect 27752 2626 27803 2633
rect 29384 2626 29435 2633
rect 31016 2626 31067 2633
rect 32648 2626 32699 2633
rect 34280 2626 34331 2633
rect 35912 2626 35963 2633
rect 37544 2626 37595 2633
rect 39176 2626 39227 2633
rect 40808 2626 40859 2633
rect 42440 2626 42491 2633
rect 44072 2626 44123 2633
rect 45704 2626 45755 2633
rect 47336 2626 47387 2633
rect 48968 2626 49019 2633
rect 50600 2626 50651 2633
rect 52232 2626 52283 2633
rect 8 2481 59 2488
rect 1640 2481 1691 2488
rect 3272 2481 3323 2488
rect 4904 2481 4955 2488
rect 6536 2481 6587 2488
rect 8168 2481 8219 2488
rect 9800 2481 9851 2488
rect 11432 2481 11483 2488
rect 13064 2481 13115 2488
rect 14696 2481 14747 2488
rect 16328 2481 16379 2488
rect 17960 2481 18011 2488
rect 19592 2481 19643 2488
rect 21224 2481 21275 2488
rect 22856 2481 22907 2488
rect 24488 2481 24539 2488
rect 26120 2481 26171 2488
rect 27752 2481 27803 2488
rect 29384 2481 29435 2488
rect 31016 2481 31067 2488
rect 32648 2481 32699 2488
rect 34280 2481 34331 2488
rect 35912 2481 35963 2488
rect 37544 2481 37595 2488
rect 39176 2481 39227 2488
rect 40808 2481 40859 2488
rect 42440 2481 42491 2488
rect 44072 2481 44123 2488
rect 45704 2481 45755 2488
rect 47336 2481 47387 2488
rect 48968 2481 49019 2488
rect 50600 2481 50651 2488
rect 52232 2481 52283 2488
rect 1 2429 7 2481
rect 59 2429 65 2481
rect 1633 2429 1639 2481
rect 1691 2429 1697 2481
rect 3265 2429 3271 2481
rect 3323 2429 3329 2481
rect 4897 2429 4903 2481
rect 4955 2429 4961 2481
rect 6529 2429 6535 2481
rect 6587 2429 6593 2481
rect 8161 2429 8167 2481
rect 8219 2429 8225 2481
rect 9793 2429 9799 2481
rect 9851 2429 9857 2481
rect 11425 2429 11431 2481
rect 11483 2429 11489 2481
rect 13057 2429 13063 2481
rect 13115 2429 13121 2481
rect 14689 2429 14695 2481
rect 14747 2429 14753 2481
rect 16321 2429 16327 2481
rect 16379 2429 16385 2481
rect 17953 2429 17959 2481
rect 18011 2429 18017 2481
rect 19585 2429 19591 2481
rect 19643 2429 19649 2481
rect 21217 2429 21223 2481
rect 21275 2429 21281 2481
rect 22849 2429 22855 2481
rect 22907 2429 22913 2481
rect 24481 2429 24487 2481
rect 24539 2429 24545 2481
rect 26113 2429 26119 2481
rect 26171 2429 26177 2481
rect 27745 2429 27751 2481
rect 27803 2429 27809 2481
rect 29377 2429 29383 2481
rect 29435 2429 29441 2481
rect 31009 2429 31015 2481
rect 31067 2429 31073 2481
rect 32641 2429 32647 2481
rect 32699 2429 32705 2481
rect 34273 2429 34279 2481
rect 34331 2429 34337 2481
rect 35905 2429 35911 2481
rect 35963 2429 35969 2481
rect 37537 2429 37543 2481
rect 37595 2429 37601 2481
rect 39169 2429 39175 2481
rect 39227 2429 39233 2481
rect 40801 2429 40807 2481
rect 40859 2429 40865 2481
rect 42433 2429 42439 2481
rect 42491 2429 42497 2481
rect 44065 2429 44071 2481
rect 44123 2429 44129 2481
rect 45697 2429 45703 2481
rect 45755 2429 45761 2481
rect 47329 2429 47335 2481
rect 47387 2429 47393 2481
rect 48961 2429 48967 2481
rect 49019 2429 49025 2481
rect 50593 2429 50599 2481
rect 50651 2429 50657 2481
rect 52225 2429 52231 2481
rect 52283 2429 52289 2481
rect 8 2422 59 2429
rect 1640 2422 1691 2429
rect 3272 2422 3323 2429
rect 4904 2422 4955 2429
rect 6536 2422 6587 2429
rect 8168 2422 8219 2429
rect 9800 2422 9851 2429
rect 11432 2422 11483 2429
rect 13064 2422 13115 2429
rect 14696 2422 14747 2429
rect 16328 2422 16379 2429
rect 17960 2422 18011 2429
rect 19592 2422 19643 2429
rect 21224 2422 21275 2429
rect 22856 2422 22907 2429
rect 24488 2422 24539 2429
rect 26120 2422 26171 2429
rect 27752 2422 27803 2429
rect 29384 2422 29435 2429
rect 31016 2422 31067 2429
rect 32648 2422 32699 2429
rect 34280 2422 34331 2429
rect 35912 2422 35963 2429
rect 37544 2422 37595 2429
rect 39176 2422 39227 2429
rect 40808 2422 40859 2429
rect 42440 2422 42491 2429
rect 44072 2422 44123 2429
rect 45704 2422 45755 2429
rect 47336 2422 47387 2429
rect 48968 2422 49019 2429
rect 50600 2422 50651 2429
rect 52232 2422 52283 2429
rect 8 2277 59 2284
rect 1640 2277 1691 2284
rect 3272 2277 3323 2284
rect 4904 2277 4955 2284
rect 6536 2277 6587 2284
rect 8168 2277 8219 2284
rect 9800 2277 9851 2284
rect 11432 2277 11483 2284
rect 13064 2277 13115 2284
rect 14696 2277 14747 2284
rect 16328 2277 16379 2284
rect 17960 2277 18011 2284
rect 19592 2277 19643 2284
rect 21224 2277 21275 2284
rect 22856 2277 22907 2284
rect 24488 2277 24539 2284
rect 26120 2277 26171 2284
rect 27752 2277 27803 2284
rect 29384 2277 29435 2284
rect 31016 2277 31067 2284
rect 32648 2277 32699 2284
rect 34280 2277 34331 2284
rect 35912 2277 35963 2284
rect 37544 2277 37595 2284
rect 39176 2277 39227 2284
rect 40808 2277 40859 2284
rect 42440 2277 42491 2284
rect 44072 2277 44123 2284
rect 45704 2277 45755 2284
rect 47336 2277 47387 2284
rect 48968 2277 49019 2284
rect 50600 2277 50651 2284
rect 52232 2277 52283 2284
rect 1 2225 7 2277
rect 59 2225 65 2277
rect 1633 2225 1639 2277
rect 1691 2225 1697 2277
rect 3265 2225 3271 2277
rect 3323 2225 3329 2277
rect 4897 2225 4903 2277
rect 4955 2225 4961 2277
rect 6529 2225 6535 2277
rect 6587 2225 6593 2277
rect 8161 2225 8167 2277
rect 8219 2225 8225 2277
rect 9793 2225 9799 2277
rect 9851 2225 9857 2277
rect 11425 2225 11431 2277
rect 11483 2225 11489 2277
rect 13057 2225 13063 2277
rect 13115 2225 13121 2277
rect 14689 2225 14695 2277
rect 14747 2225 14753 2277
rect 16321 2225 16327 2277
rect 16379 2225 16385 2277
rect 17953 2225 17959 2277
rect 18011 2225 18017 2277
rect 19585 2225 19591 2277
rect 19643 2225 19649 2277
rect 21217 2225 21223 2277
rect 21275 2225 21281 2277
rect 22849 2225 22855 2277
rect 22907 2225 22913 2277
rect 24481 2225 24487 2277
rect 24539 2225 24545 2277
rect 26113 2225 26119 2277
rect 26171 2225 26177 2277
rect 27745 2225 27751 2277
rect 27803 2225 27809 2277
rect 29377 2225 29383 2277
rect 29435 2225 29441 2277
rect 31009 2225 31015 2277
rect 31067 2225 31073 2277
rect 32641 2225 32647 2277
rect 32699 2225 32705 2277
rect 34273 2225 34279 2277
rect 34331 2225 34337 2277
rect 35905 2225 35911 2277
rect 35963 2225 35969 2277
rect 37537 2225 37543 2277
rect 37595 2225 37601 2277
rect 39169 2225 39175 2277
rect 39227 2225 39233 2277
rect 40801 2225 40807 2277
rect 40859 2225 40865 2277
rect 42433 2225 42439 2277
rect 42491 2225 42497 2277
rect 44065 2225 44071 2277
rect 44123 2225 44129 2277
rect 45697 2225 45703 2277
rect 45755 2225 45761 2277
rect 47329 2225 47335 2277
rect 47387 2225 47393 2277
rect 48961 2225 48967 2277
rect 49019 2225 49025 2277
rect 50593 2225 50599 2277
rect 50651 2225 50657 2277
rect 52225 2225 52231 2277
rect 52283 2225 52289 2277
rect 8 2218 59 2225
rect 1640 2218 1691 2225
rect 3272 2218 3323 2225
rect 4904 2218 4955 2225
rect 6536 2218 6587 2225
rect 8168 2218 8219 2225
rect 9800 2218 9851 2225
rect 11432 2218 11483 2225
rect 13064 2218 13115 2225
rect 14696 2218 14747 2225
rect 16328 2218 16379 2225
rect 17960 2218 18011 2225
rect 19592 2218 19643 2225
rect 21224 2218 21275 2225
rect 22856 2218 22907 2225
rect 24488 2218 24539 2225
rect 26120 2218 26171 2225
rect 27752 2218 27803 2225
rect 29384 2218 29435 2225
rect 31016 2218 31067 2225
rect 32648 2218 32699 2225
rect 34280 2218 34331 2225
rect 35912 2218 35963 2225
rect 37544 2218 37595 2225
rect 39176 2218 39227 2225
rect 40808 2218 40859 2225
rect 42440 2218 42491 2225
rect 44072 2218 44123 2225
rect 45704 2218 45755 2225
rect 47336 2218 47387 2225
rect 48968 2218 49019 2225
rect 50600 2218 50651 2225
rect 52232 2218 52283 2225
rect 8 2073 59 2080
rect 1640 2073 1691 2080
rect 3272 2073 3323 2080
rect 4904 2073 4955 2080
rect 6536 2073 6587 2080
rect 8168 2073 8219 2080
rect 9800 2073 9851 2080
rect 11432 2073 11483 2080
rect 13064 2073 13115 2080
rect 14696 2073 14747 2080
rect 16328 2073 16379 2080
rect 17960 2073 18011 2080
rect 19592 2073 19643 2080
rect 21224 2073 21275 2080
rect 22856 2073 22907 2080
rect 24488 2073 24539 2080
rect 26120 2073 26171 2080
rect 27752 2073 27803 2080
rect 29384 2073 29435 2080
rect 31016 2073 31067 2080
rect 32648 2073 32699 2080
rect 34280 2073 34331 2080
rect 35912 2073 35963 2080
rect 37544 2073 37595 2080
rect 39176 2073 39227 2080
rect 40808 2073 40859 2080
rect 42440 2073 42491 2080
rect 44072 2073 44123 2080
rect 45704 2073 45755 2080
rect 47336 2073 47387 2080
rect 48968 2073 49019 2080
rect 50600 2073 50651 2080
rect 52232 2073 52283 2080
rect 1 2021 7 2073
rect 59 2021 65 2073
rect 1633 2021 1639 2073
rect 1691 2021 1697 2073
rect 3265 2021 3271 2073
rect 3323 2021 3329 2073
rect 4897 2021 4903 2073
rect 4955 2021 4961 2073
rect 6529 2021 6535 2073
rect 6587 2021 6593 2073
rect 8161 2021 8167 2073
rect 8219 2021 8225 2073
rect 9793 2021 9799 2073
rect 9851 2021 9857 2073
rect 11425 2021 11431 2073
rect 11483 2021 11489 2073
rect 13057 2021 13063 2073
rect 13115 2021 13121 2073
rect 14689 2021 14695 2073
rect 14747 2021 14753 2073
rect 16321 2021 16327 2073
rect 16379 2021 16385 2073
rect 17953 2021 17959 2073
rect 18011 2021 18017 2073
rect 19585 2021 19591 2073
rect 19643 2021 19649 2073
rect 21217 2021 21223 2073
rect 21275 2021 21281 2073
rect 22849 2021 22855 2073
rect 22907 2021 22913 2073
rect 24481 2021 24487 2073
rect 24539 2021 24545 2073
rect 26113 2021 26119 2073
rect 26171 2021 26177 2073
rect 27745 2021 27751 2073
rect 27803 2021 27809 2073
rect 29377 2021 29383 2073
rect 29435 2021 29441 2073
rect 31009 2021 31015 2073
rect 31067 2021 31073 2073
rect 32641 2021 32647 2073
rect 32699 2021 32705 2073
rect 34273 2021 34279 2073
rect 34331 2021 34337 2073
rect 35905 2021 35911 2073
rect 35963 2021 35969 2073
rect 37537 2021 37543 2073
rect 37595 2021 37601 2073
rect 39169 2021 39175 2073
rect 39227 2021 39233 2073
rect 40801 2021 40807 2073
rect 40859 2021 40865 2073
rect 42433 2021 42439 2073
rect 42491 2021 42497 2073
rect 44065 2021 44071 2073
rect 44123 2021 44129 2073
rect 45697 2021 45703 2073
rect 45755 2021 45761 2073
rect 47329 2021 47335 2073
rect 47387 2021 47393 2073
rect 48961 2021 48967 2073
rect 49019 2021 49025 2073
rect 50593 2021 50599 2073
rect 50651 2021 50657 2073
rect 52225 2021 52231 2073
rect 52283 2021 52289 2073
rect 8 2014 59 2021
rect 1640 2014 1691 2021
rect 3272 2014 3323 2021
rect 4904 2014 4955 2021
rect 6536 2014 6587 2021
rect 8168 2014 8219 2021
rect 9800 2014 9851 2021
rect 11432 2014 11483 2021
rect 13064 2014 13115 2021
rect 14696 2014 14747 2021
rect 16328 2014 16379 2021
rect 17960 2014 18011 2021
rect 19592 2014 19643 2021
rect 21224 2014 21275 2021
rect 22856 2014 22907 2021
rect 24488 2014 24539 2021
rect 26120 2014 26171 2021
rect 27752 2014 27803 2021
rect 29384 2014 29435 2021
rect 31016 2014 31067 2021
rect 32648 2014 32699 2021
rect 34280 2014 34331 2021
rect 35912 2014 35963 2021
rect 37544 2014 37595 2021
rect 39176 2014 39227 2021
rect 40808 2014 40859 2021
rect 42440 2014 42491 2021
rect 44072 2014 44123 2021
rect 45704 2014 45755 2021
rect 47336 2014 47387 2021
rect 48968 2014 49019 2021
rect 50600 2014 50651 2021
rect 52232 2014 52283 2021
rect 8 1869 59 1876
rect 1640 1869 1691 1876
rect 3272 1869 3323 1876
rect 4904 1869 4955 1876
rect 6536 1869 6587 1876
rect 8168 1869 8219 1876
rect 9800 1869 9851 1876
rect 11432 1869 11483 1876
rect 13064 1869 13115 1876
rect 14696 1869 14747 1876
rect 16328 1869 16379 1876
rect 17960 1869 18011 1876
rect 19592 1869 19643 1876
rect 21224 1869 21275 1876
rect 22856 1869 22907 1876
rect 24488 1869 24539 1876
rect 26120 1869 26171 1876
rect 27752 1869 27803 1876
rect 29384 1869 29435 1876
rect 31016 1869 31067 1876
rect 32648 1869 32699 1876
rect 34280 1869 34331 1876
rect 35912 1869 35963 1876
rect 37544 1869 37595 1876
rect 39176 1869 39227 1876
rect 40808 1869 40859 1876
rect 42440 1869 42491 1876
rect 44072 1869 44123 1876
rect 45704 1869 45755 1876
rect 47336 1869 47387 1876
rect 48968 1869 49019 1876
rect 50600 1869 50651 1876
rect 52232 1869 52283 1876
rect 1 1817 7 1869
rect 59 1817 65 1869
rect 1633 1817 1639 1869
rect 1691 1817 1697 1869
rect 3265 1817 3271 1869
rect 3323 1817 3329 1869
rect 4897 1817 4903 1869
rect 4955 1817 4961 1869
rect 6529 1817 6535 1869
rect 6587 1817 6593 1869
rect 8161 1817 8167 1869
rect 8219 1817 8225 1869
rect 9793 1817 9799 1869
rect 9851 1817 9857 1869
rect 11425 1817 11431 1869
rect 11483 1817 11489 1869
rect 13057 1817 13063 1869
rect 13115 1817 13121 1869
rect 14689 1817 14695 1869
rect 14747 1817 14753 1869
rect 16321 1817 16327 1869
rect 16379 1817 16385 1869
rect 17953 1817 17959 1869
rect 18011 1817 18017 1869
rect 19585 1817 19591 1869
rect 19643 1817 19649 1869
rect 21217 1817 21223 1869
rect 21275 1817 21281 1869
rect 22849 1817 22855 1869
rect 22907 1817 22913 1869
rect 24481 1817 24487 1869
rect 24539 1817 24545 1869
rect 26113 1817 26119 1869
rect 26171 1817 26177 1869
rect 27745 1817 27751 1869
rect 27803 1817 27809 1869
rect 29377 1817 29383 1869
rect 29435 1817 29441 1869
rect 31009 1817 31015 1869
rect 31067 1817 31073 1869
rect 32641 1817 32647 1869
rect 32699 1817 32705 1869
rect 34273 1817 34279 1869
rect 34331 1817 34337 1869
rect 35905 1817 35911 1869
rect 35963 1817 35969 1869
rect 37537 1817 37543 1869
rect 37595 1817 37601 1869
rect 39169 1817 39175 1869
rect 39227 1817 39233 1869
rect 40801 1817 40807 1869
rect 40859 1817 40865 1869
rect 42433 1817 42439 1869
rect 42491 1817 42497 1869
rect 44065 1817 44071 1869
rect 44123 1817 44129 1869
rect 45697 1817 45703 1869
rect 45755 1817 45761 1869
rect 47329 1817 47335 1869
rect 47387 1817 47393 1869
rect 48961 1817 48967 1869
rect 49019 1817 49025 1869
rect 50593 1817 50599 1869
rect 50651 1817 50657 1869
rect 52225 1817 52231 1869
rect 52283 1817 52289 1869
rect 8 1810 59 1817
rect 1640 1810 1691 1817
rect 3272 1810 3323 1817
rect 4904 1810 4955 1817
rect 6536 1810 6587 1817
rect 8168 1810 8219 1817
rect 9800 1810 9851 1817
rect 11432 1810 11483 1817
rect 13064 1810 13115 1817
rect 14696 1810 14747 1817
rect 16328 1810 16379 1817
rect 17960 1810 18011 1817
rect 19592 1810 19643 1817
rect 21224 1810 21275 1817
rect 22856 1810 22907 1817
rect 24488 1810 24539 1817
rect 26120 1810 26171 1817
rect 27752 1810 27803 1817
rect 29384 1810 29435 1817
rect 31016 1810 31067 1817
rect 32648 1810 32699 1817
rect 34280 1810 34331 1817
rect 35912 1810 35963 1817
rect 37544 1810 37595 1817
rect 39176 1810 39227 1817
rect 40808 1810 40859 1817
rect 42440 1810 42491 1817
rect 44072 1810 44123 1817
rect 45704 1810 45755 1817
rect 47336 1810 47387 1817
rect 48968 1810 49019 1817
rect 50600 1810 50651 1817
rect 52232 1810 52283 1817
rect 8 1665 59 1672
rect 1640 1665 1691 1672
rect 3272 1665 3323 1672
rect 4904 1665 4955 1672
rect 6536 1665 6587 1672
rect 8168 1665 8219 1672
rect 9800 1665 9851 1672
rect 11432 1665 11483 1672
rect 13064 1665 13115 1672
rect 14696 1665 14747 1672
rect 16328 1665 16379 1672
rect 17960 1665 18011 1672
rect 19592 1665 19643 1672
rect 21224 1665 21275 1672
rect 22856 1665 22907 1672
rect 24488 1665 24539 1672
rect 26120 1665 26171 1672
rect 27752 1665 27803 1672
rect 29384 1665 29435 1672
rect 31016 1665 31067 1672
rect 32648 1665 32699 1672
rect 34280 1665 34331 1672
rect 35912 1665 35963 1672
rect 37544 1665 37595 1672
rect 39176 1665 39227 1672
rect 40808 1665 40859 1672
rect 42440 1665 42491 1672
rect 44072 1665 44123 1672
rect 45704 1665 45755 1672
rect 47336 1665 47387 1672
rect 48968 1665 49019 1672
rect 50600 1665 50651 1672
rect 52232 1665 52283 1672
rect 1 1613 7 1665
rect 59 1613 65 1665
rect 1633 1613 1639 1665
rect 1691 1613 1697 1665
rect 3265 1613 3271 1665
rect 3323 1613 3329 1665
rect 4897 1613 4903 1665
rect 4955 1613 4961 1665
rect 6529 1613 6535 1665
rect 6587 1613 6593 1665
rect 8161 1613 8167 1665
rect 8219 1613 8225 1665
rect 9793 1613 9799 1665
rect 9851 1613 9857 1665
rect 11425 1613 11431 1665
rect 11483 1613 11489 1665
rect 13057 1613 13063 1665
rect 13115 1613 13121 1665
rect 14689 1613 14695 1665
rect 14747 1613 14753 1665
rect 16321 1613 16327 1665
rect 16379 1613 16385 1665
rect 17953 1613 17959 1665
rect 18011 1613 18017 1665
rect 19585 1613 19591 1665
rect 19643 1613 19649 1665
rect 21217 1613 21223 1665
rect 21275 1613 21281 1665
rect 22849 1613 22855 1665
rect 22907 1613 22913 1665
rect 24481 1613 24487 1665
rect 24539 1613 24545 1665
rect 26113 1613 26119 1665
rect 26171 1613 26177 1665
rect 27745 1613 27751 1665
rect 27803 1613 27809 1665
rect 29377 1613 29383 1665
rect 29435 1613 29441 1665
rect 31009 1613 31015 1665
rect 31067 1613 31073 1665
rect 32641 1613 32647 1665
rect 32699 1613 32705 1665
rect 34273 1613 34279 1665
rect 34331 1613 34337 1665
rect 35905 1613 35911 1665
rect 35963 1613 35969 1665
rect 37537 1613 37543 1665
rect 37595 1613 37601 1665
rect 39169 1613 39175 1665
rect 39227 1613 39233 1665
rect 40801 1613 40807 1665
rect 40859 1613 40865 1665
rect 42433 1613 42439 1665
rect 42491 1613 42497 1665
rect 44065 1613 44071 1665
rect 44123 1613 44129 1665
rect 45697 1613 45703 1665
rect 45755 1613 45761 1665
rect 47329 1613 47335 1665
rect 47387 1613 47393 1665
rect 48961 1613 48967 1665
rect 49019 1613 49025 1665
rect 50593 1613 50599 1665
rect 50651 1613 50657 1665
rect 52225 1613 52231 1665
rect 52283 1613 52289 1665
rect 8 1606 59 1613
rect 1640 1606 1691 1613
rect 3272 1606 3323 1613
rect 4904 1606 4955 1613
rect 6536 1606 6587 1613
rect 8168 1606 8219 1613
rect 9800 1606 9851 1613
rect 11432 1606 11483 1613
rect 13064 1606 13115 1613
rect 14696 1606 14747 1613
rect 16328 1606 16379 1613
rect 17960 1606 18011 1613
rect 19592 1606 19643 1613
rect 21224 1606 21275 1613
rect 22856 1606 22907 1613
rect 24488 1606 24539 1613
rect 26120 1606 26171 1613
rect 27752 1606 27803 1613
rect 29384 1606 29435 1613
rect 31016 1606 31067 1613
rect 32648 1606 32699 1613
rect 34280 1606 34331 1613
rect 35912 1606 35963 1613
rect 37544 1606 37595 1613
rect 39176 1606 39227 1613
rect 40808 1606 40859 1613
rect 42440 1606 42491 1613
rect 44072 1606 44123 1613
rect 45704 1606 45755 1613
rect 47336 1606 47387 1613
rect 48968 1606 49019 1613
rect 50600 1606 50651 1613
rect 52232 1606 52283 1613
rect 8 1461 59 1468
rect 1640 1461 1691 1468
rect 3272 1461 3323 1468
rect 4904 1461 4955 1468
rect 6536 1461 6587 1468
rect 8168 1461 8219 1468
rect 9800 1461 9851 1468
rect 11432 1461 11483 1468
rect 13064 1461 13115 1468
rect 14696 1461 14747 1468
rect 16328 1461 16379 1468
rect 17960 1461 18011 1468
rect 19592 1461 19643 1468
rect 21224 1461 21275 1468
rect 22856 1461 22907 1468
rect 24488 1461 24539 1468
rect 26120 1461 26171 1468
rect 27752 1461 27803 1468
rect 29384 1461 29435 1468
rect 31016 1461 31067 1468
rect 32648 1461 32699 1468
rect 34280 1461 34331 1468
rect 35912 1461 35963 1468
rect 37544 1461 37595 1468
rect 39176 1461 39227 1468
rect 40808 1461 40859 1468
rect 42440 1461 42491 1468
rect 44072 1461 44123 1468
rect 45704 1461 45755 1468
rect 47336 1461 47387 1468
rect 48968 1461 49019 1468
rect 50600 1461 50651 1468
rect 52232 1461 52283 1468
rect 1 1409 7 1461
rect 59 1409 65 1461
rect 1633 1409 1639 1461
rect 1691 1409 1697 1461
rect 3265 1409 3271 1461
rect 3323 1409 3329 1461
rect 4897 1409 4903 1461
rect 4955 1409 4961 1461
rect 6529 1409 6535 1461
rect 6587 1409 6593 1461
rect 8161 1409 8167 1461
rect 8219 1409 8225 1461
rect 9793 1409 9799 1461
rect 9851 1409 9857 1461
rect 11425 1409 11431 1461
rect 11483 1409 11489 1461
rect 13057 1409 13063 1461
rect 13115 1409 13121 1461
rect 14689 1409 14695 1461
rect 14747 1409 14753 1461
rect 16321 1409 16327 1461
rect 16379 1409 16385 1461
rect 17953 1409 17959 1461
rect 18011 1409 18017 1461
rect 19585 1409 19591 1461
rect 19643 1409 19649 1461
rect 21217 1409 21223 1461
rect 21275 1409 21281 1461
rect 22849 1409 22855 1461
rect 22907 1409 22913 1461
rect 24481 1409 24487 1461
rect 24539 1409 24545 1461
rect 26113 1409 26119 1461
rect 26171 1409 26177 1461
rect 27745 1409 27751 1461
rect 27803 1409 27809 1461
rect 29377 1409 29383 1461
rect 29435 1409 29441 1461
rect 31009 1409 31015 1461
rect 31067 1409 31073 1461
rect 32641 1409 32647 1461
rect 32699 1409 32705 1461
rect 34273 1409 34279 1461
rect 34331 1409 34337 1461
rect 35905 1409 35911 1461
rect 35963 1409 35969 1461
rect 37537 1409 37543 1461
rect 37595 1409 37601 1461
rect 39169 1409 39175 1461
rect 39227 1409 39233 1461
rect 40801 1409 40807 1461
rect 40859 1409 40865 1461
rect 42433 1409 42439 1461
rect 42491 1409 42497 1461
rect 44065 1409 44071 1461
rect 44123 1409 44129 1461
rect 45697 1409 45703 1461
rect 45755 1409 45761 1461
rect 47329 1409 47335 1461
rect 47387 1409 47393 1461
rect 48961 1409 48967 1461
rect 49019 1409 49025 1461
rect 50593 1409 50599 1461
rect 50651 1409 50657 1461
rect 52225 1409 52231 1461
rect 52283 1409 52289 1461
rect 8 1402 59 1409
rect 1640 1402 1691 1409
rect 3272 1402 3323 1409
rect 4904 1402 4955 1409
rect 6536 1402 6587 1409
rect 8168 1402 8219 1409
rect 9800 1402 9851 1409
rect 11432 1402 11483 1409
rect 13064 1402 13115 1409
rect 14696 1402 14747 1409
rect 16328 1402 16379 1409
rect 17960 1402 18011 1409
rect 19592 1402 19643 1409
rect 21224 1402 21275 1409
rect 22856 1402 22907 1409
rect 24488 1402 24539 1409
rect 26120 1402 26171 1409
rect 27752 1402 27803 1409
rect 29384 1402 29435 1409
rect 31016 1402 31067 1409
rect 32648 1402 32699 1409
rect 34280 1402 34331 1409
rect 35912 1402 35963 1409
rect 37544 1402 37595 1409
rect 39176 1402 39227 1409
rect 40808 1402 40859 1409
rect 42440 1402 42491 1409
rect 44072 1402 44123 1409
rect 45704 1402 45755 1409
rect 47336 1402 47387 1409
rect 48968 1402 49019 1409
rect 50600 1402 50651 1409
rect 52232 1402 52283 1409
rect 8 1257 59 1264
rect 1640 1257 1691 1264
rect 3272 1257 3323 1264
rect 4904 1257 4955 1264
rect 6536 1257 6587 1264
rect 8168 1257 8219 1264
rect 9800 1257 9851 1264
rect 11432 1257 11483 1264
rect 13064 1257 13115 1264
rect 14696 1257 14747 1264
rect 16328 1257 16379 1264
rect 17960 1257 18011 1264
rect 19592 1257 19643 1264
rect 21224 1257 21275 1264
rect 22856 1257 22907 1264
rect 24488 1257 24539 1264
rect 26120 1257 26171 1264
rect 27752 1257 27803 1264
rect 29384 1257 29435 1264
rect 31016 1257 31067 1264
rect 32648 1257 32699 1264
rect 34280 1257 34331 1264
rect 35912 1257 35963 1264
rect 37544 1257 37595 1264
rect 39176 1257 39227 1264
rect 40808 1257 40859 1264
rect 42440 1257 42491 1264
rect 44072 1257 44123 1264
rect 45704 1257 45755 1264
rect 47336 1257 47387 1264
rect 48968 1257 49019 1264
rect 50600 1257 50651 1264
rect 52232 1257 52283 1264
rect 1 1205 7 1257
rect 59 1205 65 1257
rect 1633 1205 1639 1257
rect 1691 1205 1697 1257
rect 3265 1205 3271 1257
rect 3323 1205 3329 1257
rect 4897 1205 4903 1257
rect 4955 1205 4961 1257
rect 6529 1205 6535 1257
rect 6587 1205 6593 1257
rect 8161 1205 8167 1257
rect 8219 1205 8225 1257
rect 9793 1205 9799 1257
rect 9851 1205 9857 1257
rect 11425 1205 11431 1257
rect 11483 1205 11489 1257
rect 13057 1205 13063 1257
rect 13115 1205 13121 1257
rect 14689 1205 14695 1257
rect 14747 1205 14753 1257
rect 16321 1205 16327 1257
rect 16379 1205 16385 1257
rect 17953 1205 17959 1257
rect 18011 1205 18017 1257
rect 19585 1205 19591 1257
rect 19643 1205 19649 1257
rect 21217 1205 21223 1257
rect 21275 1205 21281 1257
rect 22849 1205 22855 1257
rect 22907 1205 22913 1257
rect 24481 1205 24487 1257
rect 24539 1205 24545 1257
rect 26113 1205 26119 1257
rect 26171 1205 26177 1257
rect 27745 1205 27751 1257
rect 27803 1205 27809 1257
rect 29377 1205 29383 1257
rect 29435 1205 29441 1257
rect 31009 1205 31015 1257
rect 31067 1205 31073 1257
rect 32641 1205 32647 1257
rect 32699 1205 32705 1257
rect 34273 1205 34279 1257
rect 34331 1205 34337 1257
rect 35905 1205 35911 1257
rect 35963 1205 35969 1257
rect 37537 1205 37543 1257
rect 37595 1205 37601 1257
rect 39169 1205 39175 1257
rect 39227 1205 39233 1257
rect 40801 1205 40807 1257
rect 40859 1205 40865 1257
rect 42433 1205 42439 1257
rect 42491 1205 42497 1257
rect 44065 1205 44071 1257
rect 44123 1205 44129 1257
rect 45697 1205 45703 1257
rect 45755 1205 45761 1257
rect 47329 1205 47335 1257
rect 47387 1205 47393 1257
rect 48961 1205 48967 1257
rect 49019 1205 49025 1257
rect 50593 1205 50599 1257
rect 50651 1205 50657 1257
rect 52225 1205 52231 1257
rect 52283 1205 52289 1257
rect 8 1198 59 1205
rect 1640 1198 1691 1205
rect 3272 1198 3323 1205
rect 4904 1198 4955 1205
rect 6536 1198 6587 1205
rect 8168 1198 8219 1205
rect 9800 1198 9851 1205
rect 11432 1198 11483 1205
rect 13064 1198 13115 1205
rect 14696 1198 14747 1205
rect 16328 1198 16379 1205
rect 17960 1198 18011 1205
rect 19592 1198 19643 1205
rect 21224 1198 21275 1205
rect 22856 1198 22907 1205
rect 24488 1198 24539 1205
rect 26120 1198 26171 1205
rect 27752 1198 27803 1205
rect 29384 1198 29435 1205
rect 31016 1198 31067 1205
rect 32648 1198 32699 1205
rect 34280 1198 34331 1205
rect 35912 1198 35963 1205
rect 37544 1198 37595 1205
rect 39176 1198 39227 1205
rect 40808 1198 40859 1205
rect 42440 1198 42491 1205
rect 44072 1198 44123 1205
rect 45704 1198 45755 1205
rect 47336 1198 47387 1205
rect 48968 1198 49019 1205
rect 50600 1198 50651 1205
rect 52232 1198 52283 1205
rect 8 1053 59 1060
rect 1640 1053 1691 1060
rect 3272 1053 3323 1060
rect 4904 1053 4955 1060
rect 6536 1053 6587 1060
rect 8168 1053 8219 1060
rect 9800 1053 9851 1060
rect 11432 1053 11483 1060
rect 13064 1053 13115 1060
rect 14696 1053 14747 1060
rect 16328 1053 16379 1060
rect 17960 1053 18011 1060
rect 19592 1053 19643 1060
rect 21224 1053 21275 1060
rect 22856 1053 22907 1060
rect 24488 1053 24539 1060
rect 26120 1053 26171 1060
rect 27752 1053 27803 1060
rect 29384 1053 29435 1060
rect 31016 1053 31067 1060
rect 32648 1053 32699 1060
rect 34280 1053 34331 1060
rect 35912 1053 35963 1060
rect 37544 1053 37595 1060
rect 39176 1053 39227 1060
rect 40808 1053 40859 1060
rect 42440 1053 42491 1060
rect 44072 1053 44123 1060
rect 45704 1053 45755 1060
rect 47336 1053 47387 1060
rect 48968 1053 49019 1060
rect 50600 1053 50651 1060
rect 52232 1053 52283 1060
rect 1 1001 7 1053
rect 59 1001 65 1053
rect 1633 1001 1639 1053
rect 1691 1001 1697 1053
rect 3265 1001 3271 1053
rect 3323 1001 3329 1053
rect 4897 1001 4903 1053
rect 4955 1001 4961 1053
rect 6529 1001 6535 1053
rect 6587 1001 6593 1053
rect 8161 1001 8167 1053
rect 8219 1001 8225 1053
rect 9793 1001 9799 1053
rect 9851 1001 9857 1053
rect 11425 1001 11431 1053
rect 11483 1001 11489 1053
rect 13057 1001 13063 1053
rect 13115 1001 13121 1053
rect 14689 1001 14695 1053
rect 14747 1001 14753 1053
rect 16321 1001 16327 1053
rect 16379 1001 16385 1053
rect 17953 1001 17959 1053
rect 18011 1001 18017 1053
rect 19585 1001 19591 1053
rect 19643 1001 19649 1053
rect 21217 1001 21223 1053
rect 21275 1001 21281 1053
rect 22849 1001 22855 1053
rect 22907 1001 22913 1053
rect 24481 1001 24487 1053
rect 24539 1001 24545 1053
rect 26113 1001 26119 1053
rect 26171 1001 26177 1053
rect 27745 1001 27751 1053
rect 27803 1001 27809 1053
rect 29377 1001 29383 1053
rect 29435 1001 29441 1053
rect 31009 1001 31015 1053
rect 31067 1001 31073 1053
rect 32641 1001 32647 1053
rect 32699 1001 32705 1053
rect 34273 1001 34279 1053
rect 34331 1001 34337 1053
rect 35905 1001 35911 1053
rect 35963 1001 35969 1053
rect 37537 1001 37543 1053
rect 37595 1001 37601 1053
rect 39169 1001 39175 1053
rect 39227 1001 39233 1053
rect 40801 1001 40807 1053
rect 40859 1001 40865 1053
rect 42433 1001 42439 1053
rect 42491 1001 42497 1053
rect 44065 1001 44071 1053
rect 44123 1001 44129 1053
rect 45697 1001 45703 1053
rect 45755 1001 45761 1053
rect 47329 1001 47335 1053
rect 47387 1001 47393 1053
rect 48961 1001 48967 1053
rect 49019 1001 49025 1053
rect 50593 1001 50599 1053
rect 50651 1001 50657 1053
rect 52225 1001 52231 1053
rect 52283 1001 52289 1053
rect 8 994 59 1001
rect 1640 994 1691 1001
rect 3272 994 3323 1001
rect 4904 994 4955 1001
rect 6536 994 6587 1001
rect 8168 994 8219 1001
rect 9800 994 9851 1001
rect 11432 994 11483 1001
rect 13064 994 13115 1001
rect 14696 994 14747 1001
rect 16328 994 16379 1001
rect 17960 994 18011 1001
rect 19592 994 19643 1001
rect 21224 994 21275 1001
rect 22856 994 22907 1001
rect 24488 994 24539 1001
rect 26120 994 26171 1001
rect 27752 994 27803 1001
rect 29384 994 29435 1001
rect 31016 994 31067 1001
rect 32648 994 32699 1001
rect 34280 994 34331 1001
rect 35912 994 35963 1001
rect 37544 994 37595 1001
rect 39176 994 39227 1001
rect 40808 994 40859 1001
rect 42440 994 42491 1001
rect 44072 994 44123 1001
rect 45704 994 45755 1001
rect 47336 994 47387 1001
rect 48968 994 49019 1001
rect 50600 994 50651 1001
rect 52232 994 52283 1001
rect 128 -14 156 977
rect 218 899 270 905
rect 218 841 270 847
rect 332 -14 360 977
rect 422 899 474 905
rect 422 841 474 847
rect 536 -14 564 977
rect 626 899 678 905
rect 626 841 678 847
rect 740 -14 768 977
rect 830 899 882 905
rect 830 841 882 847
rect 944 -14 972 977
rect 1034 899 1086 905
rect 1034 841 1086 847
rect 1148 -14 1176 977
rect 1238 899 1290 905
rect 1238 841 1290 847
rect 1352 -14 1380 977
rect 1442 899 1494 905
rect 1442 841 1494 847
rect 1556 -14 1584 977
rect 1646 899 1698 905
rect 1646 841 1698 847
rect 1760 -14 1788 977
rect 1850 899 1902 905
rect 1850 841 1902 847
rect 1964 -14 1992 977
rect 2054 899 2106 905
rect 2054 841 2106 847
rect 2168 -14 2196 977
rect 2258 899 2310 905
rect 2258 841 2310 847
rect 2372 -14 2400 977
rect 2462 899 2514 905
rect 2462 841 2514 847
rect 2576 -14 2604 977
rect 2666 899 2718 905
rect 2666 841 2718 847
rect 2780 -14 2808 977
rect 2870 899 2922 905
rect 2870 841 2922 847
rect 2984 -14 3012 977
rect 3074 899 3126 905
rect 3074 841 3126 847
rect 3188 -14 3216 977
rect 3278 899 3330 905
rect 3278 841 3330 847
rect 3392 -14 3420 977
rect 3482 899 3534 905
rect 3482 841 3534 847
rect 3596 -14 3624 977
rect 3686 899 3738 905
rect 3686 841 3738 847
rect 3800 -14 3828 977
rect 3890 899 3942 905
rect 3890 841 3942 847
rect 4004 -14 4032 977
rect 4094 899 4146 905
rect 4094 841 4146 847
rect 4208 -14 4236 977
rect 4298 899 4350 905
rect 4298 841 4350 847
rect 4412 -14 4440 977
rect 4502 899 4554 905
rect 4502 841 4554 847
rect 4616 -14 4644 977
rect 4706 899 4758 905
rect 4706 841 4758 847
rect 4820 -14 4848 977
rect 4910 899 4962 905
rect 4910 841 4962 847
rect 5024 -14 5052 977
rect 5114 899 5166 905
rect 5114 841 5166 847
rect 5228 -14 5256 977
rect 5318 899 5370 905
rect 5318 841 5370 847
rect 5432 -14 5460 977
rect 5522 899 5574 905
rect 5522 841 5574 847
rect 5636 -14 5664 977
rect 5726 899 5778 905
rect 5726 841 5778 847
rect 5840 -14 5868 977
rect 5930 899 5982 905
rect 5930 841 5982 847
rect 6044 -14 6072 977
rect 6134 899 6186 905
rect 6134 841 6186 847
rect 6248 -14 6276 977
rect 6338 899 6390 905
rect 6338 841 6390 847
rect 6452 -14 6480 977
rect 6542 899 6594 905
rect 6542 841 6594 847
rect 6656 -14 6684 977
rect 6746 899 6798 905
rect 6746 841 6798 847
rect 6860 -14 6888 977
rect 6950 899 7002 905
rect 6950 841 7002 847
rect 7064 -14 7092 977
rect 7154 899 7206 905
rect 7154 841 7206 847
rect 7268 -14 7296 977
rect 7358 899 7410 905
rect 7358 841 7410 847
rect 7472 -14 7500 977
rect 7562 899 7614 905
rect 7562 841 7614 847
rect 7676 -14 7704 977
rect 7766 899 7818 905
rect 7766 841 7818 847
rect 7880 -14 7908 977
rect 7970 899 8022 905
rect 7970 841 8022 847
rect 8084 -14 8112 977
rect 8174 899 8226 905
rect 8174 841 8226 847
rect 8288 -14 8316 977
rect 8378 899 8430 905
rect 8378 841 8430 847
rect 8492 -14 8520 977
rect 8582 899 8634 905
rect 8582 841 8634 847
rect 8696 -14 8724 977
rect 8786 899 8838 905
rect 8786 841 8838 847
rect 8900 -14 8928 977
rect 8990 899 9042 905
rect 8990 841 9042 847
rect 9104 -14 9132 977
rect 9194 899 9246 905
rect 9194 841 9246 847
rect 9308 -14 9336 977
rect 9398 899 9450 905
rect 9398 841 9450 847
rect 9512 -14 9540 977
rect 9602 899 9654 905
rect 9602 841 9654 847
rect 9716 -14 9744 977
rect 9806 899 9858 905
rect 9806 841 9858 847
rect 9920 -14 9948 977
rect 10010 899 10062 905
rect 10010 841 10062 847
rect 10124 -14 10152 977
rect 10214 899 10266 905
rect 10214 841 10266 847
rect 10328 -14 10356 977
rect 10418 899 10470 905
rect 10418 841 10470 847
rect 10532 -14 10560 977
rect 10622 899 10674 905
rect 10622 841 10674 847
rect 10736 -14 10764 977
rect 10826 899 10878 905
rect 10826 841 10878 847
rect 10940 -14 10968 977
rect 11030 899 11082 905
rect 11030 841 11082 847
rect 11144 -14 11172 977
rect 11234 899 11286 905
rect 11234 841 11286 847
rect 11348 -14 11376 977
rect 11438 899 11490 905
rect 11438 841 11490 847
rect 11552 -14 11580 977
rect 11642 899 11694 905
rect 11642 841 11694 847
rect 11756 -14 11784 977
rect 11846 899 11898 905
rect 11846 841 11898 847
rect 11960 -14 11988 977
rect 12050 899 12102 905
rect 12050 841 12102 847
rect 12164 -14 12192 977
rect 12254 899 12306 905
rect 12254 841 12306 847
rect 12368 -14 12396 977
rect 12458 899 12510 905
rect 12458 841 12510 847
rect 12572 -14 12600 977
rect 12662 899 12714 905
rect 12662 841 12714 847
rect 12776 -14 12804 977
rect 12866 899 12918 905
rect 12866 841 12918 847
rect 12980 -14 13008 977
rect 13070 899 13122 905
rect 13070 841 13122 847
rect 13184 -14 13212 977
rect 13274 899 13326 905
rect 13274 841 13326 847
rect 13388 -14 13416 977
rect 13478 899 13530 905
rect 13478 841 13530 847
rect 13592 -14 13620 977
rect 13682 899 13734 905
rect 13682 841 13734 847
rect 13796 -14 13824 977
rect 13886 899 13938 905
rect 13886 841 13938 847
rect 14000 -14 14028 977
rect 14090 899 14142 905
rect 14090 841 14142 847
rect 14204 -14 14232 977
rect 14294 899 14346 905
rect 14294 841 14346 847
rect 14408 -14 14436 977
rect 14498 899 14550 905
rect 14498 841 14550 847
rect 14612 -14 14640 977
rect 14702 899 14754 905
rect 14702 841 14754 847
rect 14816 -14 14844 977
rect 14906 899 14958 905
rect 14906 841 14958 847
rect 15020 -14 15048 977
rect 15110 899 15162 905
rect 15110 841 15162 847
rect 15224 -14 15252 977
rect 15314 899 15366 905
rect 15314 841 15366 847
rect 15428 -14 15456 977
rect 15518 899 15570 905
rect 15518 841 15570 847
rect 15632 -14 15660 977
rect 15722 899 15774 905
rect 15722 841 15774 847
rect 15836 -14 15864 977
rect 15926 899 15978 905
rect 15926 841 15978 847
rect 16040 -14 16068 977
rect 16130 899 16182 905
rect 16130 841 16182 847
rect 16244 -14 16272 977
rect 16334 899 16386 905
rect 16334 841 16386 847
rect 16448 -14 16476 977
rect 16538 899 16590 905
rect 16538 841 16590 847
rect 16652 -14 16680 977
rect 16742 899 16794 905
rect 16742 841 16794 847
rect 16856 -14 16884 977
rect 16946 899 16998 905
rect 16946 841 16998 847
rect 17060 -14 17088 977
rect 17150 899 17202 905
rect 17150 841 17202 847
rect 17264 -14 17292 977
rect 17354 899 17406 905
rect 17354 841 17406 847
rect 17468 -14 17496 977
rect 17558 899 17610 905
rect 17558 841 17610 847
rect 17672 -14 17700 977
rect 17762 899 17814 905
rect 17762 841 17814 847
rect 17876 -14 17904 977
rect 17966 899 18018 905
rect 17966 841 18018 847
rect 18080 -14 18108 977
rect 18170 899 18222 905
rect 18170 841 18222 847
rect 18284 -14 18312 977
rect 18374 899 18426 905
rect 18374 841 18426 847
rect 18488 -14 18516 977
rect 18578 899 18630 905
rect 18578 841 18630 847
rect 18692 -14 18720 977
rect 18782 899 18834 905
rect 18782 841 18834 847
rect 18896 -14 18924 977
rect 18986 899 19038 905
rect 18986 841 19038 847
rect 19100 -14 19128 977
rect 19190 899 19242 905
rect 19190 841 19242 847
rect 19304 -14 19332 977
rect 19394 899 19446 905
rect 19394 841 19446 847
rect 19508 -14 19536 977
rect 19598 899 19650 905
rect 19598 841 19650 847
rect 19712 -14 19740 977
rect 19802 899 19854 905
rect 19802 841 19854 847
rect 19916 -14 19944 977
rect 20006 899 20058 905
rect 20006 841 20058 847
rect 20120 -14 20148 977
rect 20210 899 20262 905
rect 20210 841 20262 847
rect 20324 -14 20352 977
rect 20414 899 20466 905
rect 20414 841 20466 847
rect 20528 -14 20556 977
rect 20618 899 20670 905
rect 20618 841 20670 847
rect 20732 -14 20760 977
rect 20822 899 20874 905
rect 20822 841 20874 847
rect 20936 -14 20964 977
rect 21026 899 21078 905
rect 21026 841 21078 847
rect 21140 -14 21168 977
rect 21230 899 21282 905
rect 21230 841 21282 847
rect 21344 -14 21372 977
rect 21434 899 21486 905
rect 21434 841 21486 847
rect 21548 -14 21576 977
rect 21638 899 21690 905
rect 21638 841 21690 847
rect 21752 -14 21780 977
rect 21842 899 21894 905
rect 21842 841 21894 847
rect 21956 -14 21984 977
rect 22046 899 22098 905
rect 22046 841 22098 847
rect 22160 -14 22188 977
rect 22250 899 22302 905
rect 22250 841 22302 847
rect 22364 -14 22392 977
rect 22454 899 22506 905
rect 22454 841 22506 847
rect 22568 -14 22596 977
rect 22658 899 22710 905
rect 22658 841 22710 847
rect 22772 -14 22800 977
rect 22862 899 22914 905
rect 22862 841 22914 847
rect 22976 -14 23004 977
rect 23066 899 23118 905
rect 23066 841 23118 847
rect 23180 -14 23208 977
rect 23270 899 23322 905
rect 23270 841 23322 847
rect 23384 -14 23412 977
rect 23474 899 23526 905
rect 23474 841 23526 847
rect 23588 -14 23616 977
rect 23678 899 23730 905
rect 23678 841 23730 847
rect 23792 -14 23820 977
rect 23882 899 23934 905
rect 23882 841 23934 847
rect 23996 -14 24024 977
rect 24086 899 24138 905
rect 24086 841 24138 847
rect 24200 -14 24228 977
rect 24290 899 24342 905
rect 24290 841 24342 847
rect 24404 -14 24432 977
rect 24494 899 24546 905
rect 24494 841 24546 847
rect 24608 -14 24636 977
rect 24698 899 24750 905
rect 24698 841 24750 847
rect 24812 -14 24840 977
rect 24902 899 24954 905
rect 24902 841 24954 847
rect 25016 -14 25044 977
rect 25106 899 25158 905
rect 25106 841 25158 847
rect 25220 -14 25248 977
rect 25310 899 25362 905
rect 25310 841 25362 847
rect 25424 -14 25452 977
rect 25514 899 25566 905
rect 25514 841 25566 847
rect 25628 -14 25656 977
rect 25718 899 25770 905
rect 25718 841 25770 847
rect 25832 -14 25860 977
rect 25922 899 25974 905
rect 25922 841 25974 847
rect 26036 -14 26064 977
rect 26126 899 26178 905
rect 26126 841 26178 847
rect 26240 -14 26268 977
rect 26330 899 26382 905
rect 26330 841 26382 847
rect 26444 -14 26472 977
rect 26534 899 26586 905
rect 26534 841 26586 847
rect 26648 -14 26676 977
rect 26738 899 26790 905
rect 26738 841 26790 847
rect 26852 -14 26880 977
rect 26942 899 26994 905
rect 26942 841 26994 847
rect 27056 -14 27084 977
rect 27146 899 27198 905
rect 27146 841 27198 847
rect 27260 -14 27288 977
rect 27350 899 27402 905
rect 27350 841 27402 847
rect 27464 -14 27492 977
rect 27554 899 27606 905
rect 27554 841 27606 847
rect 27668 -14 27696 977
rect 27758 899 27810 905
rect 27758 841 27810 847
rect 27872 -14 27900 977
rect 27962 899 28014 905
rect 27962 841 28014 847
rect 28076 -14 28104 977
rect 28166 899 28218 905
rect 28166 841 28218 847
rect 28280 -14 28308 977
rect 28370 899 28422 905
rect 28370 841 28422 847
rect 28484 -14 28512 977
rect 28574 899 28626 905
rect 28574 841 28626 847
rect 28688 -14 28716 977
rect 28778 899 28830 905
rect 28778 841 28830 847
rect 28892 -14 28920 977
rect 28982 899 29034 905
rect 28982 841 29034 847
rect 29096 -14 29124 977
rect 29186 899 29238 905
rect 29186 841 29238 847
rect 29300 -14 29328 977
rect 29390 899 29442 905
rect 29390 841 29442 847
rect 29504 -14 29532 977
rect 29594 899 29646 905
rect 29594 841 29646 847
rect 29708 -14 29736 977
rect 29798 899 29850 905
rect 29798 841 29850 847
rect 29912 -14 29940 977
rect 30002 899 30054 905
rect 30002 841 30054 847
rect 30116 -14 30144 977
rect 30206 899 30258 905
rect 30206 841 30258 847
rect 30320 -14 30348 977
rect 30410 899 30462 905
rect 30410 841 30462 847
rect 30524 -14 30552 977
rect 30614 899 30666 905
rect 30614 841 30666 847
rect 30728 -14 30756 977
rect 30818 899 30870 905
rect 30818 841 30870 847
rect 30932 -14 30960 977
rect 31022 899 31074 905
rect 31022 841 31074 847
rect 31136 -14 31164 977
rect 31226 899 31278 905
rect 31226 841 31278 847
rect 31340 -14 31368 977
rect 31430 899 31482 905
rect 31430 841 31482 847
rect 31544 -14 31572 977
rect 31634 899 31686 905
rect 31634 841 31686 847
rect 31748 -14 31776 977
rect 31838 899 31890 905
rect 31838 841 31890 847
rect 31952 -14 31980 977
rect 32042 899 32094 905
rect 32042 841 32094 847
rect 32156 -14 32184 977
rect 32246 899 32298 905
rect 32246 841 32298 847
rect 32360 -14 32388 977
rect 32450 899 32502 905
rect 32450 841 32502 847
rect 32564 -14 32592 977
rect 32654 899 32706 905
rect 32654 841 32706 847
rect 32768 -14 32796 977
rect 32858 899 32910 905
rect 32858 841 32910 847
rect 32972 -14 33000 977
rect 33062 899 33114 905
rect 33062 841 33114 847
rect 33176 -14 33204 977
rect 33266 899 33318 905
rect 33266 841 33318 847
rect 33380 -14 33408 977
rect 33470 899 33522 905
rect 33470 841 33522 847
rect 33584 -14 33612 977
rect 33674 899 33726 905
rect 33674 841 33726 847
rect 33788 -14 33816 977
rect 33878 899 33930 905
rect 33878 841 33930 847
rect 33992 -14 34020 977
rect 34082 899 34134 905
rect 34082 841 34134 847
rect 34196 -14 34224 977
rect 34286 899 34338 905
rect 34286 841 34338 847
rect 34400 -14 34428 977
rect 34490 899 34542 905
rect 34490 841 34542 847
rect 34604 -14 34632 977
rect 34694 899 34746 905
rect 34694 841 34746 847
rect 34808 -14 34836 977
rect 34898 899 34950 905
rect 34898 841 34950 847
rect 35012 -14 35040 977
rect 35102 899 35154 905
rect 35102 841 35154 847
rect 35216 -14 35244 977
rect 35306 899 35358 905
rect 35306 841 35358 847
rect 35420 -14 35448 977
rect 35510 899 35562 905
rect 35510 841 35562 847
rect 35624 -14 35652 977
rect 35714 899 35766 905
rect 35714 841 35766 847
rect 35828 -14 35856 977
rect 35918 899 35970 905
rect 35918 841 35970 847
rect 36032 -14 36060 977
rect 36122 899 36174 905
rect 36122 841 36174 847
rect 36236 -14 36264 977
rect 36326 899 36378 905
rect 36326 841 36378 847
rect 36440 -14 36468 977
rect 36530 899 36582 905
rect 36530 841 36582 847
rect 36644 -14 36672 977
rect 36734 899 36786 905
rect 36734 841 36786 847
rect 36848 -14 36876 977
rect 36938 899 36990 905
rect 36938 841 36990 847
rect 37052 -14 37080 977
rect 37142 899 37194 905
rect 37142 841 37194 847
rect 37256 -14 37284 977
rect 37346 899 37398 905
rect 37346 841 37398 847
rect 37460 -14 37488 977
rect 37550 899 37602 905
rect 37550 841 37602 847
rect 37664 -14 37692 977
rect 37754 899 37806 905
rect 37754 841 37806 847
rect 37868 -14 37896 977
rect 37958 899 38010 905
rect 37958 841 38010 847
rect 38072 -14 38100 977
rect 38162 899 38214 905
rect 38162 841 38214 847
rect 38276 -14 38304 977
rect 38366 899 38418 905
rect 38366 841 38418 847
rect 38480 -14 38508 977
rect 38570 899 38622 905
rect 38570 841 38622 847
rect 38684 -14 38712 977
rect 38774 899 38826 905
rect 38774 841 38826 847
rect 38888 -14 38916 977
rect 38978 899 39030 905
rect 38978 841 39030 847
rect 39092 -14 39120 977
rect 39182 899 39234 905
rect 39182 841 39234 847
rect 39296 -14 39324 977
rect 39386 899 39438 905
rect 39386 841 39438 847
rect 39500 -14 39528 977
rect 39590 899 39642 905
rect 39590 841 39642 847
rect 39704 -14 39732 977
rect 39794 899 39846 905
rect 39794 841 39846 847
rect 39908 -14 39936 977
rect 39998 899 40050 905
rect 39998 841 40050 847
rect 40112 -14 40140 977
rect 40202 899 40254 905
rect 40202 841 40254 847
rect 40316 -14 40344 977
rect 40406 899 40458 905
rect 40406 841 40458 847
rect 40520 -14 40548 977
rect 40610 899 40662 905
rect 40610 841 40662 847
rect 40724 -14 40752 977
rect 40814 899 40866 905
rect 40814 841 40866 847
rect 40928 -14 40956 977
rect 41018 899 41070 905
rect 41018 841 41070 847
rect 41132 -14 41160 977
rect 41222 899 41274 905
rect 41222 841 41274 847
rect 41336 -14 41364 977
rect 41426 899 41478 905
rect 41426 841 41478 847
rect 41540 -14 41568 977
rect 41630 899 41682 905
rect 41630 841 41682 847
rect 41744 -14 41772 977
rect 41834 899 41886 905
rect 41834 841 41886 847
rect 41948 -14 41976 977
rect 42038 899 42090 905
rect 42038 841 42090 847
rect 42152 -14 42180 977
rect 42242 899 42294 905
rect 42242 841 42294 847
rect 42356 -14 42384 977
rect 42446 899 42498 905
rect 42446 841 42498 847
rect 42560 -14 42588 977
rect 42650 899 42702 905
rect 42650 841 42702 847
rect 42764 -14 42792 977
rect 42854 899 42906 905
rect 42854 841 42906 847
rect 42968 -14 42996 977
rect 43058 899 43110 905
rect 43058 841 43110 847
rect 43172 -14 43200 977
rect 43262 899 43314 905
rect 43262 841 43314 847
rect 43376 -14 43404 977
rect 43466 899 43518 905
rect 43466 841 43518 847
rect 43580 -14 43608 977
rect 43670 899 43722 905
rect 43670 841 43722 847
rect 43784 -14 43812 977
rect 43874 899 43926 905
rect 43874 841 43926 847
rect 43988 -14 44016 977
rect 44078 899 44130 905
rect 44078 841 44130 847
rect 44192 -14 44220 977
rect 44282 899 44334 905
rect 44282 841 44334 847
rect 44396 -14 44424 977
rect 44486 899 44538 905
rect 44486 841 44538 847
rect 44600 -14 44628 977
rect 44690 899 44742 905
rect 44690 841 44742 847
rect 44804 -14 44832 977
rect 44894 899 44946 905
rect 44894 841 44946 847
rect 45008 -14 45036 977
rect 45098 899 45150 905
rect 45098 841 45150 847
rect 45212 -14 45240 977
rect 45302 899 45354 905
rect 45302 841 45354 847
rect 45416 -14 45444 977
rect 45506 899 45558 905
rect 45506 841 45558 847
rect 45620 -14 45648 977
rect 45710 899 45762 905
rect 45710 841 45762 847
rect 45824 -14 45852 977
rect 45914 899 45966 905
rect 45914 841 45966 847
rect 46028 -14 46056 977
rect 46118 899 46170 905
rect 46118 841 46170 847
rect 46232 -14 46260 977
rect 46322 899 46374 905
rect 46322 841 46374 847
rect 46436 -14 46464 977
rect 46526 899 46578 905
rect 46526 841 46578 847
rect 46640 -14 46668 977
rect 46730 899 46782 905
rect 46730 841 46782 847
rect 46844 -14 46872 977
rect 46934 899 46986 905
rect 46934 841 46986 847
rect 47048 -14 47076 977
rect 47138 899 47190 905
rect 47138 841 47190 847
rect 47252 -14 47280 977
rect 47342 899 47394 905
rect 47342 841 47394 847
rect 47456 -14 47484 977
rect 47546 899 47598 905
rect 47546 841 47598 847
rect 47660 -14 47688 977
rect 47750 899 47802 905
rect 47750 841 47802 847
rect 47864 -14 47892 977
rect 47954 899 48006 905
rect 47954 841 48006 847
rect 48068 -14 48096 977
rect 48158 899 48210 905
rect 48158 841 48210 847
rect 48272 -14 48300 977
rect 48362 899 48414 905
rect 48362 841 48414 847
rect 48476 -14 48504 977
rect 48566 899 48618 905
rect 48566 841 48618 847
rect 48680 -14 48708 977
rect 48770 899 48822 905
rect 48770 841 48822 847
rect 48884 -14 48912 977
rect 48974 899 49026 905
rect 48974 841 49026 847
rect 49088 -14 49116 977
rect 49178 899 49230 905
rect 49178 841 49230 847
rect 49292 -14 49320 977
rect 49382 899 49434 905
rect 49382 841 49434 847
rect 49496 -14 49524 977
rect 49586 899 49638 905
rect 49586 841 49638 847
rect 49700 -14 49728 977
rect 49790 899 49842 905
rect 49790 841 49842 847
rect 49904 -14 49932 977
rect 49994 899 50046 905
rect 49994 841 50046 847
rect 50108 -14 50136 977
rect 50198 899 50250 905
rect 50198 841 50250 847
rect 50312 -14 50340 977
rect 50402 899 50454 905
rect 50402 841 50454 847
rect 50516 -14 50544 977
rect 50606 899 50658 905
rect 50606 841 50658 847
rect 50720 -14 50748 977
rect 50810 899 50862 905
rect 50810 841 50862 847
rect 50924 -14 50952 977
rect 51014 899 51066 905
rect 51014 841 51066 847
rect 51128 -14 51156 977
rect 51218 899 51270 905
rect 51218 841 51270 847
rect 51332 -14 51360 977
rect 51422 899 51474 905
rect 51422 841 51474 847
rect 51536 -14 51564 977
rect 51626 899 51678 905
rect 51626 841 51678 847
rect 51740 -14 51768 977
rect 51830 899 51882 905
rect 51830 841 51882 847
rect 51944 -14 51972 977
rect 52034 899 52086 905
rect 52034 841 52086 847
rect 52148 -14 52176 977
rect 52252 899 52304 905
rect 52252 841 52304 847
rect 52445 396 52473 2645
rect 52299 368 52473 396
<< via1 >>
rect 7 2676 59 2685
rect 7 2642 16 2676
rect 16 2642 50 2676
rect 50 2642 59 2676
rect 7 2633 59 2642
rect 1639 2676 1691 2685
rect 1639 2642 1648 2676
rect 1648 2642 1682 2676
rect 1682 2642 1691 2676
rect 1639 2633 1691 2642
rect 3271 2676 3323 2685
rect 3271 2642 3280 2676
rect 3280 2642 3314 2676
rect 3314 2642 3323 2676
rect 3271 2633 3323 2642
rect 4903 2676 4955 2685
rect 4903 2642 4912 2676
rect 4912 2642 4946 2676
rect 4946 2642 4955 2676
rect 4903 2633 4955 2642
rect 6535 2676 6587 2685
rect 6535 2642 6544 2676
rect 6544 2642 6578 2676
rect 6578 2642 6587 2676
rect 6535 2633 6587 2642
rect 8167 2676 8219 2685
rect 8167 2642 8176 2676
rect 8176 2642 8210 2676
rect 8210 2642 8219 2676
rect 8167 2633 8219 2642
rect 9799 2676 9851 2685
rect 9799 2642 9808 2676
rect 9808 2642 9842 2676
rect 9842 2642 9851 2676
rect 9799 2633 9851 2642
rect 11431 2676 11483 2685
rect 11431 2642 11440 2676
rect 11440 2642 11474 2676
rect 11474 2642 11483 2676
rect 11431 2633 11483 2642
rect 13063 2676 13115 2685
rect 13063 2642 13072 2676
rect 13072 2642 13106 2676
rect 13106 2642 13115 2676
rect 13063 2633 13115 2642
rect 14695 2676 14747 2685
rect 14695 2642 14704 2676
rect 14704 2642 14738 2676
rect 14738 2642 14747 2676
rect 14695 2633 14747 2642
rect 16327 2676 16379 2685
rect 16327 2642 16336 2676
rect 16336 2642 16370 2676
rect 16370 2642 16379 2676
rect 16327 2633 16379 2642
rect 17959 2676 18011 2685
rect 17959 2642 17968 2676
rect 17968 2642 18002 2676
rect 18002 2642 18011 2676
rect 17959 2633 18011 2642
rect 19591 2676 19643 2685
rect 19591 2642 19600 2676
rect 19600 2642 19634 2676
rect 19634 2642 19643 2676
rect 19591 2633 19643 2642
rect 21223 2676 21275 2685
rect 21223 2642 21232 2676
rect 21232 2642 21266 2676
rect 21266 2642 21275 2676
rect 21223 2633 21275 2642
rect 22855 2676 22907 2685
rect 22855 2642 22864 2676
rect 22864 2642 22898 2676
rect 22898 2642 22907 2676
rect 22855 2633 22907 2642
rect 24487 2676 24539 2685
rect 24487 2642 24496 2676
rect 24496 2642 24530 2676
rect 24530 2642 24539 2676
rect 24487 2633 24539 2642
rect 26119 2676 26171 2685
rect 26119 2642 26128 2676
rect 26128 2642 26162 2676
rect 26162 2642 26171 2676
rect 26119 2633 26171 2642
rect 27751 2676 27803 2685
rect 27751 2642 27760 2676
rect 27760 2642 27794 2676
rect 27794 2642 27803 2676
rect 27751 2633 27803 2642
rect 29383 2676 29435 2685
rect 29383 2642 29392 2676
rect 29392 2642 29426 2676
rect 29426 2642 29435 2676
rect 29383 2633 29435 2642
rect 31015 2676 31067 2685
rect 31015 2642 31024 2676
rect 31024 2642 31058 2676
rect 31058 2642 31067 2676
rect 31015 2633 31067 2642
rect 32647 2676 32699 2685
rect 32647 2642 32656 2676
rect 32656 2642 32690 2676
rect 32690 2642 32699 2676
rect 32647 2633 32699 2642
rect 34279 2676 34331 2685
rect 34279 2642 34288 2676
rect 34288 2642 34322 2676
rect 34322 2642 34331 2676
rect 34279 2633 34331 2642
rect 35911 2676 35963 2685
rect 35911 2642 35920 2676
rect 35920 2642 35954 2676
rect 35954 2642 35963 2676
rect 35911 2633 35963 2642
rect 37543 2676 37595 2685
rect 37543 2642 37552 2676
rect 37552 2642 37586 2676
rect 37586 2642 37595 2676
rect 37543 2633 37595 2642
rect 39175 2676 39227 2685
rect 39175 2642 39184 2676
rect 39184 2642 39218 2676
rect 39218 2642 39227 2676
rect 39175 2633 39227 2642
rect 40807 2676 40859 2685
rect 40807 2642 40816 2676
rect 40816 2642 40850 2676
rect 40850 2642 40859 2676
rect 40807 2633 40859 2642
rect 42439 2676 42491 2685
rect 42439 2642 42448 2676
rect 42448 2642 42482 2676
rect 42482 2642 42491 2676
rect 42439 2633 42491 2642
rect 44071 2676 44123 2685
rect 44071 2642 44080 2676
rect 44080 2642 44114 2676
rect 44114 2642 44123 2676
rect 44071 2633 44123 2642
rect 45703 2676 45755 2685
rect 45703 2642 45712 2676
rect 45712 2642 45746 2676
rect 45746 2642 45755 2676
rect 45703 2633 45755 2642
rect 47335 2676 47387 2685
rect 47335 2642 47344 2676
rect 47344 2642 47378 2676
rect 47378 2642 47387 2676
rect 47335 2633 47387 2642
rect 48967 2676 49019 2685
rect 48967 2642 48976 2676
rect 48976 2642 49010 2676
rect 49010 2642 49019 2676
rect 48967 2633 49019 2642
rect 50599 2676 50651 2685
rect 50599 2642 50608 2676
rect 50608 2642 50642 2676
rect 50642 2642 50651 2676
rect 50599 2633 50651 2642
rect 52231 2676 52283 2685
rect 52231 2642 52240 2676
rect 52240 2642 52274 2676
rect 52274 2642 52283 2676
rect 52231 2633 52283 2642
rect 7 2472 59 2481
rect 7 2438 16 2472
rect 16 2438 50 2472
rect 50 2438 59 2472
rect 7 2429 59 2438
rect 1639 2472 1691 2481
rect 1639 2438 1648 2472
rect 1648 2438 1682 2472
rect 1682 2438 1691 2472
rect 1639 2429 1691 2438
rect 3271 2472 3323 2481
rect 3271 2438 3280 2472
rect 3280 2438 3314 2472
rect 3314 2438 3323 2472
rect 3271 2429 3323 2438
rect 4903 2472 4955 2481
rect 4903 2438 4912 2472
rect 4912 2438 4946 2472
rect 4946 2438 4955 2472
rect 4903 2429 4955 2438
rect 6535 2472 6587 2481
rect 6535 2438 6544 2472
rect 6544 2438 6578 2472
rect 6578 2438 6587 2472
rect 6535 2429 6587 2438
rect 8167 2472 8219 2481
rect 8167 2438 8176 2472
rect 8176 2438 8210 2472
rect 8210 2438 8219 2472
rect 8167 2429 8219 2438
rect 9799 2472 9851 2481
rect 9799 2438 9808 2472
rect 9808 2438 9842 2472
rect 9842 2438 9851 2472
rect 9799 2429 9851 2438
rect 11431 2472 11483 2481
rect 11431 2438 11440 2472
rect 11440 2438 11474 2472
rect 11474 2438 11483 2472
rect 11431 2429 11483 2438
rect 13063 2472 13115 2481
rect 13063 2438 13072 2472
rect 13072 2438 13106 2472
rect 13106 2438 13115 2472
rect 13063 2429 13115 2438
rect 14695 2472 14747 2481
rect 14695 2438 14704 2472
rect 14704 2438 14738 2472
rect 14738 2438 14747 2472
rect 14695 2429 14747 2438
rect 16327 2472 16379 2481
rect 16327 2438 16336 2472
rect 16336 2438 16370 2472
rect 16370 2438 16379 2472
rect 16327 2429 16379 2438
rect 17959 2472 18011 2481
rect 17959 2438 17968 2472
rect 17968 2438 18002 2472
rect 18002 2438 18011 2472
rect 17959 2429 18011 2438
rect 19591 2472 19643 2481
rect 19591 2438 19600 2472
rect 19600 2438 19634 2472
rect 19634 2438 19643 2472
rect 19591 2429 19643 2438
rect 21223 2472 21275 2481
rect 21223 2438 21232 2472
rect 21232 2438 21266 2472
rect 21266 2438 21275 2472
rect 21223 2429 21275 2438
rect 22855 2472 22907 2481
rect 22855 2438 22864 2472
rect 22864 2438 22898 2472
rect 22898 2438 22907 2472
rect 22855 2429 22907 2438
rect 24487 2472 24539 2481
rect 24487 2438 24496 2472
rect 24496 2438 24530 2472
rect 24530 2438 24539 2472
rect 24487 2429 24539 2438
rect 26119 2472 26171 2481
rect 26119 2438 26128 2472
rect 26128 2438 26162 2472
rect 26162 2438 26171 2472
rect 26119 2429 26171 2438
rect 27751 2472 27803 2481
rect 27751 2438 27760 2472
rect 27760 2438 27794 2472
rect 27794 2438 27803 2472
rect 27751 2429 27803 2438
rect 29383 2472 29435 2481
rect 29383 2438 29392 2472
rect 29392 2438 29426 2472
rect 29426 2438 29435 2472
rect 29383 2429 29435 2438
rect 31015 2472 31067 2481
rect 31015 2438 31024 2472
rect 31024 2438 31058 2472
rect 31058 2438 31067 2472
rect 31015 2429 31067 2438
rect 32647 2472 32699 2481
rect 32647 2438 32656 2472
rect 32656 2438 32690 2472
rect 32690 2438 32699 2472
rect 32647 2429 32699 2438
rect 34279 2472 34331 2481
rect 34279 2438 34288 2472
rect 34288 2438 34322 2472
rect 34322 2438 34331 2472
rect 34279 2429 34331 2438
rect 35911 2472 35963 2481
rect 35911 2438 35920 2472
rect 35920 2438 35954 2472
rect 35954 2438 35963 2472
rect 35911 2429 35963 2438
rect 37543 2472 37595 2481
rect 37543 2438 37552 2472
rect 37552 2438 37586 2472
rect 37586 2438 37595 2472
rect 37543 2429 37595 2438
rect 39175 2472 39227 2481
rect 39175 2438 39184 2472
rect 39184 2438 39218 2472
rect 39218 2438 39227 2472
rect 39175 2429 39227 2438
rect 40807 2472 40859 2481
rect 40807 2438 40816 2472
rect 40816 2438 40850 2472
rect 40850 2438 40859 2472
rect 40807 2429 40859 2438
rect 42439 2472 42491 2481
rect 42439 2438 42448 2472
rect 42448 2438 42482 2472
rect 42482 2438 42491 2472
rect 42439 2429 42491 2438
rect 44071 2472 44123 2481
rect 44071 2438 44080 2472
rect 44080 2438 44114 2472
rect 44114 2438 44123 2472
rect 44071 2429 44123 2438
rect 45703 2472 45755 2481
rect 45703 2438 45712 2472
rect 45712 2438 45746 2472
rect 45746 2438 45755 2472
rect 45703 2429 45755 2438
rect 47335 2472 47387 2481
rect 47335 2438 47344 2472
rect 47344 2438 47378 2472
rect 47378 2438 47387 2472
rect 47335 2429 47387 2438
rect 48967 2472 49019 2481
rect 48967 2438 48976 2472
rect 48976 2438 49010 2472
rect 49010 2438 49019 2472
rect 48967 2429 49019 2438
rect 50599 2472 50651 2481
rect 50599 2438 50608 2472
rect 50608 2438 50642 2472
rect 50642 2438 50651 2472
rect 50599 2429 50651 2438
rect 52231 2472 52283 2481
rect 52231 2438 52240 2472
rect 52240 2438 52274 2472
rect 52274 2438 52283 2472
rect 52231 2429 52283 2438
rect 7 2268 59 2277
rect 7 2234 16 2268
rect 16 2234 50 2268
rect 50 2234 59 2268
rect 7 2225 59 2234
rect 1639 2268 1691 2277
rect 1639 2234 1648 2268
rect 1648 2234 1682 2268
rect 1682 2234 1691 2268
rect 1639 2225 1691 2234
rect 3271 2268 3323 2277
rect 3271 2234 3280 2268
rect 3280 2234 3314 2268
rect 3314 2234 3323 2268
rect 3271 2225 3323 2234
rect 4903 2268 4955 2277
rect 4903 2234 4912 2268
rect 4912 2234 4946 2268
rect 4946 2234 4955 2268
rect 4903 2225 4955 2234
rect 6535 2268 6587 2277
rect 6535 2234 6544 2268
rect 6544 2234 6578 2268
rect 6578 2234 6587 2268
rect 6535 2225 6587 2234
rect 8167 2268 8219 2277
rect 8167 2234 8176 2268
rect 8176 2234 8210 2268
rect 8210 2234 8219 2268
rect 8167 2225 8219 2234
rect 9799 2268 9851 2277
rect 9799 2234 9808 2268
rect 9808 2234 9842 2268
rect 9842 2234 9851 2268
rect 9799 2225 9851 2234
rect 11431 2268 11483 2277
rect 11431 2234 11440 2268
rect 11440 2234 11474 2268
rect 11474 2234 11483 2268
rect 11431 2225 11483 2234
rect 13063 2268 13115 2277
rect 13063 2234 13072 2268
rect 13072 2234 13106 2268
rect 13106 2234 13115 2268
rect 13063 2225 13115 2234
rect 14695 2268 14747 2277
rect 14695 2234 14704 2268
rect 14704 2234 14738 2268
rect 14738 2234 14747 2268
rect 14695 2225 14747 2234
rect 16327 2268 16379 2277
rect 16327 2234 16336 2268
rect 16336 2234 16370 2268
rect 16370 2234 16379 2268
rect 16327 2225 16379 2234
rect 17959 2268 18011 2277
rect 17959 2234 17968 2268
rect 17968 2234 18002 2268
rect 18002 2234 18011 2268
rect 17959 2225 18011 2234
rect 19591 2268 19643 2277
rect 19591 2234 19600 2268
rect 19600 2234 19634 2268
rect 19634 2234 19643 2268
rect 19591 2225 19643 2234
rect 21223 2268 21275 2277
rect 21223 2234 21232 2268
rect 21232 2234 21266 2268
rect 21266 2234 21275 2268
rect 21223 2225 21275 2234
rect 22855 2268 22907 2277
rect 22855 2234 22864 2268
rect 22864 2234 22898 2268
rect 22898 2234 22907 2268
rect 22855 2225 22907 2234
rect 24487 2268 24539 2277
rect 24487 2234 24496 2268
rect 24496 2234 24530 2268
rect 24530 2234 24539 2268
rect 24487 2225 24539 2234
rect 26119 2268 26171 2277
rect 26119 2234 26128 2268
rect 26128 2234 26162 2268
rect 26162 2234 26171 2268
rect 26119 2225 26171 2234
rect 27751 2268 27803 2277
rect 27751 2234 27760 2268
rect 27760 2234 27794 2268
rect 27794 2234 27803 2268
rect 27751 2225 27803 2234
rect 29383 2268 29435 2277
rect 29383 2234 29392 2268
rect 29392 2234 29426 2268
rect 29426 2234 29435 2268
rect 29383 2225 29435 2234
rect 31015 2268 31067 2277
rect 31015 2234 31024 2268
rect 31024 2234 31058 2268
rect 31058 2234 31067 2268
rect 31015 2225 31067 2234
rect 32647 2268 32699 2277
rect 32647 2234 32656 2268
rect 32656 2234 32690 2268
rect 32690 2234 32699 2268
rect 32647 2225 32699 2234
rect 34279 2268 34331 2277
rect 34279 2234 34288 2268
rect 34288 2234 34322 2268
rect 34322 2234 34331 2268
rect 34279 2225 34331 2234
rect 35911 2268 35963 2277
rect 35911 2234 35920 2268
rect 35920 2234 35954 2268
rect 35954 2234 35963 2268
rect 35911 2225 35963 2234
rect 37543 2268 37595 2277
rect 37543 2234 37552 2268
rect 37552 2234 37586 2268
rect 37586 2234 37595 2268
rect 37543 2225 37595 2234
rect 39175 2268 39227 2277
rect 39175 2234 39184 2268
rect 39184 2234 39218 2268
rect 39218 2234 39227 2268
rect 39175 2225 39227 2234
rect 40807 2268 40859 2277
rect 40807 2234 40816 2268
rect 40816 2234 40850 2268
rect 40850 2234 40859 2268
rect 40807 2225 40859 2234
rect 42439 2268 42491 2277
rect 42439 2234 42448 2268
rect 42448 2234 42482 2268
rect 42482 2234 42491 2268
rect 42439 2225 42491 2234
rect 44071 2268 44123 2277
rect 44071 2234 44080 2268
rect 44080 2234 44114 2268
rect 44114 2234 44123 2268
rect 44071 2225 44123 2234
rect 45703 2268 45755 2277
rect 45703 2234 45712 2268
rect 45712 2234 45746 2268
rect 45746 2234 45755 2268
rect 45703 2225 45755 2234
rect 47335 2268 47387 2277
rect 47335 2234 47344 2268
rect 47344 2234 47378 2268
rect 47378 2234 47387 2268
rect 47335 2225 47387 2234
rect 48967 2268 49019 2277
rect 48967 2234 48976 2268
rect 48976 2234 49010 2268
rect 49010 2234 49019 2268
rect 48967 2225 49019 2234
rect 50599 2268 50651 2277
rect 50599 2234 50608 2268
rect 50608 2234 50642 2268
rect 50642 2234 50651 2268
rect 50599 2225 50651 2234
rect 52231 2268 52283 2277
rect 52231 2234 52240 2268
rect 52240 2234 52274 2268
rect 52274 2234 52283 2268
rect 52231 2225 52283 2234
rect 7 2064 59 2073
rect 7 2030 16 2064
rect 16 2030 50 2064
rect 50 2030 59 2064
rect 7 2021 59 2030
rect 1639 2064 1691 2073
rect 1639 2030 1648 2064
rect 1648 2030 1682 2064
rect 1682 2030 1691 2064
rect 1639 2021 1691 2030
rect 3271 2064 3323 2073
rect 3271 2030 3280 2064
rect 3280 2030 3314 2064
rect 3314 2030 3323 2064
rect 3271 2021 3323 2030
rect 4903 2064 4955 2073
rect 4903 2030 4912 2064
rect 4912 2030 4946 2064
rect 4946 2030 4955 2064
rect 4903 2021 4955 2030
rect 6535 2064 6587 2073
rect 6535 2030 6544 2064
rect 6544 2030 6578 2064
rect 6578 2030 6587 2064
rect 6535 2021 6587 2030
rect 8167 2064 8219 2073
rect 8167 2030 8176 2064
rect 8176 2030 8210 2064
rect 8210 2030 8219 2064
rect 8167 2021 8219 2030
rect 9799 2064 9851 2073
rect 9799 2030 9808 2064
rect 9808 2030 9842 2064
rect 9842 2030 9851 2064
rect 9799 2021 9851 2030
rect 11431 2064 11483 2073
rect 11431 2030 11440 2064
rect 11440 2030 11474 2064
rect 11474 2030 11483 2064
rect 11431 2021 11483 2030
rect 13063 2064 13115 2073
rect 13063 2030 13072 2064
rect 13072 2030 13106 2064
rect 13106 2030 13115 2064
rect 13063 2021 13115 2030
rect 14695 2064 14747 2073
rect 14695 2030 14704 2064
rect 14704 2030 14738 2064
rect 14738 2030 14747 2064
rect 14695 2021 14747 2030
rect 16327 2064 16379 2073
rect 16327 2030 16336 2064
rect 16336 2030 16370 2064
rect 16370 2030 16379 2064
rect 16327 2021 16379 2030
rect 17959 2064 18011 2073
rect 17959 2030 17968 2064
rect 17968 2030 18002 2064
rect 18002 2030 18011 2064
rect 17959 2021 18011 2030
rect 19591 2064 19643 2073
rect 19591 2030 19600 2064
rect 19600 2030 19634 2064
rect 19634 2030 19643 2064
rect 19591 2021 19643 2030
rect 21223 2064 21275 2073
rect 21223 2030 21232 2064
rect 21232 2030 21266 2064
rect 21266 2030 21275 2064
rect 21223 2021 21275 2030
rect 22855 2064 22907 2073
rect 22855 2030 22864 2064
rect 22864 2030 22898 2064
rect 22898 2030 22907 2064
rect 22855 2021 22907 2030
rect 24487 2064 24539 2073
rect 24487 2030 24496 2064
rect 24496 2030 24530 2064
rect 24530 2030 24539 2064
rect 24487 2021 24539 2030
rect 26119 2064 26171 2073
rect 26119 2030 26128 2064
rect 26128 2030 26162 2064
rect 26162 2030 26171 2064
rect 26119 2021 26171 2030
rect 27751 2064 27803 2073
rect 27751 2030 27760 2064
rect 27760 2030 27794 2064
rect 27794 2030 27803 2064
rect 27751 2021 27803 2030
rect 29383 2064 29435 2073
rect 29383 2030 29392 2064
rect 29392 2030 29426 2064
rect 29426 2030 29435 2064
rect 29383 2021 29435 2030
rect 31015 2064 31067 2073
rect 31015 2030 31024 2064
rect 31024 2030 31058 2064
rect 31058 2030 31067 2064
rect 31015 2021 31067 2030
rect 32647 2064 32699 2073
rect 32647 2030 32656 2064
rect 32656 2030 32690 2064
rect 32690 2030 32699 2064
rect 32647 2021 32699 2030
rect 34279 2064 34331 2073
rect 34279 2030 34288 2064
rect 34288 2030 34322 2064
rect 34322 2030 34331 2064
rect 34279 2021 34331 2030
rect 35911 2064 35963 2073
rect 35911 2030 35920 2064
rect 35920 2030 35954 2064
rect 35954 2030 35963 2064
rect 35911 2021 35963 2030
rect 37543 2064 37595 2073
rect 37543 2030 37552 2064
rect 37552 2030 37586 2064
rect 37586 2030 37595 2064
rect 37543 2021 37595 2030
rect 39175 2064 39227 2073
rect 39175 2030 39184 2064
rect 39184 2030 39218 2064
rect 39218 2030 39227 2064
rect 39175 2021 39227 2030
rect 40807 2064 40859 2073
rect 40807 2030 40816 2064
rect 40816 2030 40850 2064
rect 40850 2030 40859 2064
rect 40807 2021 40859 2030
rect 42439 2064 42491 2073
rect 42439 2030 42448 2064
rect 42448 2030 42482 2064
rect 42482 2030 42491 2064
rect 42439 2021 42491 2030
rect 44071 2064 44123 2073
rect 44071 2030 44080 2064
rect 44080 2030 44114 2064
rect 44114 2030 44123 2064
rect 44071 2021 44123 2030
rect 45703 2064 45755 2073
rect 45703 2030 45712 2064
rect 45712 2030 45746 2064
rect 45746 2030 45755 2064
rect 45703 2021 45755 2030
rect 47335 2064 47387 2073
rect 47335 2030 47344 2064
rect 47344 2030 47378 2064
rect 47378 2030 47387 2064
rect 47335 2021 47387 2030
rect 48967 2064 49019 2073
rect 48967 2030 48976 2064
rect 48976 2030 49010 2064
rect 49010 2030 49019 2064
rect 48967 2021 49019 2030
rect 50599 2064 50651 2073
rect 50599 2030 50608 2064
rect 50608 2030 50642 2064
rect 50642 2030 50651 2064
rect 50599 2021 50651 2030
rect 52231 2064 52283 2073
rect 52231 2030 52240 2064
rect 52240 2030 52274 2064
rect 52274 2030 52283 2064
rect 52231 2021 52283 2030
rect 7 1860 59 1869
rect 7 1826 16 1860
rect 16 1826 50 1860
rect 50 1826 59 1860
rect 7 1817 59 1826
rect 1639 1860 1691 1869
rect 1639 1826 1648 1860
rect 1648 1826 1682 1860
rect 1682 1826 1691 1860
rect 1639 1817 1691 1826
rect 3271 1860 3323 1869
rect 3271 1826 3280 1860
rect 3280 1826 3314 1860
rect 3314 1826 3323 1860
rect 3271 1817 3323 1826
rect 4903 1860 4955 1869
rect 4903 1826 4912 1860
rect 4912 1826 4946 1860
rect 4946 1826 4955 1860
rect 4903 1817 4955 1826
rect 6535 1860 6587 1869
rect 6535 1826 6544 1860
rect 6544 1826 6578 1860
rect 6578 1826 6587 1860
rect 6535 1817 6587 1826
rect 8167 1860 8219 1869
rect 8167 1826 8176 1860
rect 8176 1826 8210 1860
rect 8210 1826 8219 1860
rect 8167 1817 8219 1826
rect 9799 1860 9851 1869
rect 9799 1826 9808 1860
rect 9808 1826 9842 1860
rect 9842 1826 9851 1860
rect 9799 1817 9851 1826
rect 11431 1860 11483 1869
rect 11431 1826 11440 1860
rect 11440 1826 11474 1860
rect 11474 1826 11483 1860
rect 11431 1817 11483 1826
rect 13063 1860 13115 1869
rect 13063 1826 13072 1860
rect 13072 1826 13106 1860
rect 13106 1826 13115 1860
rect 13063 1817 13115 1826
rect 14695 1860 14747 1869
rect 14695 1826 14704 1860
rect 14704 1826 14738 1860
rect 14738 1826 14747 1860
rect 14695 1817 14747 1826
rect 16327 1860 16379 1869
rect 16327 1826 16336 1860
rect 16336 1826 16370 1860
rect 16370 1826 16379 1860
rect 16327 1817 16379 1826
rect 17959 1860 18011 1869
rect 17959 1826 17968 1860
rect 17968 1826 18002 1860
rect 18002 1826 18011 1860
rect 17959 1817 18011 1826
rect 19591 1860 19643 1869
rect 19591 1826 19600 1860
rect 19600 1826 19634 1860
rect 19634 1826 19643 1860
rect 19591 1817 19643 1826
rect 21223 1860 21275 1869
rect 21223 1826 21232 1860
rect 21232 1826 21266 1860
rect 21266 1826 21275 1860
rect 21223 1817 21275 1826
rect 22855 1860 22907 1869
rect 22855 1826 22864 1860
rect 22864 1826 22898 1860
rect 22898 1826 22907 1860
rect 22855 1817 22907 1826
rect 24487 1860 24539 1869
rect 24487 1826 24496 1860
rect 24496 1826 24530 1860
rect 24530 1826 24539 1860
rect 24487 1817 24539 1826
rect 26119 1860 26171 1869
rect 26119 1826 26128 1860
rect 26128 1826 26162 1860
rect 26162 1826 26171 1860
rect 26119 1817 26171 1826
rect 27751 1860 27803 1869
rect 27751 1826 27760 1860
rect 27760 1826 27794 1860
rect 27794 1826 27803 1860
rect 27751 1817 27803 1826
rect 29383 1860 29435 1869
rect 29383 1826 29392 1860
rect 29392 1826 29426 1860
rect 29426 1826 29435 1860
rect 29383 1817 29435 1826
rect 31015 1860 31067 1869
rect 31015 1826 31024 1860
rect 31024 1826 31058 1860
rect 31058 1826 31067 1860
rect 31015 1817 31067 1826
rect 32647 1860 32699 1869
rect 32647 1826 32656 1860
rect 32656 1826 32690 1860
rect 32690 1826 32699 1860
rect 32647 1817 32699 1826
rect 34279 1860 34331 1869
rect 34279 1826 34288 1860
rect 34288 1826 34322 1860
rect 34322 1826 34331 1860
rect 34279 1817 34331 1826
rect 35911 1860 35963 1869
rect 35911 1826 35920 1860
rect 35920 1826 35954 1860
rect 35954 1826 35963 1860
rect 35911 1817 35963 1826
rect 37543 1860 37595 1869
rect 37543 1826 37552 1860
rect 37552 1826 37586 1860
rect 37586 1826 37595 1860
rect 37543 1817 37595 1826
rect 39175 1860 39227 1869
rect 39175 1826 39184 1860
rect 39184 1826 39218 1860
rect 39218 1826 39227 1860
rect 39175 1817 39227 1826
rect 40807 1860 40859 1869
rect 40807 1826 40816 1860
rect 40816 1826 40850 1860
rect 40850 1826 40859 1860
rect 40807 1817 40859 1826
rect 42439 1860 42491 1869
rect 42439 1826 42448 1860
rect 42448 1826 42482 1860
rect 42482 1826 42491 1860
rect 42439 1817 42491 1826
rect 44071 1860 44123 1869
rect 44071 1826 44080 1860
rect 44080 1826 44114 1860
rect 44114 1826 44123 1860
rect 44071 1817 44123 1826
rect 45703 1860 45755 1869
rect 45703 1826 45712 1860
rect 45712 1826 45746 1860
rect 45746 1826 45755 1860
rect 45703 1817 45755 1826
rect 47335 1860 47387 1869
rect 47335 1826 47344 1860
rect 47344 1826 47378 1860
rect 47378 1826 47387 1860
rect 47335 1817 47387 1826
rect 48967 1860 49019 1869
rect 48967 1826 48976 1860
rect 48976 1826 49010 1860
rect 49010 1826 49019 1860
rect 48967 1817 49019 1826
rect 50599 1860 50651 1869
rect 50599 1826 50608 1860
rect 50608 1826 50642 1860
rect 50642 1826 50651 1860
rect 50599 1817 50651 1826
rect 52231 1860 52283 1869
rect 52231 1826 52240 1860
rect 52240 1826 52274 1860
rect 52274 1826 52283 1860
rect 52231 1817 52283 1826
rect 7 1656 59 1665
rect 7 1622 16 1656
rect 16 1622 50 1656
rect 50 1622 59 1656
rect 7 1613 59 1622
rect 1639 1656 1691 1665
rect 1639 1622 1648 1656
rect 1648 1622 1682 1656
rect 1682 1622 1691 1656
rect 1639 1613 1691 1622
rect 3271 1656 3323 1665
rect 3271 1622 3280 1656
rect 3280 1622 3314 1656
rect 3314 1622 3323 1656
rect 3271 1613 3323 1622
rect 4903 1656 4955 1665
rect 4903 1622 4912 1656
rect 4912 1622 4946 1656
rect 4946 1622 4955 1656
rect 4903 1613 4955 1622
rect 6535 1656 6587 1665
rect 6535 1622 6544 1656
rect 6544 1622 6578 1656
rect 6578 1622 6587 1656
rect 6535 1613 6587 1622
rect 8167 1656 8219 1665
rect 8167 1622 8176 1656
rect 8176 1622 8210 1656
rect 8210 1622 8219 1656
rect 8167 1613 8219 1622
rect 9799 1656 9851 1665
rect 9799 1622 9808 1656
rect 9808 1622 9842 1656
rect 9842 1622 9851 1656
rect 9799 1613 9851 1622
rect 11431 1656 11483 1665
rect 11431 1622 11440 1656
rect 11440 1622 11474 1656
rect 11474 1622 11483 1656
rect 11431 1613 11483 1622
rect 13063 1656 13115 1665
rect 13063 1622 13072 1656
rect 13072 1622 13106 1656
rect 13106 1622 13115 1656
rect 13063 1613 13115 1622
rect 14695 1656 14747 1665
rect 14695 1622 14704 1656
rect 14704 1622 14738 1656
rect 14738 1622 14747 1656
rect 14695 1613 14747 1622
rect 16327 1656 16379 1665
rect 16327 1622 16336 1656
rect 16336 1622 16370 1656
rect 16370 1622 16379 1656
rect 16327 1613 16379 1622
rect 17959 1656 18011 1665
rect 17959 1622 17968 1656
rect 17968 1622 18002 1656
rect 18002 1622 18011 1656
rect 17959 1613 18011 1622
rect 19591 1656 19643 1665
rect 19591 1622 19600 1656
rect 19600 1622 19634 1656
rect 19634 1622 19643 1656
rect 19591 1613 19643 1622
rect 21223 1656 21275 1665
rect 21223 1622 21232 1656
rect 21232 1622 21266 1656
rect 21266 1622 21275 1656
rect 21223 1613 21275 1622
rect 22855 1656 22907 1665
rect 22855 1622 22864 1656
rect 22864 1622 22898 1656
rect 22898 1622 22907 1656
rect 22855 1613 22907 1622
rect 24487 1656 24539 1665
rect 24487 1622 24496 1656
rect 24496 1622 24530 1656
rect 24530 1622 24539 1656
rect 24487 1613 24539 1622
rect 26119 1656 26171 1665
rect 26119 1622 26128 1656
rect 26128 1622 26162 1656
rect 26162 1622 26171 1656
rect 26119 1613 26171 1622
rect 27751 1656 27803 1665
rect 27751 1622 27760 1656
rect 27760 1622 27794 1656
rect 27794 1622 27803 1656
rect 27751 1613 27803 1622
rect 29383 1656 29435 1665
rect 29383 1622 29392 1656
rect 29392 1622 29426 1656
rect 29426 1622 29435 1656
rect 29383 1613 29435 1622
rect 31015 1656 31067 1665
rect 31015 1622 31024 1656
rect 31024 1622 31058 1656
rect 31058 1622 31067 1656
rect 31015 1613 31067 1622
rect 32647 1656 32699 1665
rect 32647 1622 32656 1656
rect 32656 1622 32690 1656
rect 32690 1622 32699 1656
rect 32647 1613 32699 1622
rect 34279 1656 34331 1665
rect 34279 1622 34288 1656
rect 34288 1622 34322 1656
rect 34322 1622 34331 1656
rect 34279 1613 34331 1622
rect 35911 1656 35963 1665
rect 35911 1622 35920 1656
rect 35920 1622 35954 1656
rect 35954 1622 35963 1656
rect 35911 1613 35963 1622
rect 37543 1656 37595 1665
rect 37543 1622 37552 1656
rect 37552 1622 37586 1656
rect 37586 1622 37595 1656
rect 37543 1613 37595 1622
rect 39175 1656 39227 1665
rect 39175 1622 39184 1656
rect 39184 1622 39218 1656
rect 39218 1622 39227 1656
rect 39175 1613 39227 1622
rect 40807 1656 40859 1665
rect 40807 1622 40816 1656
rect 40816 1622 40850 1656
rect 40850 1622 40859 1656
rect 40807 1613 40859 1622
rect 42439 1656 42491 1665
rect 42439 1622 42448 1656
rect 42448 1622 42482 1656
rect 42482 1622 42491 1656
rect 42439 1613 42491 1622
rect 44071 1656 44123 1665
rect 44071 1622 44080 1656
rect 44080 1622 44114 1656
rect 44114 1622 44123 1656
rect 44071 1613 44123 1622
rect 45703 1656 45755 1665
rect 45703 1622 45712 1656
rect 45712 1622 45746 1656
rect 45746 1622 45755 1656
rect 45703 1613 45755 1622
rect 47335 1656 47387 1665
rect 47335 1622 47344 1656
rect 47344 1622 47378 1656
rect 47378 1622 47387 1656
rect 47335 1613 47387 1622
rect 48967 1656 49019 1665
rect 48967 1622 48976 1656
rect 48976 1622 49010 1656
rect 49010 1622 49019 1656
rect 48967 1613 49019 1622
rect 50599 1656 50651 1665
rect 50599 1622 50608 1656
rect 50608 1622 50642 1656
rect 50642 1622 50651 1656
rect 50599 1613 50651 1622
rect 52231 1656 52283 1665
rect 52231 1622 52240 1656
rect 52240 1622 52274 1656
rect 52274 1622 52283 1656
rect 52231 1613 52283 1622
rect 7 1452 59 1461
rect 7 1418 16 1452
rect 16 1418 50 1452
rect 50 1418 59 1452
rect 7 1409 59 1418
rect 1639 1452 1691 1461
rect 1639 1418 1648 1452
rect 1648 1418 1682 1452
rect 1682 1418 1691 1452
rect 1639 1409 1691 1418
rect 3271 1452 3323 1461
rect 3271 1418 3280 1452
rect 3280 1418 3314 1452
rect 3314 1418 3323 1452
rect 3271 1409 3323 1418
rect 4903 1452 4955 1461
rect 4903 1418 4912 1452
rect 4912 1418 4946 1452
rect 4946 1418 4955 1452
rect 4903 1409 4955 1418
rect 6535 1452 6587 1461
rect 6535 1418 6544 1452
rect 6544 1418 6578 1452
rect 6578 1418 6587 1452
rect 6535 1409 6587 1418
rect 8167 1452 8219 1461
rect 8167 1418 8176 1452
rect 8176 1418 8210 1452
rect 8210 1418 8219 1452
rect 8167 1409 8219 1418
rect 9799 1452 9851 1461
rect 9799 1418 9808 1452
rect 9808 1418 9842 1452
rect 9842 1418 9851 1452
rect 9799 1409 9851 1418
rect 11431 1452 11483 1461
rect 11431 1418 11440 1452
rect 11440 1418 11474 1452
rect 11474 1418 11483 1452
rect 11431 1409 11483 1418
rect 13063 1452 13115 1461
rect 13063 1418 13072 1452
rect 13072 1418 13106 1452
rect 13106 1418 13115 1452
rect 13063 1409 13115 1418
rect 14695 1452 14747 1461
rect 14695 1418 14704 1452
rect 14704 1418 14738 1452
rect 14738 1418 14747 1452
rect 14695 1409 14747 1418
rect 16327 1452 16379 1461
rect 16327 1418 16336 1452
rect 16336 1418 16370 1452
rect 16370 1418 16379 1452
rect 16327 1409 16379 1418
rect 17959 1452 18011 1461
rect 17959 1418 17968 1452
rect 17968 1418 18002 1452
rect 18002 1418 18011 1452
rect 17959 1409 18011 1418
rect 19591 1452 19643 1461
rect 19591 1418 19600 1452
rect 19600 1418 19634 1452
rect 19634 1418 19643 1452
rect 19591 1409 19643 1418
rect 21223 1452 21275 1461
rect 21223 1418 21232 1452
rect 21232 1418 21266 1452
rect 21266 1418 21275 1452
rect 21223 1409 21275 1418
rect 22855 1452 22907 1461
rect 22855 1418 22864 1452
rect 22864 1418 22898 1452
rect 22898 1418 22907 1452
rect 22855 1409 22907 1418
rect 24487 1452 24539 1461
rect 24487 1418 24496 1452
rect 24496 1418 24530 1452
rect 24530 1418 24539 1452
rect 24487 1409 24539 1418
rect 26119 1452 26171 1461
rect 26119 1418 26128 1452
rect 26128 1418 26162 1452
rect 26162 1418 26171 1452
rect 26119 1409 26171 1418
rect 27751 1452 27803 1461
rect 27751 1418 27760 1452
rect 27760 1418 27794 1452
rect 27794 1418 27803 1452
rect 27751 1409 27803 1418
rect 29383 1452 29435 1461
rect 29383 1418 29392 1452
rect 29392 1418 29426 1452
rect 29426 1418 29435 1452
rect 29383 1409 29435 1418
rect 31015 1452 31067 1461
rect 31015 1418 31024 1452
rect 31024 1418 31058 1452
rect 31058 1418 31067 1452
rect 31015 1409 31067 1418
rect 32647 1452 32699 1461
rect 32647 1418 32656 1452
rect 32656 1418 32690 1452
rect 32690 1418 32699 1452
rect 32647 1409 32699 1418
rect 34279 1452 34331 1461
rect 34279 1418 34288 1452
rect 34288 1418 34322 1452
rect 34322 1418 34331 1452
rect 34279 1409 34331 1418
rect 35911 1452 35963 1461
rect 35911 1418 35920 1452
rect 35920 1418 35954 1452
rect 35954 1418 35963 1452
rect 35911 1409 35963 1418
rect 37543 1452 37595 1461
rect 37543 1418 37552 1452
rect 37552 1418 37586 1452
rect 37586 1418 37595 1452
rect 37543 1409 37595 1418
rect 39175 1452 39227 1461
rect 39175 1418 39184 1452
rect 39184 1418 39218 1452
rect 39218 1418 39227 1452
rect 39175 1409 39227 1418
rect 40807 1452 40859 1461
rect 40807 1418 40816 1452
rect 40816 1418 40850 1452
rect 40850 1418 40859 1452
rect 40807 1409 40859 1418
rect 42439 1452 42491 1461
rect 42439 1418 42448 1452
rect 42448 1418 42482 1452
rect 42482 1418 42491 1452
rect 42439 1409 42491 1418
rect 44071 1452 44123 1461
rect 44071 1418 44080 1452
rect 44080 1418 44114 1452
rect 44114 1418 44123 1452
rect 44071 1409 44123 1418
rect 45703 1452 45755 1461
rect 45703 1418 45712 1452
rect 45712 1418 45746 1452
rect 45746 1418 45755 1452
rect 45703 1409 45755 1418
rect 47335 1452 47387 1461
rect 47335 1418 47344 1452
rect 47344 1418 47378 1452
rect 47378 1418 47387 1452
rect 47335 1409 47387 1418
rect 48967 1452 49019 1461
rect 48967 1418 48976 1452
rect 48976 1418 49010 1452
rect 49010 1418 49019 1452
rect 48967 1409 49019 1418
rect 50599 1452 50651 1461
rect 50599 1418 50608 1452
rect 50608 1418 50642 1452
rect 50642 1418 50651 1452
rect 50599 1409 50651 1418
rect 52231 1452 52283 1461
rect 52231 1418 52240 1452
rect 52240 1418 52274 1452
rect 52274 1418 52283 1452
rect 52231 1409 52283 1418
rect 7 1248 59 1257
rect 7 1214 16 1248
rect 16 1214 50 1248
rect 50 1214 59 1248
rect 7 1205 59 1214
rect 1639 1248 1691 1257
rect 1639 1214 1648 1248
rect 1648 1214 1682 1248
rect 1682 1214 1691 1248
rect 1639 1205 1691 1214
rect 3271 1248 3323 1257
rect 3271 1214 3280 1248
rect 3280 1214 3314 1248
rect 3314 1214 3323 1248
rect 3271 1205 3323 1214
rect 4903 1248 4955 1257
rect 4903 1214 4912 1248
rect 4912 1214 4946 1248
rect 4946 1214 4955 1248
rect 4903 1205 4955 1214
rect 6535 1248 6587 1257
rect 6535 1214 6544 1248
rect 6544 1214 6578 1248
rect 6578 1214 6587 1248
rect 6535 1205 6587 1214
rect 8167 1248 8219 1257
rect 8167 1214 8176 1248
rect 8176 1214 8210 1248
rect 8210 1214 8219 1248
rect 8167 1205 8219 1214
rect 9799 1248 9851 1257
rect 9799 1214 9808 1248
rect 9808 1214 9842 1248
rect 9842 1214 9851 1248
rect 9799 1205 9851 1214
rect 11431 1248 11483 1257
rect 11431 1214 11440 1248
rect 11440 1214 11474 1248
rect 11474 1214 11483 1248
rect 11431 1205 11483 1214
rect 13063 1248 13115 1257
rect 13063 1214 13072 1248
rect 13072 1214 13106 1248
rect 13106 1214 13115 1248
rect 13063 1205 13115 1214
rect 14695 1248 14747 1257
rect 14695 1214 14704 1248
rect 14704 1214 14738 1248
rect 14738 1214 14747 1248
rect 14695 1205 14747 1214
rect 16327 1248 16379 1257
rect 16327 1214 16336 1248
rect 16336 1214 16370 1248
rect 16370 1214 16379 1248
rect 16327 1205 16379 1214
rect 17959 1248 18011 1257
rect 17959 1214 17968 1248
rect 17968 1214 18002 1248
rect 18002 1214 18011 1248
rect 17959 1205 18011 1214
rect 19591 1248 19643 1257
rect 19591 1214 19600 1248
rect 19600 1214 19634 1248
rect 19634 1214 19643 1248
rect 19591 1205 19643 1214
rect 21223 1248 21275 1257
rect 21223 1214 21232 1248
rect 21232 1214 21266 1248
rect 21266 1214 21275 1248
rect 21223 1205 21275 1214
rect 22855 1248 22907 1257
rect 22855 1214 22864 1248
rect 22864 1214 22898 1248
rect 22898 1214 22907 1248
rect 22855 1205 22907 1214
rect 24487 1248 24539 1257
rect 24487 1214 24496 1248
rect 24496 1214 24530 1248
rect 24530 1214 24539 1248
rect 24487 1205 24539 1214
rect 26119 1248 26171 1257
rect 26119 1214 26128 1248
rect 26128 1214 26162 1248
rect 26162 1214 26171 1248
rect 26119 1205 26171 1214
rect 27751 1248 27803 1257
rect 27751 1214 27760 1248
rect 27760 1214 27794 1248
rect 27794 1214 27803 1248
rect 27751 1205 27803 1214
rect 29383 1248 29435 1257
rect 29383 1214 29392 1248
rect 29392 1214 29426 1248
rect 29426 1214 29435 1248
rect 29383 1205 29435 1214
rect 31015 1248 31067 1257
rect 31015 1214 31024 1248
rect 31024 1214 31058 1248
rect 31058 1214 31067 1248
rect 31015 1205 31067 1214
rect 32647 1248 32699 1257
rect 32647 1214 32656 1248
rect 32656 1214 32690 1248
rect 32690 1214 32699 1248
rect 32647 1205 32699 1214
rect 34279 1248 34331 1257
rect 34279 1214 34288 1248
rect 34288 1214 34322 1248
rect 34322 1214 34331 1248
rect 34279 1205 34331 1214
rect 35911 1248 35963 1257
rect 35911 1214 35920 1248
rect 35920 1214 35954 1248
rect 35954 1214 35963 1248
rect 35911 1205 35963 1214
rect 37543 1248 37595 1257
rect 37543 1214 37552 1248
rect 37552 1214 37586 1248
rect 37586 1214 37595 1248
rect 37543 1205 37595 1214
rect 39175 1248 39227 1257
rect 39175 1214 39184 1248
rect 39184 1214 39218 1248
rect 39218 1214 39227 1248
rect 39175 1205 39227 1214
rect 40807 1248 40859 1257
rect 40807 1214 40816 1248
rect 40816 1214 40850 1248
rect 40850 1214 40859 1248
rect 40807 1205 40859 1214
rect 42439 1248 42491 1257
rect 42439 1214 42448 1248
rect 42448 1214 42482 1248
rect 42482 1214 42491 1248
rect 42439 1205 42491 1214
rect 44071 1248 44123 1257
rect 44071 1214 44080 1248
rect 44080 1214 44114 1248
rect 44114 1214 44123 1248
rect 44071 1205 44123 1214
rect 45703 1248 45755 1257
rect 45703 1214 45712 1248
rect 45712 1214 45746 1248
rect 45746 1214 45755 1248
rect 45703 1205 45755 1214
rect 47335 1248 47387 1257
rect 47335 1214 47344 1248
rect 47344 1214 47378 1248
rect 47378 1214 47387 1248
rect 47335 1205 47387 1214
rect 48967 1248 49019 1257
rect 48967 1214 48976 1248
rect 48976 1214 49010 1248
rect 49010 1214 49019 1248
rect 48967 1205 49019 1214
rect 50599 1248 50651 1257
rect 50599 1214 50608 1248
rect 50608 1214 50642 1248
rect 50642 1214 50651 1248
rect 50599 1205 50651 1214
rect 52231 1248 52283 1257
rect 52231 1214 52240 1248
rect 52240 1214 52274 1248
rect 52274 1214 52283 1248
rect 52231 1205 52283 1214
rect 7 1044 59 1053
rect 7 1010 16 1044
rect 16 1010 50 1044
rect 50 1010 59 1044
rect 7 1001 59 1010
rect 1639 1044 1691 1053
rect 1639 1010 1648 1044
rect 1648 1010 1682 1044
rect 1682 1010 1691 1044
rect 1639 1001 1691 1010
rect 3271 1044 3323 1053
rect 3271 1010 3280 1044
rect 3280 1010 3314 1044
rect 3314 1010 3323 1044
rect 3271 1001 3323 1010
rect 4903 1044 4955 1053
rect 4903 1010 4912 1044
rect 4912 1010 4946 1044
rect 4946 1010 4955 1044
rect 4903 1001 4955 1010
rect 6535 1044 6587 1053
rect 6535 1010 6544 1044
rect 6544 1010 6578 1044
rect 6578 1010 6587 1044
rect 6535 1001 6587 1010
rect 8167 1044 8219 1053
rect 8167 1010 8176 1044
rect 8176 1010 8210 1044
rect 8210 1010 8219 1044
rect 8167 1001 8219 1010
rect 9799 1044 9851 1053
rect 9799 1010 9808 1044
rect 9808 1010 9842 1044
rect 9842 1010 9851 1044
rect 9799 1001 9851 1010
rect 11431 1044 11483 1053
rect 11431 1010 11440 1044
rect 11440 1010 11474 1044
rect 11474 1010 11483 1044
rect 11431 1001 11483 1010
rect 13063 1044 13115 1053
rect 13063 1010 13072 1044
rect 13072 1010 13106 1044
rect 13106 1010 13115 1044
rect 13063 1001 13115 1010
rect 14695 1044 14747 1053
rect 14695 1010 14704 1044
rect 14704 1010 14738 1044
rect 14738 1010 14747 1044
rect 14695 1001 14747 1010
rect 16327 1044 16379 1053
rect 16327 1010 16336 1044
rect 16336 1010 16370 1044
rect 16370 1010 16379 1044
rect 16327 1001 16379 1010
rect 17959 1044 18011 1053
rect 17959 1010 17968 1044
rect 17968 1010 18002 1044
rect 18002 1010 18011 1044
rect 17959 1001 18011 1010
rect 19591 1044 19643 1053
rect 19591 1010 19600 1044
rect 19600 1010 19634 1044
rect 19634 1010 19643 1044
rect 19591 1001 19643 1010
rect 21223 1044 21275 1053
rect 21223 1010 21232 1044
rect 21232 1010 21266 1044
rect 21266 1010 21275 1044
rect 21223 1001 21275 1010
rect 22855 1044 22907 1053
rect 22855 1010 22864 1044
rect 22864 1010 22898 1044
rect 22898 1010 22907 1044
rect 22855 1001 22907 1010
rect 24487 1044 24539 1053
rect 24487 1010 24496 1044
rect 24496 1010 24530 1044
rect 24530 1010 24539 1044
rect 24487 1001 24539 1010
rect 26119 1044 26171 1053
rect 26119 1010 26128 1044
rect 26128 1010 26162 1044
rect 26162 1010 26171 1044
rect 26119 1001 26171 1010
rect 27751 1044 27803 1053
rect 27751 1010 27760 1044
rect 27760 1010 27794 1044
rect 27794 1010 27803 1044
rect 27751 1001 27803 1010
rect 29383 1044 29435 1053
rect 29383 1010 29392 1044
rect 29392 1010 29426 1044
rect 29426 1010 29435 1044
rect 29383 1001 29435 1010
rect 31015 1044 31067 1053
rect 31015 1010 31024 1044
rect 31024 1010 31058 1044
rect 31058 1010 31067 1044
rect 31015 1001 31067 1010
rect 32647 1044 32699 1053
rect 32647 1010 32656 1044
rect 32656 1010 32690 1044
rect 32690 1010 32699 1044
rect 32647 1001 32699 1010
rect 34279 1044 34331 1053
rect 34279 1010 34288 1044
rect 34288 1010 34322 1044
rect 34322 1010 34331 1044
rect 34279 1001 34331 1010
rect 35911 1044 35963 1053
rect 35911 1010 35920 1044
rect 35920 1010 35954 1044
rect 35954 1010 35963 1044
rect 35911 1001 35963 1010
rect 37543 1044 37595 1053
rect 37543 1010 37552 1044
rect 37552 1010 37586 1044
rect 37586 1010 37595 1044
rect 37543 1001 37595 1010
rect 39175 1044 39227 1053
rect 39175 1010 39184 1044
rect 39184 1010 39218 1044
rect 39218 1010 39227 1044
rect 39175 1001 39227 1010
rect 40807 1044 40859 1053
rect 40807 1010 40816 1044
rect 40816 1010 40850 1044
rect 40850 1010 40859 1044
rect 40807 1001 40859 1010
rect 42439 1044 42491 1053
rect 42439 1010 42448 1044
rect 42448 1010 42482 1044
rect 42482 1010 42491 1044
rect 42439 1001 42491 1010
rect 44071 1044 44123 1053
rect 44071 1010 44080 1044
rect 44080 1010 44114 1044
rect 44114 1010 44123 1044
rect 44071 1001 44123 1010
rect 45703 1044 45755 1053
rect 45703 1010 45712 1044
rect 45712 1010 45746 1044
rect 45746 1010 45755 1044
rect 45703 1001 45755 1010
rect 47335 1044 47387 1053
rect 47335 1010 47344 1044
rect 47344 1010 47378 1044
rect 47378 1010 47387 1044
rect 47335 1001 47387 1010
rect 48967 1044 49019 1053
rect 48967 1010 48976 1044
rect 48976 1010 49010 1044
rect 49010 1010 49019 1044
rect 48967 1001 49019 1010
rect 50599 1044 50651 1053
rect 50599 1010 50608 1044
rect 50608 1010 50642 1044
rect 50642 1010 50651 1044
rect 50599 1001 50651 1010
rect 52231 1044 52283 1053
rect 52231 1010 52240 1044
rect 52240 1010 52274 1044
rect 52274 1010 52283 1044
rect 52231 1001 52283 1010
rect 218 890 270 899
rect 218 856 227 890
rect 227 856 261 890
rect 261 856 270 890
rect 218 847 270 856
rect 422 890 474 899
rect 422 856 431 890
rect 431 856 465 890
rect 465 856 474 890
rect 422 847 474 856
rect 626 890 678 899
rect 626 856 635 890
rect 635 856 669 890
rect 669 856 678 890
rect 626 847 678 856
rect 830 890 882 899
rect 830 856 839 890
rect 839 856 873 890
rect 873 856 882 890
rect 830 847 882 856
rect 1034 890 1086 899
rect 1034 856 1043 890
rect 1043 856 1077 890
rect 1077 856 1086 890
rect 1034 847 1086 856
rect 1238 890 1290 899
rect 1238 856 1247 890
rect 1247 856 1281 890
rect 1281 856 1290 890
rect 1238 847 1290 856
rect 1442 890 1494 899
rect 1442 856 1451 890
rect 1451 856 1485 890
rect 1485 856 1494 890
rect 1442 847 1494 856
rect 1646 890 1698 899
rect 1646 856 1655 890
rect 1655 856 1689 890
rect 1689 856 1698 890
rect 1646 847 1698 856
rect 1850 890 1902 899
rect 1850 856 1859 890
rect 1859 856 1893 890
rect 1893 856 1902 890
rect 1850 847 1902 856
rect 2054 890 2106 899
rect 2054 856 2063 890
rect 2063 856 2097 890
rect 2097 856 2106 890
rect 2054 847 2106 856
rect 2258 890 2310 899
rect 2258 856 2267 890
rect 2267 856 2301 890
rect 2301 856 2310 890
rect 2258 847 2310 856
rect 2462 890 2514 899
rect 2462 856 2471 890
rect 2471 856 2505 890
rect 2505 856 2514 890
rect 2462 847 2514 856
rect 2666 890 2718 899
rect 2666 856 2675 890
rect 2675 856 2709 890
rect 2709 856 2718 890
rect 2666 847 2718 856
rect 2870 890 2922 899
rect 2870 856 2879 890
rect 2879 856 2913 890
rect 2913 856 2922 890
rect 2870 847 2922 856
rect 3074 890 3126 899
rect 3074 856 3083 890
rect 3083 856 3117 890
rect 3117 856 3126 890
rect 3074 847 3126 856
rect 3278 890 3330 899
rect 3278 856 3287 890
rect 3287 856 3321 890
rect 3321 856 3330 890
rect 3278 847 3330 856
rect 3482 890 3534 899
rect 3482 856 3491 890
rect 3491 856 3525 890
rect 3525 856 3534 890
rect 3482 847 3534 856
rect 3686 890 3738 899
rect 3686 856 3695 890
rect 3695 856 3729 890
rect 3729 856 3738 890
rect 3686 847 3738 856
rect 3890 890 3942 899
rect 3890 856 3899 890
rect 3899 856 3933 890
rect 3933 856 3942 890
rect 3890 847 3942 856
rect 4094 890 4146 899
rect 4094 856 4103 890
rect 4103 856 4137 890
rect 4137 856 4146 890
rect 4094 847 4146 856
rect 4298 890 4350 899
rect 4298 856 4307 890
rect 4307 856 4341 890
rect 4341 856 4350 890
rect 4298 847 4350 856
rect 4502 890 4554 899
rect 4502 856 4511 890
rect 4511 856 4545 890
rect 4545 856 4554 890
rect 4502 847 4554 856
rect 4706 890 4758 899
rect 4706 856 4715 890
rect 4715 856 4749 890
rect 4749 856 4758 890
rect 4706 847 4758 856
rect 4910 890 4962 899
rect 4910 856 4919 890
rect 4919 856 4953 890
rect 4953 856 4962 890
rect 4910 847 4962 856
rect 5114 890 5166 899
rect 5114 856 5123 890
rect 5123 856 5157 890
rect 5157 856 5166 890
rect 5114 847 5166 856
rect 5318 890 5370 899
rect 5318 856 5327 890
rect 5327 856 5361 890
rect 5361 856 5370 890
rect 5318 847 5370 856
rect 5522 890 5574 899
rect 5522 856 5531 890
rect 5531 856 5565 890
rect 5565 856 5574 890
rect 5522 847 5574 856
rect 5726 890 5778 899
rect 5726 856 5735 890
rect 5735 856 5769 890
rect 5769 856 5778 890
rect 5726 847 5778 856
rect 5930 890 5982 899
rect 5930 856 5939 890
rect 5939 856 5973 890
rect 5973 856 5982 890
rect 5930 847 5982 856
rect 6134 890 6186 899
rect 6134 856 6143 890
rect 6143 856 6177 890
rect 6177 856 6186 890
rect 6134 847 6186 856
rect 6338 890 6390 899
rect 6338 856 6347 890
rect 6347 856 6381 890
rect 6381 856 6390 890
rect 6338 847 6390 856
rect 6542 890 6594 899
rect 6542 856 6551 890
rect 6551 856 6585 890
rect 6585 856 6594 890
rect 6542 847 6594 856
rect 6746 890 6798 899
rect 6746 856 6755 890
rect 6755 856 6789 890
rect 6789 856 6798 890
rect 6746 847 6798 856
rect 6950 890 7002 899
rect 6950 856 6959 890
rect 6959 856 6993 890
rect 6993 856 7002 890
rect 6950 847 7002 856
rect 7154 890 7206 899
rect 7154 856 7163 890
rect 7163 856 7197 890
rect 7197 856 7206 890
rect 7154 847 7206 856
rect 7358 890 7410 899
rect 7358 856 7367 890
rect 7367 856 7401 890
rect 7401 856 7410 890
rect 7358 847 7410 856
rect 7562 890 7614 899
rect 7562 856 7571 890
rect 7571 856 7605 890
rect 7605 856 7614 890
rect 7562 847 7614 856
rect 7766 890 7818 899
rect 7766 856 7775 890
rect 7775 856 7809 890
rect 7809 856 7818 890
rect 7766 847 7818 856
rect 7970 890 8022 899
rect 7970 856 7979 890
rect 7979 856 8013 890
rect 8013 856 8022 890
rect 7970 847 8022 856
rect 8174 890 8226 899
rect 8174 856 8183 890
rect 8183 856 8217 890
rect 8217 856 8226 890
rect 8174 847 8226 856
rect 8378 890 8430 899
rect 8378 856 8387 890
rect 8387 856 8421 890
rect 8421 856 8430 890
rect 8378 847 8430 856
rect 8582 890 8634 899
rect 8582 856 8591 890
rect 8591 856 8625 890
rect 8625 856 8634 890
rect 8582 847 8634 856
rect 8786 890 8838 899
rect 8786 856 8795 890
rect 8795 856 8829 890
rect 8829 856 8838 890
rect 8786 847 8838 856
rect 8990 890 9042 899
rect 8990 856 8999 890
rect 8999 856 9033 890
rect 9033 856 9042 890
rect 8990 847 9042 856
rect 9194 890 9246 899
rect 9194 856 9203 890
rect 9203 856 9237 890
rect 9237 856 9246 890
rect 9194 847 9246 856
rect 9398 890 9450 899
rect 9398 856 9407 890
rect 9407 856 9441 890
rect 9441 856 9450 890
rect 9398 847 9450 856
rect 9602 890 9654 899
rect 9602 856 9611 890
rect 9611 856 9645 890
rect 9645 856 9654 890
rect 9602 847 9654 856
rect 9806 890 9858 899
rect 9806 856 9815 890
rect 9815 856 9849 890
rect 9849 856 9858 890
rect 9806 847 9858 856
rect 10010 890 10062 899
rect 10010 856 10019 890
rect 10019 856 10053 890
rect 10053 856 10062 890
rect 10010 847 10062 856
rect 10214 890 10266 899
rect 10214 856 10223 890
rect 10223 856 10257 890
rect 10257 856 10266 890
rect 10214 847 10266 856
rect 10418 890 10470 899
rect 10418 856 10427 890
rect 10427 856 10461 890
rect 10461 856 10470 890
rect 10418 847 10470 856
rect 10622 890 10674 899
rect 10622 856 10631 890
rect 10631 856 10665 890
rect 10665 856 10674 890
rect 10622 847 10674 856
rect 10826 890 10878 899
rect 10826 856 10835 890
rect 10835 856 10869 890
rect 10869 856 10878 890
rect 10826 847 10878 856
rect 11030 890 11082 899
rect 11030 856 11039 890
rect 11039 856 11073 890
rect 11073 856 11082 890
rect 11030 847 11082 856
rect 11234 890 11286 899
rect 11234 856 11243 890
rect 11243 856 11277 890
rect 11277 856 11286 890
rect 11234 847 11286 856
rect 11438 890 11490 899
rect 11438 856 11447 890
rect 11447 856 11481 890
rect 11481 856 11490 890
rect 11438 847 11490 856
rect 11642 890 11694 899
rect 11642 856 11651 890
rect 11651 856 11685 890
rect 11685 856 11694 890
rect 11642 847 11694 856
rect 11846 890 11898 899
rect 11846 856 11855 890
rect 11855 856 11889 890
rect 11889 856 11898 890
rect 11846 847 11898 856
rect 12050 890 12102 899
rect 12050 856 12059 890
rect 12059 856 12093 890
rect 12093 856 12102 890
rect 12050 847 12102 856
rect 12254 890 12306 899
rect 12254 856 12263 890
rect 12263 856 12297 890
rect 12297 856 12306 890
rect 12254 847 12306 856
rect 12458 890 12510 899
rect 12458 856 12467 890
rect 12467 856 12501 890
rect 12501 856 12510 890
rect 12458 847 12510 856
rect 12662 890 12714 899
rect 12662 856 12671 890
rect 12671 856 12705 890
rect 12705 856 12714 890
rect 12662 847 12714 856
rect 12866 890 12918 899
rect 12866 856 12875 890
rect 12875 856 12909 890
rect 12909 856 12918 890
rect 12866 847 12918 856
rect 13070 890 13122 899
rect 13070 856 13079 890
rect 13079 856 13113 890
rect 13113 856 13122 890
rect 13070 847 13122 856
rect 13274 890 13326 899
rect 13274 856 13283 890
rect 13283 856 13317 890
rect 13317 856 13326 890
rect 13274 847 13326 856
rect 13478 890 13530 899
rect 13478 856 13487 890
rect 13487 856 13521 890
rect 13521 856 13530 890
rect 13478 847 13530 856
rect 13682 890 13734 899
rect 13682 856 13691 890
rect 13691 856 13725 890
rect 13725 856 13734 890
rect 13682 847 13734 856
rect 13886 890 13938 899
rect 13886 856 13895 890
rect 13895 856 13929 890
rect 13929 856 13938 890
rect 13886 847 13938 856
rect 14090 890 14142 899
rect 14090 856 14099 890
rect 14099 856 14133 890
rect 14133 856 14142 890
rect 14090 847 14142 856
rect 14294 890 14346 899
rect 14294 856 14303 890
rect 14303 856 14337 890
rect 14337 856 14346 890
rect 14294 847 14346 856
rect 14498 890 14550 899
rect 14498 856 14507 890
rect 14507 856 14541 890
rect 14541 856 14550 890
rect 14498 847 14550 856
rect 14702 890 14754 899
rect 14702 856 14711 890
rect 14711 856 14745 890
rect 14745 856 14754 890
rect 14702 847 14754 856
rect 14906 890 14958 899
rect 14906 856 14915 890
rect 14915 856 14949 890
rect 14949 856 14958 890
rect 14906 847 14958 856
rect 15110 890 15162 899
rect 15110 856 15119 890
rect 15119 856 15153 890
rect 15153 856 15162 890
rect 15110 847 15162 856
rect 15314 890 15366 899
rect 15314 856 15323 890
rect 15323 856 15357 890
rect 15357 856 15366 890
rect 15314 847 15366 856
rect 15518 890 15570 899
rect 15518 856 15527 890
rect 15527 856 15561 890
rect 15561 856 15570 890
rect 15518 847 15570 856
rect 15722 890 15774 899
rect 15722 856 15731 890
rect 15731 856 15765 890
rect 15765 856 15774 890
rect 15722 847 15774 856
rect 15926 890 15978 899
rect 15926 856 15935 890
rect 15935 856 15969 890
rect 15969 856 15978 890
rect 15926 847 15978 856
rect 16130 890 16182 899
rect 16130 856 16139 890
rect 16139 856 16173 890
rect 16173 856 16182 890
rect 16130 847 16182 856
rect 16334 890 16386 899
rect 16334 856 16343 890
rect 16343 856 16377 890
rect 16377 856 16386 890
rect 16334 847 16386 856
rect 16538 890 16590 899
rect 16538 856 16547 890
rect 16547 856 16581 890
rect 16581 856 16590 890
rect 16538 847 16590 856
rect 16742 890 16794 899
rect 16742 856 16751 890
rect 16751 856 16785 890
rect 16785 856 16794 890
rect 16742 847 16794 856
rect 16946 890 16998 899
rect 16946 856 16955 890
rect 16955 856 16989 890
rect 16989 856 16998 890
rect 16946 847 16998 856
rect 17150 890 17202 899
rect 17150 856 17159 890
rect 17159 856 17193 890
rect 17193 856 17202 890
rect 17150 847 17202 856
rect 17354 890 17406 899
rect 17354 856 17363 890
rect 17363 856 17397 890
rect 17397 856 17406 890
rect 17354 847 17406 856
rect 17558 890 17610 899
rect 17558 856 17567 890
rect 17567 856 17601 890
rect 17601 856 17610 890
rect 17558 847 17610 856
rect 17762 890 17814 899
rect 17762 856 17771 890
rect 17771 856 17805 890
rect 17805 856 17814 890
rect 17762 847 17814 856
rect 17966 890 18018 899
rect 17966 856 17975 890
rect 17975 856 18009 890
rect 18009 856 18018 890
rect 17966 847 18018 856
rect 18170 890 18222 899
rect 18170 856 18179 890
rect 18179 856 18213 890
rect 18213 856 18222 890
rect 18170 847 18222 856
rect 18374 890 18426 899
rect 18374 856 18383 890
rect 18383 856 18417 890
rect 18417 856 18426 890
rect 18374 847 18426 856
rect 18578 890 18630 899
rect 18578 856 18587 890
rect 18587 856 18621 890
rect 18621 856 18630 890
rect 18578 847 18630 856
rect 18782 890 18834 899
rect 18782 856 18791 890
rect 18791 856 18825 890
rect 18825 856 18834 890
rect 18782 847 18834 856
rect 18986 890 19038 899
rect 18986 856 18995 890
rect 18995 856 19029 890
rect 19029 856 19038 890
rect 18986 847 19038 856
rect 19190 890 19242 899
rect 19190 856 19199 890
rect 19199 856 19233 890
rect 19233 856 19242 890
rect 19190 847 19242 856
rect 19394 890 19446 899
rect 19394 856 19403 890
rect 19403 856 19437 890
rect 19437 856 19446 890
rect 19394 847 19446 856
rect 19598 890 19650 899
rect 19598 856 19607 890
rect 19607 856 19641 890
rect 19641 856 19650 890
rect 19598 847 19650 856
rect 19802 890 19854 899
rect 19802 856 19811 890
rect 19811 856 19845 890
rect 19845 856 19854 890
rect 19802 847 19854 856
rect 20006 890 20058 899
rect 20006 856 20015 890
rect 20015 856 20049 890
rect 20049 856 20058 890
rect 20006 847 20058 856
rect 20210 890 20262 899
rect 20210 856 20219 890
rect 20219 856 20253 890
rect 20253 856 20262 890
rect 20210 847 20262 856
rect 20414 890 20466 899
rect 20414 856 20423 890
rect 20423 856 20457 890
rect 20457 856 20466 890
rect 20414 847 20466 856
rect 20618 890 20670 899
rect 20618 856 20627 890
rect 20627 856 20661 890
rect 20661 856 20670 890
rect 20618 847 20670 856
rect 20822 890 20874 899
rect 20822 856 20831 890
rect 20831 856 20865 890
rect 20865 856 20874 890
rect 20822 847 20874 856
rect 21026 890 21078 899
rect 21026 856 21035 890
rect 21035 856 21069 890
rect 21069 856 21078 890
rect 21026 847 21078 856
rect 21230 890 21282 899
rect 21230 856 21239 890
rect 21239 856 21273 890
rect 21273 856 21282 890
rect 21230 847 21282 856
rect 21434 890 21486 899
rect 21434 856 21443 890
rect 21443 856 21477 890
rect 21477 856 21486 890
rect 21434 847 21486 856
rect 21638 890 21690 899
rect 21638 856 21647 890
rect 21647 856 21681 890
rect 21681 856 21690 890
rect 21638 847 21690 856
rect 21842 890 21894 899
rect 21842 856 21851 890
rect 21851 856 21885 890
rect 21885 856 21894 890
rect 21842 847 21894 856
rect 22046 890 22098 899
rect 22046 856 22055 890
rect 22055 856 22089 890
rect 22089 856 22098 890
rect 22046 847 22098 856
rect 22250 890 22302 899
rect 22250 856 22259 890
rect 22259 856 22293 890
rect 22293 856 22302 890
rect 22250 847 22302 856
rect 22454 890 22506 899
rect 22454 856 22463 890
rect 22463 856 22497 890
rect 22497 856 22506 890
rect 22454 847 22506 856
rect 22658 890 22710 899
rect 22658 856 22667 890
rect 22667 856 22701 890
rect 22701 856 22710 890
rect 22658 847 22710 856
rect 22862 890 22914 899
rect 22862 856 22871 890
rect 22871 856 22905 890
rect 22905 856 22914 890
rect 22862 847 22914 856
rect 23066 890 23118 899
rect 23066 856 23075 890
rect 23075 856 23109 890
rect 23109 856 23118 890
rect 23066 847 23118 856
rect 23270 890 23322 899
rect 23270 856 23279 890
rect 23279 856 23313 890
rect 23313 856 23322 890
rect 23270 847 23322 856
rect 23474 890 23526 899
rect 23474 856 23483 890
rect 23483 856 23517 890
rect 23517 856 23526 890
rect 23474 847 23526 856
rect 23678 890 23730 899
rect 23678 856 23687 890
rect 23687 856 23721 890
rect 23721 856 23730 890
rect 23678 847 23730 856
rect 23882 890 23934 899
rect 23882 856 23891 890
rect 23891 856 23925 890
rect 23925 856 23934 890
rect 23882 847 23934 856
rect 24086 890 24138 899
rect 24086 856 24095 890
rect 24095 856 24129 890
rect 24129 856 24138 890
rect 24086 847 24138 856
rect 24290 890 24342 899
rect 24290 856 24299 890
rect 24299 856 24333 890
rect 24333 856 24342 890
rect 24290 847 24342 856
rect 24494 890 24546 899
rect 24494 856 24503 890
rect 24503 856 24537 890
rect 24537 856 24546 890
rect 24494 847 24546 856
rect 24698 890 24750 899
rect 24698 856 24707 890
rect 24707 856 24741 890
rect 24741 856 24750 890
rect 24698 847 24750 856
rect 24902 890 24954 899
rect 24902 856 24911 890
rect 24911 856 24945 890
rect 24945 856 24954 890
rect 24902 847 24954 856
rect 25106 890 25158 899
rect 25106 856 25115 890
rect 25115 856 25149 890
rect 25149 856 25158 890
rect 25106 847 25158 856
rect 25310 890 25362 899
rect 25310 856 25319 890
rect 25319 856 25353 890
rect 25353 856 25362 890
rect 25310 847 25362 856
rect 25514 890 25566 899
rect 25514 856 25523 890
rect 25523 856 25557 890
rect 25557 856 25566 890
rect 25514 847 25566 856
rect 25718 890 25770 899
rect 25718 856 25727 890
rect 25727 856 25761 890
rect 25761 856 25770 890
rect 25718 847 25770 856
rect 25922 890 25974 899
rect 25922 856 25931 890
rect 25931 856 25965 890
rect 25965 856 25974 890
rect 25922 847 25974 856
rect 26126 890 26178 899
rect 26126 856 26135 890
rect 26135 856 26169 890
rect 26169 856 26178 890
rect 26126 847 26178 856
rect 26330 890 26382 899
rect 26330 856 26339 890
rect 26339 856 26373 890
rect 26373 856 26382 890
rect 26330 847 26382 856
rect 26534 890 26586 899
rect 26534 856 26543 890
rect 26543 856 26577 890
rect 26577 856 26586 890
rect 26534 847 26586 856
rect 26738 890 26790 899
rect 26738 856 26747 890
rect 26747 856 26781 890
rect 26781 856 26790 890
rect 26738 847 26790 856
rect 26942 890 26994 899
rect 26942 856 26951 890
rect 26951 856 26985 890
rect 26985 856 26994 890
rect 26942 847 26994 856
rect 27146 890 27198 899
rect 27146 856 27155 890
rect 27155 856 27189 890
rect 27189 856 27198 890
rect 27146 847 27198 856
rect 27350 890 27402 899
rect 27350 856 27359 890
rect 27359 856 27393 890
rect 27393 856 27402 890
rect 27350 847 27402 856
rect 27554 890 27606 899
rect 27554 856 27563 890
rect 27563 856 27597 890
rect 27597 856 27606 890
rect 27554 847 27606 856
rect 27758 890 27810 899
rect 27758 856 27767 890
rect 27767 856 27801 890
rect 27801 856 27810 890
rect 27758 847 27810 856
rect 27962 890 28014 899
rect 27962 856 27971 890
rect 27971 856 28005 890
rect 28005 856 28014 890
rect 27962 847 28014 856
rect 28166 890 28218 899
rect 28166 856 28175 890
rect 28175 856 28209 890
rect 28209 856 28218 890
rect 28166 847 28218 856
rect 28370 890 28422 899
rect 28370 856 28379 890
rect 28379 856 28413 890
rect 28413 856 28422 890
rect 28370 847 28422 856
rect 28574 890 28626 899
rect 28574 856 28583 890
rect 28583 856 28617 890
rect 28617 856 28626 890
rect 28574 847 28626 856
rect 28778 890 28830 899
rect 28778 856 28787 890
rect 28787 856 28821 890
rect 28821 856 28830 890
rect 28778 847 28830 856
rect 28982 890 29034 899
rect 28982 856 28991 890
rect 28991 856 29025 890
rect 29025 856 29034 890
rect 28982 847 29034 856
rect 29186 890 29238 899
rect 29186 856 29195 890
rect 29195 856 29229 890
rect 29229 856 29238 890
rect 29186 847 29238 856
rect 29390 890 29442 899
rect 29390 856 29399 890
rect 29399 856 29433 890
rect 29433 856 29442 890
rect 29390 847 29442 856
rect 29594 890 29646 899
rect 29594 856 29603 890
rect 29603 856 29637 890
rect 29637 856 29646 890
rect 29594 847 29646 856
rect 29798 890 29850 899
rect 29798 856 29807 890
rect 29807 856 29841 890
rect 29841 856 29850 890
rect 29798 847 29850 856
rect 30002 890 30054 899
rect 30002 856 30011 890
rect 30011 856 30045 890
rect 30045 856 30054 890
rect 30002 847 30054 856
rect 30206 890 30258 899
rect 30206 856 30215 890
rect 30215 856 30249 890
rect 30249 856 30258 890
rect 30206 847 30258 856
rect 30410 890 30462 899
rect 30410 856 30419 890
rect 30419 856 30453 890
rect 30453 856 30462 890
rect 30410 847 30462 856
rect 30614 890 30666 899
rect 30614 856 30623 890
rect 30623 856 30657 890
rect 30657 856 30666 890
rect 30614 847 30666 856
rect 30818 890 30870 899
rect 30818 856 30827 890
rect 30827 856 30861 890
rect 30861 856 30870 890
rect 30818 847 30870 856
rect 31022 890 31074 899
rect 31022 856 31031 890
rect 31031 856 31065 890
rect 31065 856 31074 890
rect 31022 847 31074 856
rect 31226 890 31278 899
rect 31226 856 31235 890
rect 31235 856 31269 890
rect 31269 856 31278 890
rect 31226 847 31278 856
rect 31430 890 31482 899
rect 31430 856 31439 890
rect 31439 856 31473 890
rect 31473 856 31482 890
rect 31430 847 31482 856
rect 31634 890 31686 899
rect 31634 856 31643 890
rect 31643 856 31677 890
rect 31677 856 31686 890
rect 31634 847 31686 856
rect 31838 890 31890 899
rect 31838 856 31847 890
rect 31847 856 31881 890
rect 31881 856 31890 890
rect 31838 847 31890 856
rect 32042 890 32094 899
rect 32042 856 32051 890
rect 32051 856 32085 890
rect 32085 856 32094 890
rect 32042 847 32094 856
rect 32246 890 32298 899
rect 32246 856 32255 890
rect 32255 856 32289 890
rect 32289 856 32298 890
rect 32246 847 32298 856
rect 32450 890 32502 899
rect 32450 856 32459 890
rect 32459 856 32493 890
rect 32493 856 32502 890
rect 32450 847 32502 856
rect 32654 890 32706 899
rect 32654 856 32663 890
rect 32663 856 32697 890
rect 32697 856 32706 890
rect 32654 847 32706 856
rect 32858 890 32910 899
rect 32858 856 32867 890
rect 32867 856 32901 890
rect 32901 856 32910 890
rect 32858 847 32910 856
rect 33062 890 33114 899
rect 33062 856 33071 890
rect 33071 856 33105 890
rect 33105 856 33114 890
rect 33062 847 33114 856
rect 33266 890 33318 899
rect 33266 856 33275 890
rect 33275 856 33309 890
rect 33309 856 33318 890
rect 33266 847 33318 856
rect 33470 890 33522 899
rect 33470 856 33479 890
rect 33479 856 33513 890
rect 33513 856 33522 890
rect 33470 847 33522 856
rect 33674 890 33726 899
rect 33674 856 33683 890
rect 33683 856 33717 890
rect 33717 856 33726 890
rect 33674 847 33726 856
rect 33878 890 33930 899
rect 33878 856 33887 890
rect 33887 856 33921 890
rect 33921 856 33930 890
rect 33878 847 33930 856
rect 34082 890 34134 899
rect 34082 856 34091 890
rect 34091 856 34125 890
rect 34125 856 34134 890
rect 34082 847 34134 856
rect 34286 890 34338 899
rect 34286 856 34295 890
rect 34295 856 34329 890
rect 34329 856 34338 890
rect 34286 847 34338 856
rect 34490 890 34542 899
rect 34490 856 34499 890
rect 34499 856 34533 890
rect 34533 856 34542 890
rect 34490 847 34542 856
rect 34694 890 34746 899
rect 34694 856 34703 890
rect 34703 856 34737 890
rect 34737 856 34746 890
rect 34694 847 34746 856
rect 34898 890 34950 899
rect 34898 856 34907 890
rect 34907 856 34941 890
rect 34941 856 34950 890
rect 34898 847 34950 856
rect 35102 890 35154 899
rect 35102 856 35111 890
rect 35111 856 35145 890
rect 35145 856 35154 890
rect 35102 847 35154 856
rect 35306 890 35358 899
rect 35306 856 35315 890
rect 35315 856 35349 890
rect 35349 856 35358 890
rect 35306 847 35358 856
rect 35510 890 35562 899
rect 35510 856 35519 890
rect 35519 856 35553 890
rect 35553 856 35562 890
rect 35510 847 35562 856
rect 35714 890 35766 899
rect 35714 856 35723 890
rect 35723 856 35757 890
rect 35757 856 35766 890
rect 35714 847 35766 856
rect 35918 890 35970 899
rect 35918 856 35927 890
rect 35927 856 35961 890
rect 35961 856 35970 890
rect 35918 847 35970 856
rect 36122 890 36174 899
rect 36122 856 36131 890
rect 36131 856 36165 890
rect 36165 856 36174 890
rect 36122 847 36174 856
rect 36326 890 36378 899
rect 36326 856 36335 890
rect 36335 856 36369 890
rect 36369 856 36378 890
rect 36326 847 36378 856
rect 36530 890 36582 899
rect 36530 856 36539 890
rect 36539 856 36573 890
rect 36573 856 36582 890
rect 36530 847 36582 856
rect 36734 890 36786 899
rect 36734 856 36743 890
rect 36743 856 36777 890
rect 36777 856 36786 890
rect 36734 847 36786 856
rect 36938 890 36990 899
rect 36938 856 36947 890
rect 36947 856 36981 890
rect 36981 856 36990 890
rect 36938 847 36990 856
rect 37142 890 37194 899
rect 37142 856 37151 890
rect 37151 856 37185 890
rect 37185 856 37194 890
rect 37142 847 37194 856
rect 37346 890 37398 899
rect 37346 856 37355 890
rect 37355 856 37389 890
rect 37389 856 37398 890
rect 37346 847 37398 856
rect 37550 890 37602 899
rect 37550 856 37559 890
rect 37559 856 37593 890
rect 37593 856 37602 890
rect 37550 847 37602 856
rect 37754 890 37806 899
rect 37754 856 37763 890
rect 37763 856 37797 890
rect 37797 856 37806 890
rect 37754 847 37806 856
rect 37958 890 38010 899
rect 37958 856 37967 890
rect 37967 856 38001 890
rect 38001 856 38010 890
rect 37958 847 38010 856
rect 38162 890 38214 899
rect 38162 856 38171 890
rect 38171 856 38205 890
rect 38205 856 38214 890
rect 38162 847 38214 856
rect 38366 890 38418 899
rect 38366 856 38375 890
rect 38375 856 38409 890
rect 38409 856 38418 890
rect 38366 847 38418 856
rect 38570 890 38622 899
rect 38570 856 38579 890
rect 38579 856 38613 890
rect 38613 856 38622 890
rect 38570 847 38622 856
rect 38774 890 38826 899
rect 38774 856 38783 890
rect 38783 856 38817 890
rect 38817 856 38826 890
rect 38774 847 38826 856
rect 38978 890 39030 899
rect 38978 856 38987 890
rect 38987 856 39021 890
rect 39021 856 39030 890
rect 38978 847 39030 856
rect 39182 890 39234 899
rect 39182 856 39191 890
rect 39191 856 39225 890
rect 39225 856 39234 890
rect 39182 847 39234 856
rect 39386 890 39438 899
rect 39386 856 39395 890
rect 39395 856 39429 890
rect 39429 856 39438 890
rect 39386 847 39438 856
rect 39590 890 39642 899
rect 39590 856 39599 890
rect 39599 856 39633 890
rect 39633 856 39642 890
rect 39590 847 39642 856
rect 39794 890 39846 899
rect 39794 856 39803 890
rect 39803 856 39837 890
rect 39837 856 39846 890
rect 39794 847 39846 856
rect 39998 890 40050 899
rect 39998 856 40007 890
rect 40007 856 40041 890
rect 40041 856 40050 890
rect 39998 847 40050 856
rect 40202 890 40254 899
rect 40202 856 40211 890
rect 40211 856 40245 890
rect 40245 856 40254 890
rect 40202 847 40254 856
rect 40406 890 40458 899
rect 40406 856 40415 890
rect 40415 856 40449 890
rect 40449 856 40458 890
rect 40406 847 40458 856
rect 40610 890 40662 899
rect 40610 856 40619 890
rect 40619 856 40653 890
rect 40653 856 40662 890
rect 40610 847 40662 856
rect 40814 890 40866 899
rect 40814 856 40823 890
rect 40823 856 40857 890
rect 40857 856 40866 890
rect 40814 847 40866 856
rect 41018 890 41070 899
rect 41018 856 41027 890
rect 41027 856 41061 890
rect 41061 856 41070 890
rect 41018 847 41070 856
rect 41222 890 41274 899
rect 41222 856 41231 890
rect 41231 856 41265 890
rect 41265 856 41274 890
rect 41222 847 41274 856
rect 41426 890 41478 899
rect 41426 856 41435 890
rect 41435 856 41469 890
rect 41469 856 41478 890
rect 41426 847 41478 856
rect 41630 890 41682 899
rect 41630 856 41639 890
rect 41639 856 41673 890
rect 41673 856 41682 890
rect 41630 847 41682 856
rect 41834 890 41886 899
rect 41834 856 41843 890
rect 41843 856 41877 890
rect 41877 856 41886 890
rect 41834 847 41886 856
rect 42038 890 42090 899
rect 42038 856 42047 890
rect 42047 856 42081 890
rect 42081 856 42090 890
rect 42038 847 42090 856
rect 42242 890 42294 899
rect 42242 856 42251 890
rect 42251 856 42285 890
rect 42285 856 42294 890
rect 42242 847 42294 856
rect 42446 890 42498 899
rect 42446 856 42455 890
rect 42455 856 42489 890
rect 42489 856 42498 890
rect 42446 847 42498 856
rect 42650 890 42702 899
rect 42650 856 42659 890
rect 42659 856 42693 890
rect 42693 856 42702 890
rect 42650 847 42702 856
rect 42854 890 42906 899
rect 42854 856 42863 890
rect 42863 856 42897 890
rect 42897 856 42906 890
rect 42854 847 42906 856
rect 43058 890 43110 899
rect 43058 856 43067 890
rect 43067 856 43101 890
rect 43101 856 43110 890
rect 43058 847 43110 856
rect 43262 890 43314 899
rect 43262 856 43271 890
rect 43271 856 43305 890
rect 43305 856 43314 890
rect 43262 847 43314 856
rect 43466 890 43518 899
rect 43466 856 43475 890
rect 43475 856 43509 890
rect 43509 856 43518 890
rect 43466 847 43518 856
rect 43670 890 43722 899
rect 43670 856 43679 890
rect 43679 856 43713 890
rect 43713 856 43722 890
rect 43670 847 43722 856
rect 43874 890 43926 899
rect 43874 856 43883 890
rect 43883 856 43917 890
rect 43917 856 43926 890
rect 43874 847 43926 856
rect 44078 890 44130 899
rect 44078 856 44087 890
rect 44087 856 44121 890
rect 44121 856 44130 890
rect 44078 847 44130 856
rect 44282 890 44334 899
rect 44282 856 44291 890
rect 44291 856 44325 890
rect 44325 856 44334 890
rect 44282 847 44334 856
rect 44486 890 44538 899
rect 44486 856 44495 890
rect 44495 856 44529 890
rect 44529 856 44538 890
rect 44486 847 44538 856
rect 44690 890 44742 899
rect 44690 856 44699 890
rect 44699 856 44733 890
rect 44733 856 44742 890
rect 44690 847 44742 856
rect 44894 890 44946 899
rect 44894 856 44903 890
rect 44903 856 44937 890
rect 44937 856 44946 890
rect 44894 847 44946 856
rect 45098 890 45150 899
rect 45098 856 45107 890
rect 45107 856 45141 890
rect 45141 856 45150 890
rect 45098 847 45150 856
rect 45302 890 45354 899
rect 45302 856 45311 890
rect 45311 856 45345 890
rect 45345 856 45354 890
rect 45302 847 45354 856
rect 45506 890 45558 899
rect 45506 856 45515 890
rect 45515 856 45549 890
rect 45549 856 45558 890
rect 45506 847 45558 856
rect 45710 890 45762 899
rect 45710 856 45719 890
rect 45719 856 45753 890
rect 45753 856 45762 890
rect 45710 847 45762 856
rect 45914 890 45966 899
rect 45914 856 45923 890
rect 45923 856 45957 890
rect 45957 856 45966 890
rect 45914 847 45966 856
rect 46118 890 46170 899
rect 46118 856 46127 890
rect 46127 856 46161 890
rect 46161 856 46170 890
rect 46118 847 46170 856
rect 46322 890 46374 899
rect 46322 856 46331 890
rect 46331 856 46365 890
rect 46365 856 46374 890
rect 46322 847 46374 856
rect 46526 890 46578 899
rect 46526 856 46535 890
rect 46535 856 46569 890
rect 46569 856 46578 890
rect 46526 847 46578 856
rect 46730 890 46782 899
rect 46730 856 46739 890
rect 46739 856 46773 890
rect 46773 856 46782 890
rect 46730 847 46782 856
rect 46934 890 46986 899
rect 46934 856 46943 890
rect 46943 856 46977 890
rect 46977 856 46986 890
rect 46934 847 46986 856
rect 47138 890 47190 899
rect 47138 856 47147 890
rect 47147 856 47181 890
rect 47181 856 47190 890
rect 47138 847 47190 856
rect 47342 890 47394 899
rect 47342 856 47351 890
rect 47351 856 47385 890
rect 47385 856 47394 890
rect 47342 847 47394 856
rect 47546 890 47598 899
rect 47546 856 47555 890
rect 47555 856 47589 890
rect 47589 856 47598 890
rect 47546 847 47598 856
rect 47750 890 47802 899
rect 47750 856 47759 890
rect 47759 856 47793 890
rect 47793 856 47802 890
rect 47750 847 47802 856
rect 47954 890 48006 899
rect 47954 856 47963 890
rect 47963 856 47997 890
rect 47997 856 48006 890
rect 47954 847 48006 856
rect 48158 890 48210 899
rect 48158 856 48167 890
rect 48167 856 48201 890
rect 48201 856 48210 890
rect 48158 847 48210 856
rect 48362 890 48414 899
rect 48362 856 48371 890
rect 48371 856 48405 890
rect 48405 856 48414 890
rect 48362 847 48414 856
rect 48566 890 48618 899
rect 48566 856 48575 890
rect 48575 856 48609 890
rect 48609 856 48618 890
rect 48566 847 48618 856
rect 48770 890 48822 899
rect 48770 856 48779 890
rect 48779 856 48813 890
rect 48813 856 48822 890
rect 48770 847 48822 856
rect 48974 890 49026 899
rect 48974 856 48983 890
rect 48983 856 49017 890
rect 49017 856 49026 890
rect 48974 847 49026 856
rect 49178 890 49230 899
rect 49178 856 49187 890
rect 49187 856 49221 890
rect 49221 856 49230 890
rect 49178 847 49230 856
rect 49382 890 49434 899
rect 49382 856 49391 890
rect 49391 856 49425 890
rect 49425 856 49434 890
rect 49382 847 49434 856
rect 49586 890 49638 899
rect 49586 856 49595 890
rect 49595 856 49629 890
rect 49629 856 49638 890
rect 49586 847 49638 856
rect 49790 890 49842 899
rect 49790 856 49799 890
rect 49799 856 49833 890
rect 49833 856 49842 890
rect 49790 847 49842 856
rect 49994 890 50046 899
rect 49994 856 50003 890
rect 50003 856 50037 890
rect 50037 856 50046 890
rect 49994 847 50046 856
rect 50198 890 50250 899
rect 50198 856 50207 890
rect 50207 856 50241 890
rect 50241 856 50250 890
rect 50198 847 50250 856
rect 50402 890 50454 899
rect 50402 856 50411 890
rect 50411 856 50445 890
rect 50445 856 50454 890
rect 50402 847 50454 856
rect 50606 890 50658 899
rect 50606 856 50615 890
rect 50615 856 50649 890
rect 50649 856 50658 890
rect 50606 847 50658 856
rect 50810 890 50862 899
rect 50810 856 50819 890
rect 50819 856 50853 890
rect 50853 856 50862 890
rect 50810 847 50862 856
rect 51014 890 51066 899
rect 51014 856 51023 890
rect 51023 856 51057 890
rect 51057 856 51066 890
rect 51014 847 51066 856
rect 51218 890 51270 899
rect 51218 856 51227 890
rect 51227 856 51261 890
rect 51261 856 51270 890
rect 51218 847 51270 856
rect 51422 890 51474 899
rect 51422 856 51431 890
rect 51431 856 51465 890
rect 51465 856 51474 890
rect 51422 847 51474 856
rect 51626 890 51678 899
rect 51626 856 51635 890
rect 51635 856 51669 890
rect 51669 856 51678 890
rect 51626 847 51678 856
rect 51830 890 51882 899
rect 51830 856 51839 890
rect 51839 856 51873 890
rect 51873 856 51882 890
rect 51830 847 51882 856
rect 52034 890 52086 899
rect 52034 856 52043 890
rect 52043 856 52077 890
rect 52077 856 52086 890
rect 52034 847 52086 856
rect 52252 890 52304 899
rect 52252 856 52261 890
rect 52261 856 52295 890
rect 52295 856 52304 890
rect 52252 847 52304 856
<< metal2 >>
rect 7 2685 59 2691
rect 1 2638 7 2681
rect 1639 2685 1691 2691
rect 59 2673 65 2681
rect 1633 2673 1639 2681
rect 59 2645 1639 2673
rect 59 2638 65 2645
rect 1633 2638 1639 2645
rect 7 2627 59 2633
rect 3271 2685 3323 2691
rect 1691 2673 1697 2681
rect 3265 2673 3271 2681
rect 1691 2645 3271 2673
rect 1691 2638 1697 2645
rect 3265 2638 3271 2645
rect 1639 2627 1691 2633
rect 4903 2685 4955 2691
rect 3323 2673 3329 2681
rect 4897 2673 4903 2681
rect 3323 2645 4903 2673
rect 3323 2638 3329 2645
rect 4897 2638 4903 2645
rect 3271 2627 3323 2633
rect 6535 2685 6587 2691
rect 4955 2673 4961 2681
rect 6529 2673 6535 2681
rect 4955 2645 6535 2673
rect 4955 2638 4961 2645
rect 6529 2638 6535 2645
rect 4903 2627 4955 2633
rect 8167 2685 8219 2691
rect 6587 2673 6593 2681
rect 8161 2673 8167 2681
rect 6587 2645 8167 2673
rect 6587 2638 6593 2645
rect 8161 2638 8167 2645
rect 6535 2627 6587 2633
rect 9799 2685 9851 2691
rect 8219 2673 8225 2681
rect 9793 2673 9799 2681
rect 8219 2645 9799 2673
rect 8219 2638 8225 2645
rect 9793 2638 9799 2645
rect 8167 2627 8219 2633
rect 11431 2685 11483 2691
rect 9851 2673 9857 2681
rect 11425 2673 11431 2681
rect 9851 2645 11431 2673
rect 9851 2638 9857 2645
rect 11425 2638 11431 2645
rect 9799 2627 9851 2633
rect 13063 2685 13115 2691
rect 11483 2673 11489 2681
rect 13057 2673 13063 2681
rect 11483 2645 13063 2673
rect 11483 2638 11489 2645
rect 13057 2638 13063 2645
rect 11431 2627 11483 2633
rect 14695 2685 14747 2691
rect 13115 2673 13121 2681
rect 14689 2673 14695 2681
rect 13115 2645 14695 2673
rect 13115 2638 13121 2645
rect 14689 2638 14695 2645
rect 13063 2627 13115 2633
rect 16327 2685 16379 2691
rect 14747 2673 14753 2681
rect 16321 2673 16327 2681
rect 14747 2645 16327 2673
rect 14747 2638 14753 2645
rect 16321 2638 16327 2645
rect 14695 2627 14747 2633
rect 17959 2685 18011 2691
rect 16379 2673 16385 2681
rect 17953 2673 17959 2681
rect 16379 2645 17959 2673
rect 16379 2638 16385 2645
rect 17953 2638 17959 2645
rect 16327 2627 16379 2633
rect 19591 2685 19643 2691
rect 18011 2673 18017 2681
rect 19585 2673 19591 2681
rect 18011 2645 19591 2673
rect 18011 2638 18017 2645
rect 19585 2638 19591 2645
rect 17959 2627 18011 2633
rect 21223 2685 21275 2691
rect 19643 2673 19649 2681
rect 21217 2673 21223 2681
rect 19643 2645 21223 2673
rect 19643 2638 19649 2645
rect 21217 2638 21223 2645
rect 19591 2627 19643 2633
rect 22855 2685 22907 2691
rect 21275 2673 21281 2681
rect 22849 2673 22855 2681
rect 21275 2645 22855 2673
rect 21275 2638 21281 2645
rect 22849 2638 22855 2645
rect 21223 2627 21275 2633
rect 24487 2685 24539 2691
rect 22907 2673 22913 2681
rect 24481 2673 24487 2681
rect 22907 2645 24487 2673
rect 22907 2638 22913 2645
rect 24481 2638 24487 2645
rect 22855 2627 22907 2633
rect 26119 2685 26171 2691
rect 24539 2673 24545 2681
rect 26113 2673 26119 2681
rect 24539 2645 26119 2673
rect 24539 2638 24545 2645
rect 26113 2638 26119 2645
rect 24487 2627 24539 2633
rect 27751 2685 27803 2691
rect 26171 2673 26177 2681
rect 27745 2673 27751 2681
rect 26171 2645 27751 2673
rect 26171 2638 26177 2645
rect 27745 2638 27751 2645
rect 26119 2627 26171 2633
rect 29383 2685 29435 2691
rect 27803 2673 27809 2681
rect 29377 2673 29383 2681
rect 27803 2645 29383 2673
rect 27803 2638 27809 2645
rect 29377 2638 29383 2645
rect 27751 2627 27803 2633
rect 31015 2685 31067 2691
rect 29435 2673 29441 2681
rect 31009 2673 31015 2681
rect 29435 2645 31015 2673
rect 29435 2638 29441 2645
rect 31009 2638 31015 2645
rect 29383 2627 29435 2633
rect 32647 2685 32699 2691
rect 31067 2673 31073 2681
rect 32641 2673 32647 2681
rect 31067 2645 32647 2673
rect 31067 2638 31073 2645
rect 32641 2638 32647 2645
rect 31015 2627 31067 2633
rect 34279 2685 34331 2691
rect 32699 2673 32705 2681
rect 34273 2673 34279 2681
rect 32699 2645 34279 2673
rect 32699 2638 32705 2645
rect 34273 2638 34279 2645
rect 32647 2627 32699 2633
rect 35911 2685 35963 2691
rect 34331 2673 34337 2681
rect 35905 2673 35911 2681
rect 34331 2645 35911 2673
rect 34331 2638 34337 2645
rect 35905 2638 35911 2645
rect 34279 2627 34331 2633
rect 37543 2685 37595 2691
rect 35963 2673 35969 2681
rect 37537 2673 37543 2681
rect 35963 2645 37543 2673
rect 35963 2638 35969 2645
rect 37537 2638 37543 2645
rect 35911 2627 35963 2633
rect 39175 2685 39227 2691
rect 37595 2673 37601 2681
rect 39169 2673 39175 2681
rect 37595 2645 39175 2673
rect 37595 2638 37601 2645
rect 39169 2638 39175 2645
rect 37543 2627 37595 2633
rect 40807 2685 40859 2691
rect 39227 2673 39233 2681
rect 40801 2673 40807 2681
rect 39227 2645 40807 2673
rect 39227 2638 39233 2645
rect 40801 2638 40807 2645
rect 39175 2627 39227 2633
rect 42439 2685 42491 2691
rect 40859 2673 40865 2681
rect 42433 2673 42439 2681
rect 40859 2645 42439 2673
rect 40859 2638 40865 2645
rect 42433 2638 42439 2645
rect 40807 2627 40859 2633
rect 44071 2685 44123 2691
rect 42491 2673 42497 2681
rect 44065 2673 44071 2681
rect 42491 2645 44071 2673
rect 42491 2638 42497 2645
rect 44065 2638 44071 2645
rect 42439 2627 42491 2633
rect 45703 2685 45755 2691
rect 44123 2673 44129 2681
rect 45697 2673 45703 2681
rect 44123 2645 45703 2673
rect 44123 2638 44129 2645
rect 45697 2638 45703 2645
rect 44071 2627 44123 2633
rect 47335 2685 47387 2691
rect 45755 2673 45761 2681
rect 47329 2673 47335 2681
rect 45755 2645 47335 2673
rect 45755 2638 45761 2645
rect 47329 2638 47335 2645
rect 45703 2627 45755 2633
rect 48967 2685 49019 2691
rect 47387 2673 47393 2681
rect 48961 2673 48967 2681
rect 47387 2645 48967 2673
rect 47387 2638 47393 2645
rect 48961 2638 48967 2645
rect 47335 2627 47387 2633
rect 50599 2685 50651 2691
rect 49019 2673 49025 2681
rect 50593 2673 50599 2681
rect 49019 2645 50599 2673
rect 49019 2638 49025 2645
rect 50593 2638 50599 2645
rect 48967 2627 49019 2633
rect 52231 2685 52283 2691
rect 50651 2673 50657 2681
rect 52225 2673 52231 2681
rect 50651 2645 52231 2673
rect 50651 2638 50657 2645
rect 52225 2638 52231 2645
rect 50599 2627 50651 2633
rect 52283 2638 52289 2681
rect 52231 2627 52283 2633
rect 7 2481 59 2487
rect 1 2434 7 2477
rect 1639 2481 1691 2487
rect 59 2469 65 2477
rect 1633 2469 1639 2477
rect 59 2441 1639 2469
rect 59 2434 65 2441
rect 1633 2434 1639 2441
rect 7 2423 59 2429
rect 3271 2481 3323 2487
rect 1691 2469 1697 2477
rect 3265 2469 3271 2477
rect 1691 2441 3271 2469
rect 1691 2434 1697 2441
rect 3265 2434 3271 2441
rect 1639 2423 1691 2429
rect 4903 2481 4955 2487
rect 3323 2469 3329 2477
rect 4897 2469 4903 2477
rect 3323 2441 4903 2469
rect 3323 2434 3329 2441
rect 4897 2434 4903 2441
rect 3271 2423 3323 2429
rect 6535 2481 6587 2487
rect 4955 2469 4961 2477
rect 6529 2469 6535 2477
rect 4955 2441 6535 2469
rect 4955 2434 4961 2441
rect 6529 2434 6535 2441
rect 4903 2423 4955 2429
rect 8167 2481 8219 2487
rect 6587 2469 6593 2477
rect 8161 2469 8167 2477
rect 6587 2441 8167 2469
rect 6587 2434 6593 2441
rect 8161 2434 8167 2441
rect 6535 2423 6587 2429
rect 9799 2481 9851 2487
rect 8219 2469 8225 2477
rect 9793 2469 9799 2477
rect 8219 2441 9799 2469
rect 8219 2434 8225 2441
rect 9793 2434 9799 2441
rect 8167 2423 8219 2429
rect 11431 2481 11483 2487
rect 9851 2469 9857 2477
rect 11425 2469 11431 2477
rect 9851 2441 11431 2469
rect 9851 2434 9857 2441
rect 11425 2434 11431 2441
rect 9799 2423 9851 2429
rect 13063 2481 13115 2487
rect 11483 2469 11489 2477
rect 13057 2469 13063 2477
rect 11483 2441 13063 2469
rect 11483 2434 11489 2441
rect 13057 2434 13063 2441
rect 11431 2423 11483 2429
rect 14695 2481 14747 2487
rect 13115 2469 13121 2477
rect 14689 2469 14695 2477
rect 13115 2441 14695 2469
rect 13115 2434 13121 2441
rect 14689 2434 14695 2441
rect 13063 2423 13115 2429
rect 16327 2481 16379 2487
rect 14747 2469 14753 2477
rect 16321 2469 16327 2477
rect 14747 2441 16327 2469
rect 14747 2434 14753 2441
rect 16321 2434 16327 2441
rect 14695 2423 14747 2429
rect 17959 2481 18011 2487
rect 16379 2469 16385 2477
rect 17953 2469 17959 2477
rect 16379 2441 17959 2469
rect 16379 2434 16385 2441
rect 17953 2434 17959 2441
rect 16327 2423 16379 2429
rect 19591 2481 19643 2487
rect 18011 2469 18017 2477
rect 19585 2469 19591 2477
rect 18011 2441 19591 2469
rect 18011 2434 18017 2441
rect 19585 2434 19591 2441
rect 17959 2423 18011 2429
rect 21223 2481 21275 2487
rect 19643 2469 19649 2477
rect 21217 2469 21223 2477
rect 19643 2441 21223 2469
rect 19643 2434 19649 2441
rect 21217 2434 21223 2441
rect 19591 2423 19643 2429
rect 22855 2481 22907 2487
rect 21275 2469 21281 2477
rect 22849 2469 22855 2477
rect 21275 2441 22855 2469
rect 21275 2434 21281 2441
rect 22849 2434 22855 2441
rect 21223 2423 21275 2429
rect 24487 2481 24539 2487
rect 22907 2469 22913 2477
rect 24481 2469 24487 2477
rect 22907 2441 24487 2469
rect 22907 2434 22913 2441
rect 24481 2434 24487 2441
rect 22855 2423 22907 2429
rect 26119 2481 26171 2487
rect 24539 2469 24545 2477
rect 26113 2469 26119 2477
rect 24539 2441 26119 2469
rect 24539 2434 24545 2441
rect 26113 2434 26119 2441
rect 24487 2423 24539 2429
rect 27751 2481 27803 2487
rect 26171 2469 26177 2477
rect 27745 2469 27751 2477
rect 26171 2441 27751 2469
rect 26171 2434 26177 2441
rect 27745 2434 27751 2441
rect 26119 2423 26171 2429
rect 29383 2481 29435 2487
rect 27803 2469 27809 2477
rect 29377 2469 29383 2477
rect 27803 2441 29383 2469
rect 27803 2434 27809 2441
rect 29377 2434 29383 2441
rect 27751 2423 27803 2429
rect 31015 2481 31067 2487
rect 29435 2469 29441 2477
rect 31009 2469 31015 2477
rect 29435 2441 31015 2469
rect 29435 2434 29441 2441
rect 31009 2434 31015 2441
rect 29383 2423 29435 2429
rect 32647 2481 32699 2487
rect 31067 2469 31073 2477
rect 32641 2469 32647 2477
rect 31067 2441 32647 2469
rect 31067 2434 31073 2441
rect 32641 2434 32647 2441
rect 31015 2423 31067 2429
rect 34279 2481 34331 2487
rect 32699 2469 32705 2477
rect 34273 2469 34279 2477
rect 32699 2441 34279 2469
rect 32699 2434 32705 2441
rect 34273 2434 34279 2441
rect 32647 2423 32699 2429
rect 35911 2481 35963 2487
rect 34331 2469 34337 2477
rect 35905 2469 35911 2477
rect 34331 2441 35911 2469
rect 34331 2434 34337 2441
rect 35905 2434 35911 2441
rect 34279 2423 34331 2429
rect 37543 2481 37595 2487
rect 35963 2469 35969 2477
rect 37537 2469 37543 2477
rect 35963 2441 37543 2469
rect 35963 2434 35969 2441
rect 37537 2434 37543 2441
rect 35911 2423 35963 2429
rect 39175 2481 39227 2487
rect 37595 2469 37601 2477
rect 39169 2469 39175 2477
rect 37595 2441 39175 2469
rect 37595 2434 37601 2441
rect 39169 2434 39175 2441
rect 37543 2423 37595 2429
rect 40807 2481 40859 2487
rect 39227 2469 39233 2477
rect 40801 2469 40807 2477
rect 39227 2441 40807 2469
rect 39227 2434 39233 2441
rect 40801 2434 40807 2441
rect 39175 2423 39227 2429
rect 42439 2481 42491 2487
rect 40859 2469 40865 2477
rect 42433 2469 42439 2477
rect 40859 2441 42439 2469
rect 40859 2434 40865 2441
rect 42433 2434 42439 2441
rect 40807 2423 40859 2429
rect 44071 2481 44123 2487
rect 42491 2469 42497 2477
rect 44065 2469 44071 2477
rect 42491 2441 44071 2469
rect 42491 2434 42497 2441
rect 44065 2434 44071 2441
rect 42439 2423 42491 2429
rect 45703 2481 45755 2487
rect 44123 2469 44129 2477
rect 45697 2469 45703 2477
rect 44123 2441 45703 2469
rect 44123 2434 44129 2441
rect 45697 2434 45703 2441
rect 44071 2423 44123 2429
rect 47335 2481 47387 2487
rect 45755 2469 45761 2477
rect 47329 2469 47335 2477
rect 45755 2441 47335 2469
rect 45755 2434 45761 2441
rect 47329 2434 47335 2441
rect 45703 2423 45755 2429
rect 48967 2481 49019 2487
rect 47387 2469 47393 2477
rect 48961 2469 48967 2477
rect 47387 2441 48967 2469
rect 47387 2434 47393 2441
rect 48961 2434 48967 2441
rect 47335 2423 47387 2429
rect 50599 2481 50651 2487
rect 49019 2469 49025 2477
rect 50593 2469 50599 2477
rect 49019 2441 50599 2469
rect 49019 2434 49025 2441
rect 50593 2434 50599 2441
rect 48967 2423 49019 2429
rect 52231 2481 52283 2487
rect 50651 2469 50657 2477
rect 52225 2469 52231 2477
rect 50651 2441 52231 2469
rect 50651 2434 50657 2441
rect 52225 2434 52231 2441
rect 50599 2423 50651 2429
rect 52283 2434 52289 2477
rect 52231 2423 52283 2429
rect 7 2277 59 2283
rect 1 2230 7 2273
rect 1639 2277 1691 2283
rect 59 2265 65 2273
rect 1633 2265 1639 2273
rect 59 2237 1639 2265
rect 59 2230 65 2237
rect 1633 2230 1639 2237
rect 7 2219 59 2225
rect 3271 2277 3323 2283
rect 1691 2265 1697 2273
rect 3265 2265 3271 2273
rect 1691 2237 3271 2265
rect 1691 2230 1697 2237
rect 3265 2230 3271 2237
rect 1639 2219 1691 2225
rect 4903 2277 4955 2283
rect 3323 2265 3329 2273
rect 4897 2265 4903 2273
rect 3323 2237 4903 2265
rect 3323 2230 3329 2237
rect 4897 2230 4903 2237
rect 3271 2219 3323 2225
rect 6535 2277 6587 2283
rect 4955 2265 4961 2273
rect 6529 2265 6535 2273
rect 4955 2237 6535 2265
rect 4955 2230 4961 2237
rect 6529 2230 6535 2237
rect 4903 2219 4955 2225
rect 8167 2277 8219 2283
rect 6587 2265 6593 2273
rect 8161 2265 8167 2273
rect 6587 2237 8167 2265
rect 6587 2230 6593 2237
rect 8161 2230 8167 2237
rect 6535 2219 6587 2225
rect 9799 2277 9851 2283
rect 8219 2265 8225 2273
rect 9793 2265 9799 2273
rect 8219 2237 9799 2265
rect 8219 2230 8225 2237
rect 9793 2230 9799 2237
rect 8167 2219 8219 2225
rect 11431 2277 11483 2283
rect 9851 2265 9857 2273
rect 11425 2265 11431 2273
rect 9851 2237 11431 2265
rect 9851 2230 9857 2237
rect 11425 2230 11431 2237
rect 9799 2219 9851 2225
rect 13063 2277 13115 2283
rect 11483 2265 11489 2273
rect 13057 2265 13063 2273
rect 11483 2237 13063 2265
rect 11483 2230 11489 2237
rect 13057 2230 13063 2237
rect 11431 2219 11483 2225
rect 14695 2277 14747 2283
rect 13115 2265 13121 2273
rect 14689 2265 14695 2273
rect 13115 2237 14695 2265
rect 13115 2230 13121 2237
rect 14689 2230 14695 2237
rect 13063 2219 13115 2225
rect 16327 2277 16379 2283
rect 14747 2265 14753 2273
rect 16321 2265 16327 2273
rect 14747 2237 16327 2265
rect 14747 2230 14753 2237
rect 16321 2230 16327 2237
rect 14695 2219 14747 2225
rect 17959 2277 18011 2283
rect 16379 2265 16385 2273
rect 17953 2265 17959 2273
rect 16379 2237 17959 2265
rect 16379 2230 16385 2237
rect 17953 2230 17959 2237
rect 16327 2219 16379 2225
rect 19591 2277 19643 2283
rect 18011 2265 18017 2273
rect 19585 2265 19591 2273
rect 18011 2237 19591 2265
rect 18011 2230 18017 2237
rect 19585 2230 19591 2237
rect 17959 2219 18011 2225
rect 21223 2277 21275 2283
rect 19643 2265 19649 2273
rect 21217 2265 21223 2273
rect 19643 2237 21223 2265
rect 19643 2230 19649 2237
rect 21217 2230 21223 2237
rect 19591 2219 19643 2225
rect 22855 2277 22907 2283
rect 21275 2265 21281 2273
rect 22849 2265 22855 2273
rect 21275 2237 22855 2265
rect 21275 2230 21281 2237
rect 22849 2230 22855 2237
rect 21223 2219 21275 2225
rect 24487 2277 24539 2283
rect 22907 2265 22913 2273
rect 24481 2265 24487 2273
rect 22907 2237 24487 2265
rect 22907 2230 22913 2237
rect 24481 2230 24487 2237
rect 22855 2219 22907 2225
rect 26119 2277 26171 2283
rect 24539 2265 24545 2273
rect 26113 2265 26119 2273
rect 24539 2237 26119 2265
rect 24539 2230 24545 2237
rect 26113 2230 26119 2237
rect 24487 2219 24539 2225
rect 27751 2277 27803 2283
rect 26171 2265 26177 2273
rect 27745 2265 27751 2273
rect 26171 2237 27751 2265
rect 26171 2230 26177 2237
rect 27745 2230 27751 2237
rect 26119 2219 26171 2225
rect 29383 2277 29435 2283
rect 27803 2265 27809 2273
rect 29377 2265 29383 2273
rect 27803 2237 29383 2265
rect 27803 2230 27809 2237
rect 29377 2230 29383 2237
rect 27751 2219 27803 2225
rect 31015 2277 31067 2283
rect 29435 2265 29441 2273
rect 31009 2265 31015 2273
rect 29435 2237 31015 2265
rect 29435 2230 29441 2237
rect 31009 2230 31015 2237
rect 29383 2219 29435 2225
rect 32647 2277 32699 2283
rect 31067 2265 31073 2273
rect 32641 2265 32647 2273
rect 31067 2237 32647 2265
rect 31067 2230 31073 2237
rect 32641 2230 32647 2237
rect 31015 2219 31067 2225
rect 34279 2277 34331 2283
rect 32699 2265 32705 2273
rect 34273 2265 34279 2273
rect 32699 2237 34279 2265
rect 32699 2230 32705 2237
rect 34273 2230 34279 2237
rect 32647 2219 32699 2225
rect 35911 2277 35963 2283
rect 34331 2265 34337 2273
rect 35905 2265 35911 2273
rect 34331 2237 35911 2265
rect 34331 2230 34337 2237
rect 35905 2230 35911 2237
rect 34279 2219 34331 2225
rect 37543 2277 37595 2283
rect 35963 2265 35969 2273
rect 37537 2265 37543 2273
rect 35963 2237 37543 2265
rect 35963 2230 35969 2237
rect 37537 2230 37543 2237
rect 35911 2219 35963 2225
rect 39175 2277 39227 2283
rect 37595 2265 37601 2273
rect 39169 2265 39175 2273
rect 37595 2237 39175 2265
rect 37595 2230 37601 2237
rect 39169 2230 39175 2237
rect 37543 2219 37595 2225
rect 40807 2277 40859 2283
rect 39227 2265 39233 2273
rect 40801 2265 40807 2273
rect 39227 2237 40807 2265
rect 39227 2230 39233 2237
rect 40801 2230 40807 2237
rect 39175 2219 39227 2225
rect 42439 2277 42491 2283
rect 40859 2265 40865 2273
rect 42433 2265 42439 2273
rect 40859 2237 42439 2265
rect 40859 2230 40865 2237
rect 42433 2230 42439 2237
rect 40807 2219 40859 2225
rect 44071 2277 44123 2283
rect 42491 2265 42497 2273
rect 44065 2265 44071 2273
rect 42491 2237 44071 2265
rect 42491 2230 42497 2237
rect 44065 2230 44071 2237
rect 42439 2219 42491 2225
rect 45703 2277 45755 2283
rect 44123 2265 44129 2273
rect 45697 2265 45703 2273
rect 44123 2237 45703 2265
rect 44123 2230 44129 2237
rect 45697 2230 45703 2237
rect 44071 2219 44123 2225
rect 47335 2277 47387 2283
rect 45755 2265 45761 2273
rect 47329 2265 47335 2273
rect 45755 2237 47335 2265
rect 45755 2230 45761 2237
rect 47329 2230 47335 2237
rect 45703 2219 45755 2225
rect 48967 2277 49019 2283
rect 47387 2265 47393 2273
rect 48961 2265 48967 2273
rect 47387 2237 48967 2265
rect 47387 2230 47393 2237
rect 48961 2230 48967 2237
rect 47335 2219 47387 2225
rect 50599 2277 50651 2283
rect 49019 2265 49025 2273
rect 50593 2265 50599 2273
rect 49019 2237 50599 2265
rect 49019 2230 49025 2237
rect 50593 2230 50599 2237
rect 48967 2219 49019 2225
rect 52231 2277 52283 2283
rect 50651 2265 50657 2273
rect 52225 2265 52231 2273
rect 50651 2237 52231 2265
rect 50651 2230 50657 2237
rect 52225 2230 52231 2237
rect 50599 2219 50651 2225
rect 52283 2230 52289 2273
rect 52231 2219 52283 2225
rect 7 2073 59 2079
rect 1 2026 7 2069
rect 1639 2073 1691 2079
rect 59 2061 65 2069
rect 1633 2061 1639 2069
rect 59 2033 1639 2061
rect 59 2026 65 2033
rect 1633 2026 1639 2033
rect 7 2015 59 2021
rect 3271 2073 3323 2079
rect 1691 2061 1697 2069
rect 3265 2061 3271 2069
rect 1691 2033 3271 2061
rect 1691 2026 1697 2033
rect 3265 2026 3271 2033
rect 1639 2015 1691 2021
rect 4903 2073 4955 2079
rect 3323 2061 3329 2069
rect 4897 2061 4903 2069
rect 3323 2033 4903 2061
rect 3323 2026 3329 2033
rect 4897 2026 4903 2033
rect 3271 2015 3323 2021
rect 6535 2073 6587 2079
rect 4955 2061 4961 2069
rect 6529 2061 6535 2069
rect 4955 2033 6535 2061
rect 4955 2026 4961 2033
rect 6529 2026 6535 2033
rect 4903 2015 4955 2021
rect 8167 2073 8219 2079
rect 6587 2061 6593 2069
rect 8161 2061 8167 2069
rect 6587 2033 8167 2061
rect 6587 2026 6593 2033
rect 8161 2026 8167 2033
rect 6535 2015 6587 2021
rect 9799 2073 9851 2079
rect 8219 2061 8225 2069
rect 9793 2061 9799 2069
rect 8219 2033 9799 2061
rect 8219 2026 8225 2033
rect 9793 2026 9799 2033
rect 8167 2015 8219 2021
rect 11431 2073 11483 2079
rect 9851 2061 9857 2069
rect 11425 2061 11431 2069
rect 9851 2033 11431 2061
rect 9851 2026 9857 2033
rect 11425 2026 11431 2033
rect 9799 2015 9851 2021
rect 13063 2073 13115 2079
rect 11483 2061 11489 2069
rect 13057 2061 13063 2069
rect 11483 2033 13063 2061
rect 11483 2026 11489 2033
rect 13057 2026 13063 2033
rect 11431 2015 11483 2021
rect 14695 2073 14747 2079
rect 13115 2061 13121 2069
rect 14689 2061 14695 2069
rect 13115 2033 14695 2061
rect 13115 2026 13121 2033
rect 14689 2026 14695 2033
rect 13063 2015 13115 2021
rect 16327 2073 16379 2079
rect 14747 2061 14753 2069
rect 16321 2061 16327 2069
rect 14747 2033 16327 2061
rect 14747 2026 14753 2033
rect 16321 2026 16327 2033
rect 14695 2015 14747 2021
rect 17959 2073 18011 2079
rect 16379 2061 16385 2069
rect 17953 2061 17959 2069
rect 16379 2033 17959 2061
rect 16379 2026 16385 2033
rect 17953 2026 17959 2033
rect 16327 2015 16379 2021
rect 19591 2073 19643 2079
rect 18011 2061 18017 2069
rect 19585 2061 19591 2069
rect 18011 2033 19591 2061
rect 18011 2026 18017 2033
rect 19585 2026 19591 2033
rect 17959 2015 18011 2021
rect 21223 2073 21275 2079
rect 19643 2061 19649 2069
rect 21217 2061 21223 2069
rect 19643 2033 21223 2061
rect 19643 2026 19649 2033
rect 21217 2026 21223 2033
rect 19591 2015 19643 2021
rect 22855 2073 22907 2079
rect 21275 2061 21281 2069
rect 22849 2061 22855 2069
rect 21275 2033 22855 2061
rect 21275 2026 21281 2033
rect 22849 2026 22855 2033
rect 21223 2015 21275 2021
rect 24487 2073 24539 2079
rect 22907 2061 22913 2069
rect 24481 2061 24487 2069
rect 22907 2033 24487 2061
rect 22907 2026 22913 2033
rect 24481 2026 24487 2033
rect 22855 2015 22907 2021
rect 26119 2073 26171 2079
rect 24539 2061 24545 2069
rect 26113 2061 26119 2069
rect 24539 2033 26119 2061
rect 24539 2026 24545 2033
rect 26113 2026 26119 2033
rect 24487 2015 24539 2021
rect 27751 2073 27803 2079
rect 26171 2061 26177 2069
rect 27745 2061 27751 2069
rect 26171 2033 27751 2061
rect 26171 2026 26177 2033
rect 27745 2026 27751 2033
rect 26119 2015 26171 2021
rect 29383 2073 29435 2079
rect 27803 2061 27809 2069
rect 29377 2061 29383 2069
rect 27803 2033 29383 2061
rect 27803 2026 27809 2033
rect 29377 2026 29383 2033
rect 27751 2015 27803 2021
rect 31015 2073 31067 2079
rect 29435 2061 29441 2069
rect 31009 2061 31015 2069
rect 29435 2033 31015 2061
rect 29435 2026 29441 2033
rect 31009 2026 31015 2033
rect 29383 2015 29435 2021
rect 32647 2073 32699 2079
rect 31067 2061 31073 2069
rect 32641 2061 32647 2069
rect 31067 2033 32647 2061
rect 31067 2026 31073 2033
rect 32641 2026 32647 2033
rect 31015 2015 31067 2021
rect 34279 2073 34331 2079
rect 32699 2061 32705 2069
rect 34273 2061 34279 2069
rect 32699 2033 34279 2061
rect 32699 2026 32705 2033
rect 34273 2026 34279 2033
rect 32647 2015 32699 2021
rect 35911 2073 35963 2079
rect 34331 2061 34337 2069
rect 35905 2061 35911 2069
rect 34331 2033 35911 2061
rect 34331 2026 34337 2033
rect 35905 2026 35911 2033
rect 34279 2015 34331 2021
rect 37543 2073 37595 2079
rect 35963 2061 35969 2069
rect 37537 2061 37543 2069
rect 35963 2033 37543 2061
rect 35963 2026 35969 2033
rect 37537 2026 37543 2033
rect 35911 2015 35963 2021
rect 39175 2073 39227 2079
rect 37595 2061 37601 2069
rect 39169 2061 39175 2069
rect 37595 2033 39175 2061
rect 37595 2026 37601 2033
rect 39169 2026 39175 2033
rect 37543 2015 37595 2021
rect 40807 2073 40859 2079
rect 39227 2061 39233 2069
rect 40801 2061 40807 2069
rect 39227 2033 40807 2061
rect 39227 2026 39233 2033
rect 40801 2026 40807 2033
rect 39175 2015 39227 2021
rect 42439 2073 42491 2079
rect 40859 2061 40865 2069
rect 42433 2061 42439 2069
rect 40859 2033 42439 2061
rect 40859 2026 40865 2033
rect 42433 2026 42439 2033
rect 40807 2015 40859 2021
rect 44071 2073 44123 2079
rect 42491 2061 42497 2069
rect 44065 2061 44071 2069
rect 42491 2033 44071 2061
rect 42491 2026 42497 2033
rect 44065 2026 44071 2033
rect 42439 2015 42491 2021
rect 45703 2073 45755 2079
rect 44123 2061 44129 2069
rect 45697 2061 45703 2069
rect 44123 2033 45703 2061
rect 44123 2026 44129 2033
rect 45697 2026 45703 2033
rect 44071 2015 44123 2021
rect 47335 2073 47387 2079
rect 45755 2061 45761 2069
rect 47329 2061 47335 2069
rect 45755 2033 47335 2061
rect 45755 2026 45761 2033
rect 47329 2026 47335 2033
rect 45703 2015 45755 2021
rect 48967 2073 49019 2079
rect 47387 2061 47393 2069
rect 48961 2061 48967 2069
rect 47387 2033 48967 2061
rect 47387 2026 47393 2033
rect 48961 2026 48967 2033
rect 47335 2015 47387 2021
rect 50599 2073 50651 2079
rect 49019 2061 49025 2069
rect 50593 2061 50599 2069
rect 49019 2033 50599 2061
rect 49019 2026 49025 2033
rect 50593 2026 50599 2033
rect 48967 2015 49019 2021
rect 52231 2073 52283 2079
rect 50651 2061 50657 2069
rect 52225 2061 52231 2069
rect 50651 2033 52231 2061
rect 50651 2026 50657 2033
rect 52225 2026 52231 2033
rect 50599 2015 50651 2021
rect 52283 2026 52289 2069
rect 52231 2015 52283 2021
rect 7 1869 59 1875
rect 1 1822 7 1865
rect 1639 1869 1691 1875
rect 59 1857 65 1865
rect 1633 1857 1639 1865
rect 59 1829 1639 1857
rect 59 1822 65 1829
rect 1633 1822 1639 1829
rect 7 1811 59 1817
rect 3271 1869 3323 1875
rect 1691 1857 1697 1865
rect 3265 1857 3271 1865
rect 1691 1829 3271 1857
rect 1691 1822 1697 1829
rect 3265 1822 3271 1829
rect 1639 1811 1691 1817
rect 4903 1869 4955 1875
rect 3323 1857 3329 1865
rect 4897 1857 4903 1865
rect 3323 1829 4903 1857
rect 3323 1822 3329 1829
rect 4897 1822 4903 1829
rect 3271 1811 3323 1817
rect 6535 1869 6587 1875
rect 4955 1857 4961 1865
rect 6529 1857 6535 1865
rect 4955 1829 6535 1857
rect 4955 1822 4961 1829
rect 6529 1822 6535 1829
rect 4903 1811 4955 1817
rect 8167 1869 8219 1875
rect 6587 1857 6593 1865
rect 8161 1857 8167 1865
rect 6587 1829 8167 1857
rect 6587 1822 6593 1829
rect 8161 1822 8167 1829
rect 6535 1811 6587 1817
rect 9799 1869 9851 1875
rect 8219 1857 8225 1865
rect 9793 1857 9799 1865
rect 8219 1829 9799 1857
rect 8219 1822 8225 1829
rect 9793 1822 9799 1829
rect 8167 1811 8219 1817
rect 11431 1869 11483 1875
rect 9851 1857 9857 1865
rect 11425 1857 11431 1865
rect 9851 1829 11431 1857
rect 9851 1822 9857 1829
rect 11425 1822 11431 1829
rect 9799 1811 9851 1817
rect 13063 1869 13115 1875
rect 11483 1857 11489 1865
rect 13057 1857 13063 1865
rect 11483 1829 13063 1857
rect 11483 1822 11489 1829
rect 13057 1822 13063 1829
rect 11431 1811 11483 1817
rect 14695 1869 14747 1875
rect 13115 1857 13121 1865
rect 14689 1857 14695 1865
rect 13115 1829 14695 1857
rect 13115 1822 13121 1829
rect 14689 1822 14695 1829
rect 13063 1811 13115 1817
rect 16327 1869 16379 1875
rect 14747 1857 14753 1865
rect 16321 1857 16327 1865
rect 14747 1829 16327 1857
rect 14747 1822 14753 1829
rect 16321 1822 16327 1829
rect 14695 1811 14747 1817
rect 17959 1869 18011 1875
rect 16379 1857 16385 1865
rect 17953 1857 17959 1865
rect 16379 1829 17959 1857
rect 16379 1822 16385 1829
rect 17953 1822 17959 1829
rect 16327 1811 16379 1817
rect 19591 1869 19643 1875
rect 18011 1857 18017 1865
rect 19585 1857 19591 1865
rect 18011 1829 19591 1857
rect 18011 1822 18017 1829
rect 19585 1822 19591 1829
rect 17959 1811 18011 1817
rect 21223 1869 21275 1875
rect 19643 1857 19649 1865
rect 21217 1857 21223 1865
rect 19643 1829 21223 1857
rect 19643 1822 19649 1829
rect 21217 1822 21223 1829
rect 19591 1811 19643 1817
rect 22855 1869 22907 1875
rect 21275 1857 21281 1865
rect 22849 1857 22855 1865
rect 21275 1829 22855 1857
rect 21275 1822 21281 1829
rect 22849 1822 22855 1829
rect 21223 1811 21275 1817
rect 24487 1869 24539 1875
rect 22907 1857 22913 1865
rect 24481 1857 24487 1865
rect 22907 1829 24487 1857
rect 22907 1822 22913 1829
rect 24481 1822 24487 1829
rect 22855 1811 22907 1817
rect 26119 1869 26171 1875
rect 24539 1857 24545 1865
rect 26113 1857 26119 1865
rect 24539 1829 26119 1857
rect 24539 1822 24545 1829
rect 26113 1822 26119 1829
rect 24487 1811 24539 1817
rect 27751 1869 27803 1875
rect 26171 1857 26177 1865
rect 27745 1857 27751 1865
rect 26171 1829 27751 1857
rect 26171 1822 26177 1829
rect 27745 1822 27751 1829
rect 26119 1811 26171 1817
rect 29383 1869 29435 1875
rect 27803 1857 27809 1865
rect 29377 1857 29383 1865
rect 27803 1829 29383 1857
rect 27803 1822 27809 1829
rect 29377 1822 29383 1829
rect 27751 1811 27803 1817
rect 31015 1869 31067 1875
rect 29435 1857 29441 1865
rect 31009 1857 31015 1865
rect 29435 1829 31015 1857
rect 29435 1822 29441 1829
rect 31009 1822 31015 1829
rect 29383 1811 29435 1817
rect 32647 1869 32699 1875
rect 31067 1857 31073 1865
rect 32641 1857 32647 1865
rect 31067 1829 32647 1857
rect 31067 1822 31073 1829
rect 32641 1822 32647 1829
rect 31015 1811 31067 1817
rect 34279 1869 34331 1875
rect 32699 1857 32705 1865
rect 34273 1857 34279 1865
rect 32699 1829 34279 1857
rect 32699 1822 32705 1829
rect 34273 1822 34279 1829
rect 32647 1811 32699 1817
rect 35911 1869 35963 1875
rect 34331 1857 34337 1865
rect 35905 1857 35911 1865
rect 34331 1829 35911 1857
rect 34331 1822 34337 1829
rect 35905 1822 35911 1829
rect 34279 1811 34331 1817
rect 37543 1869 37595 1875
rect 35963 1857 35969 1865
rect 37537 1857 37543 1865
rect 35963 1829 37543 1857
rect 35963 1822 35969 1829
rect 37537 1822 37543 1829
rect 35911 1811 35963 1817
rect 39175 1869 39227 1875
rect 37595 1857 37601 1865
rect 39169 1857 39175 1865
rect 37595 1829 39175 1857
rect 37595 1822 37601 1829
rect 39169 1822 39175 1829
rect 37543 1811 37595 1817
rect 40807 1869 40859 1875
rect 39227 1857 39233 1865
rect 40801 1857 40807 1865
rect 39227 1829 40807 1857
rect 39227 1822 39233 1829
rect 40801 1822 40807 1829
rect 39175 1811 39227 1817
rect 42439 1869 42491 1875
rect 40859 1857 40865 1865
rect 42433 1857 42439 1865
rect 40859 1829 42439 1857
rect 40859 1822 40865 1829
rect 42433 1822 42439 1829
rect 40807 1811 40859 1817
rect 44071 1869 44123 1875
rect 42491 1857 42497 1865
rect 44065 1857 44071 1865
rect 42491 1829 44071 1857
rect 42491 1822 42497 1829
rect 44065 1822 44071 1829
rect 42439 1811 42491 1817
rect 45703 1869 45755 1875
rect 44123 1857 44129 1865
rect 45697 1857 45703 1865
rect 44123 1829 45703 1857
rect 44123 1822 44129 1829
rect 45697 1822 45703 1829
rect 44071 1811 44123 1817
rect 47335 1869 47387 1875
rect 45755 1857 45761 1865
rect 47329 1857 47335 1865
rect 45755 1829 47335 1857
rect 45755 1822 45761 1829
rect 47329 1822 47335 1829
rect 45703 1811 45755 1817
rect 48967 1869 49019 1875
rect 47387 1857 47393 1865
rect 48961 1857 48967 1865
rect 47387 1829 48967 1857
rect 47387 1822 47393 1829
rect 48961 1822 48967 1829
rect 47335 1811 47387 1817
rect 50599 1869 50651 1875
rect 49019 1857 49025 1865
rect 50593 1857 50599 1865
rect 49019 1829 50599 1857
rect 49019 1822 49025 1829
rect 50593 1822 50599 1829
rect 48967 1811 49019 1817
rect 52231 1869 52283 1875
rect 50651 1857 50657 1865
rect 52225 1857 52231 1865
rect 50651 1829 52231 1857
rect 50651 1822 50657 1829
rect 52225 1822 52231 1829
rect 50599 1811 50651 1817
rect 52283 1822 52289 1865
rect 52231 1811 52283 1817
rect 7 1665 59 1671
rect 1 1618 7 1661
rect 1639 1665 1691 1671
rect 59 1653 65 1661
rect 1633 1653 1639 1661
rect 59 1625 1639 1653
rect 59 1618 65 1625
rect 1633 1618 1639 1625
rect 7 1607 59 1613
rect 3271 1665 3323 1671
rect 1691 1653 1697 1661
rect 3265 1653 3271 1661
rect 1691 1625 3271 1653
rect 1691 1618 1697 1625
rect 3265 1618 3271 1625
rect 1639 1607 1691 1613
rect 4903 1665 4955 1671
rect 3323 1653 3329 1661
rect 4897 1653 4903 1661
rect 3323 1625 4903 1653
rect 3323 1618 3329 1625
rect 4897 1618 4903 1625
rect 3271 1607 3323 1613
rect 6535 1665 6587 1671
rect 4955 1653 4961 1661
rect 6529 1653 6535 1661
rect 4955 1625 6535 1653
rect 4955 1618 4961 1625
rect 6529 1618 6535 1625
rect 4903 1607 4955 1613
rect 8167 1665 8219 1671
rect 6587 1653 6593 1661
rect 8161 1653 8167 1661
rect 6587 1625 8167 1653
rect 6587 1618 6593 1625
rect 8161 1618 8167 1625
rect 6535 1607 6587 1613
rect 9799 1665 9851 1671
rect 8219 1653 8225 1661
rect 9793 1653 9799 1661
rect 8219 1625 9799 1653
rect 8219 1618 8225 1625
rect 9793 1618 9799 1625
rect 8167 1607 8219 1613
rect 11431 1665 11483 1671
rect 9851 1653 9857 1661
rect 11425 1653 11431 1661
rect 9851 1625 11431 1653
rect 9851 1618 9857 1625
rect 11425 1618 11431 1625
rect 9799 1607 9851 1613
rect 13063 1665 13115 1671
rect 11483 1653 11489 1661
rect 13057 1653 13063 1661
rect 11483 1625 13063 1653
rect 11483 1618 11489 1625
rect 13057 1618 13063 1625
rect 11431 1607 11483 1613
rect 14695 1665 14747 1671
rect 13115 1653 13121 1661
rect 14689 1653 14695 1661
rect 13115 1625 14695 1653
rect 13115 1618 13121 1625
rect 14689 1618 14695 1625
rect 13063 1607 13115 1613
rect 16327 1665 16379 1671
rect 14747 1653 14753 1661
rect 16321 1653 16327 1661
rect 14747 1625 16327 1653
rect 14747 1618 14753 1625
rect 16321 1618 16327 1625
rect 14695 1607 14747 1613
rect 17959 1665 18011 1671
rect 16379 1653 16385 1661
rect 17953 1653 17959 1661
rect 16379 1625 17959 1653
rect 16379 1618 16385 1625
rect 17953 1618 17959 1625
rect 16327 1607 16379 1613
rect 19591 1665 19643 1671
rect 18011 1653 18017 1661
rect 19585 1653 19591 1661
rect 18011 1625 19591 1653
rect 18011 1618 18017 1625
rect 19585 1618 19591 1625
rect 17959 1607 18011 1613
rect 21223 1665 21275 1671
rect 19643 1653 19649 1661
rect 21217 1653 21223 1661
rect 19643 1625 21223 1653
rect 19643 1618 19649 1625
rect 21217 1618 21223 1625
rect 19591 1607 19643 1613
rect 22855 1665 22907 1671
rect 21275 1653 21281 1661
rect 22849 1653 22855 1661
rect 21275 1625 22855 1653
rect 21275 1618 21281 1625
rect 22849 1618 22855 1625
rect 21223 1607 21275 1613
rect 24487 1665 24539 1671
rect 22907 1653 22913 1661
rect 24481 1653 24487 1661
rect 22907 1625 24487 1653
rect 22907 1618 22913 1625
rect 24481 1618 24487 1625
rect 22855 1607 22907 1613
rect 26119 1665 26171 1671
rect 24539 1653 24545 1661
rect 26113 1653 26119 1661
rect 24539 1625 26119 1653
rect 24539 1618 24545 1625
rect 26113 1618 26119 1625
rect 24487 1607 24539 1613
rect 27751 1665 27803 1671
rect 26171 1653 26177 1661
rect 27745 1653 27751 1661
rect 26171 1625 27751 1653
rect 26171 1618 26177 1625
rect 27745 1618 27751 1625
rect 26119 1607 26171 1613
rect 29383 1665 29435 1671
rect 27803 1653 27809 1661
rect 29377 1653 29383 1661
rect 27803 1625 29383 1653
rect 27803 1618 27809 1625
rect 29377 1618 29383 1625
rect 27751 1607 27803 1613
rect 31015 1665 31067 1671
rect 29435 1653 29441 1661
rect 31009 1653 31015 1661
rect 29435 1625 31015 1653
rect 29435 1618 29441 1625
rect 31009 1618 31015 1625
rect 29383 1607 29435 1613
rect 32647 1665 32699 1671
rect 31067 1653 31073 1661
rect 32641 1653 32647 1661
rect 31067 1625 32647 1653
rect 31067 1618 31073 1625
rect 32641 1618 32647 1625
rect 31015 1607 31067 1613
rect 34279 1665 34331 1671
rect 32699 1653 32705 1661
rect 34273 1653 34279 1661
rect 32699 1625 34279 1653
rect 32699 1618 32705 1625
rect 34273 1618 34279 1625
rect 32647 1607 32699 1613
rect 35911 1665 35963 1671
rect 34331 1653 34337 1661
rect 35905 1653 35911 1661
rect 34331 1625 35911 1653
rect 34331 1618 34337 1625
rect 35905 1618 35911 1625
rect 34279 1607 34331 1613
rect 37543 1665 37595 1671
rect 35963 1653 35969 1661
rect 37537 1653 37543 1661
rect 35963 1625 37543 1653
rect 35963 1618 35969 1625
rect 37537 1618 37543 1625
rect 35911 1607 35963 1613
rect 39175 1665 39227 1671
rect 37595 1653 37601 1661
rect 39169 1653 39175 1661
rect 37595 1625 39175 1653
rect 37595 1618 37601 1625
rect 39169 1618 39175 1625
rect 37543 1607 37595 1613
rect 40807 1665 40859 1671
rect 39227 1653 39233 1661
rect 40801 1653 40807 1661
rect 39227 1625 40807 1653
rect 39227 1618 39233 1625
rect 40801 1618 40807 1625
rect 39175 1607 39227 1613
rect 42439 1665 42491 1671
rect 40859 1653 40865 1661
rect 42433 1653 42439 1661
rect 40859 1625 42439 1653
rect 40859 1618 40865 1625
rect 42433 1618 42439 1625
rect 40807 1607 40859 1613
rect 44071 1665 44123 1671
rect 42491 1653 42497 1661
rect 44065 1653 44071 1661
rect 42491 1625 44071 1653
rect 42491 1618 42497 1625
rect 44065 1618 44071 1625
rect 42439 1607 42491 1613
rect 45703 1665 45755 1671
rect 44123 1653 44129 1661
rect 45697 1653 45703 1661
rect 44123 1625 45703 1653
rect 44123 1618 44129 1625
rect 45697 1618 45703 1625
rect 44071 1607 44123 1613
rect 47335 1665 47387 1671
rect 45755 1653 45761 1661
rect 47329 1653 47335 1661
rect 45755 1625 47335 1653
rect 45755 1618 45761 1625
rect 47329 1618 47335 1625
rect 45703 1607 45755 1613
rect 48967 1665 49019 1671
rect 47387 1653 47393 1661
rect 48961 1653 48967 1661
rect 47387 1625 48967 1653
rect 47387 1618 47393 1625
rect 48961 1618 48967 1625
rect 47335 1607 47387 1613
rect 50599 1665 50651 1671
rect 49019 1653 49025 1661
rect 50593 1653 50599 1661
rect 49019 1625 50599 1653
rect 49019 1618 49025 1625
rect 50593 1618 50599 1625
rect 48967 1607 49019 1613
rect 52231 1665 52283 1671
rect 50651 1653 50657 1661
rect 52225 1653 52231 1661
rect 50651 1625 52231 1653
rect 50651 1618 50657 1625
rect 52225 1618 52231 1625
rect 50599 1607 50651 1613
rect 52283 1618 52289 1661
rect 52231 1607 52283 1613
rect 7 1461 59 1467
rect 1 1414 7 1457
rect 1639 1461 1691 1467
rect 59 1449 65 1457
rect 1633 1449 1639 1457
rect 59 1421 1639 1449
rect 59 1414 65 1421
rect 1633 1414 1639 1421
rect 7 1403 59 1409
rect 3271 1461 3323 1467
rect 1691 1449 1697 1457
rect 3265 1449 3271 1457
rect 1691 1421 3271 1449
rect 1691 1414 1697 1421
rect 3265 1414 3271 1421
rect 1639 1403 1691 1409
rect 4903 1461 4955 1467
rect 3323 1449 3329 1457
rect 4897 1449 4903 1457
rect 3323 1421 4903 1449
rect 3323 1414 3329 1421
rect 4897 1414 4903 1421
rect 3271 1403 3323 1409
rect 6535 1461 6587 1467
rect 4955 1449 4961 1457
rect 6529 1449 6535 1457
rect 4955 1421 6535 1449
rect 4955 1414 4961 1421
rect 6529 1414 6535 1421
rect 4903 1403 4955 1409
rect 8167 1461 8219 1467
rect 6587 1449 6593 1457
rect 8161 1449 8167 1457
rect 6587 1421 8167 1449
rect 6587 1414 6593 1421
rect 8161 1414 8167 1421
rect 6535 1403 6587 1409
rect 9799 1461 9851 1467
rect 8219 1449 8225 1457
rect 9793 1449 9799 1457
rect 8219 1421 9799 1449
rect 8219 1414 8225 1421
rect 9793 1414 9799 1421
rect 8167 1403 8219 1409
rect 11431 1461 11483 1467
rect 9851 1449 9857 1457
rect 11425 1449 11431 1457
rect 9851 1421 11431 1449
rect 9851 1414 9857 1421
rect 11425 1414 11431 1421
rect 9799 1403 9851 1409
rect 13063 1461 13115 1467
rect 11483 1449 11489 1457
rect 13057 1449 13063 1457
rect 11483 1421 13063 1449
rect 11483 1414 11489 1421
rect 13057 1414 13063 1421
rect 11431 1403 11483 1409
rect 14695 1461 14747 1467
rect 13115 1449 13121 1457
rect 14689 1449 14695 1457
rect 13115 1421 14695 1449
rect 13115 1414 13121 1421
rect 14689 1414 14695 1421
rect 13063 1403 13115 1409
rect 16327 1461 16379 1467
rect 14747 1449 14753 1457
rect 16321 1449 16327 1457
rect 14747 1421 16327 1449
rect 14747 1414 14753 1421
rect 16321 1414 16327 1421
rect 14695 1403 14747 1409
rect 17959 1461 18011 1467
rect 16379 1449 16385 1457
rect 17953 1449 17959 1457
rect 16379 1421 17959 1449
rect 16379 1414 16385 1421
rect 17953 1414 17959 1421
rect 16327 1403 16379 1409
rect 19591 1461 19643 1467
rect 18011 1449 18017 1457
rect 19585 1449 19591 1457
rect 18011 1421 19591 1449
rect 18011 1414 18017 1421
rect 19585 1414 19591 1421
rect 17959 1403 18011 1409
rect 21223 1461 21275 1467
rect 19643 1449 19649 1457
rect 21217 1449 21223 1457
rect 19643 1421 21223 1449
rect 19643 1414 19649 1421
rect 21217 1414 21223 1421
rect 19591 1403 19643 1409
rect 22855 1461 22907 1467
rect 21275 1449 21281 1457
rect 22849 1449 22855 1457
rect 21275 1421 22855 1449
rect 21275 1414 21281 1421
rect 22849 1414 22855 1421
rect 21223 1403 21275 1409
rect 24487 1461 24539 1467
rect 22907 1449 22913 1457
rect 24481 1449 24487 1457
rect 22907 1421 24487 1449
rect 22907 1414 22913 1421
rect 24481 1414 24487 1421
rect 22855 1403 22907 1409
rect 26119 1461 26171 1467
rect 24539 1449 24545 1457
rect 26113 1449 26119 1457
rect 24539 1421 26119 1449
rect 24539 1414 24545 1421
rect 26113 1414 26119 1421
rect 24487 1403 24539 1409
rect 27751 1461 27803 1467
rect 26171 1449 26177 1457
rect 27745 1449 27751 1457
rect 26171 1421 27751 1449
rect 26171 1414 26177 1421
rect 27745 1414 27751 1421
rect 26119 1403 26171 1409
rect 29383 1461 29435 1467
rect 27803 1449 27809 1457
rect 29377 1449 29383 1457
rect 27803 1421 29383 1449
rect 27803 1414 27809 1421
rect 29377 1414 29383 1421
rect 27751 1403 27803 1409
rect 31015 1461 31067 1467
rect 29435 1449 29441 1457
rect 31009 1449 31015 1457
rect 29435 1421 31015 1449
rect 29435 1414 29441 1421
rect 31009 1414 31015 1421
rect 29383 1403 29435 1409
rect 32647 1461 32699 1467
rect 31067 1449 31073 1457
rect 32641 1449 32647 1457
rect 31067 1421 32647 1449
rect 31067 1414 31073 1421
rect 32641 1414 32647 1421
rect 31015 1403 31067 1409
rect 34279 1461 34331 1467
rect 32699 1449 32705 1457
rect 34273 1449 34279 1457
rect 32699 1421 34279 1449
rect 32699 1414 32705 1421
rect 34273 1414 34279 1421
rect 32647 1403 32699 1409
rect 35911 1461 35963 1467
rect 34331 1449 34337 1457
rect 35905 1449 35911 1457
rect 34331 1421 35911 1449
rect 34331 1414 34337 1421
rect 35905 1414 35911 1421
rect 34279 1403 34331 1409
rect 37543 1461 37595 1467
rect 35963 1449 35969 1457
rect 37537 1449 37543 1457
rect 35963 1421 37543 1449
rect 35963 1414 35969 1421
rect 37537 1414 37543 1421
rect 35911 1403 35963 1409
rect 39175 1461 39227 1467
rect 37595 1449 37601 1457
rect 39169 1449 39175 1457
rect 37595 1421 39175 1449
rect 37595 1414 37601 1421
rect 39169 1414 39175 1421
rect 37543 1403 37595 1409
rect 40807 1461 40859 1467
rect 39227 1449 39233 1457
rect 40801 1449 40807 1457
rect 39227 1421 40807 1449
rect 39227 1414 39233 1421
rect 40801 1414 40807 1421
rect 39175 1403 39227 1409
rect 42439 1461 42491 1467
rect 40859 1449 40865 1457
rect 42433 1449 42439 1457
rect 40859 1421 42439 1449
rect 40859 1414 40865 1421
rect 42433 1414 42439 1421
rect 40807 1403 40859 1409
rect 44071 1461 44123 1467
rect 42491 1449 42497 1457
rect 44065 1449 44071 1457
rect 42491 1421 44071 1449
rect 42491 1414 42497 1421
rect 44065 1414 44071 1421
rect 42439 1403 42491 1409
rect 45703 1461 45755 1467
rect 44123 1449 44129 1457
rect 45697 1449 45703 1457
rect 44123 1421 45703 1449
rect 44123 1414 44129 1421
rect 45697 1414 45703 1421
rect 44071 1403 44123 1409
rect 47335 1461 47387 1467
rect 45755 1449 45761 1457
rect 47329 1449 47335 1457
rect 45755 1421 47335 1449
rect 45755 1414 45761 1421
rect 47329 1414 47335 1421
rect 45703 1403 45755 1409
rect 48967 1461 49019 1467
rect 47387 1449 47393 1457
rect 48961 1449 48967 1457
rect 47387 1421 48967 1449
rect 47387 1414 47393 1421
rect 48961 1414 48967 1421
rect 47335 1403 47387 1409
rect 50599 1461 50651 1467
rect 49019 1449 49025 1457
rect 50593 1449 50599 1457
rect 49019 1421 50599 1449
rect 49019 1414 49025 1421
rect 50593 1414 50599 1421
rect 48967 1403 49019 1409
rect 52231 1461 52283 1467
rect 50651 1449 50657 1457
rect 52225 1449 52231 1457
rect 50651 1421 52231 1449
rect 50651 1414 50657 1421
rect 52225 1414 52231 1421
rect 50599 1403 50651 1409
rect 52283 1414 52289 1457
rect 52231 1403 52283 1409
rect 7 1257 59 1263
rect 1 1210 7 1253
rect 1639 1257 1691 1263
rect 59 1245 65 1253
rect 1633 1245 1639 1253
rect 59 1217 1639 1245
rect 59 1210 65 1217
rect 1633 1210 1639 1217
rect 7 1199 59 1205
rect 3271 1257 3323 1263
rect 1691 1245 1697 1253
rect 3265 1245 3271 1253
rect 1691 1217 3271 1245
rect 1691 1210 1697 1217
rect 3265 1210 3271 1217
rect 1639 1199 1691 1205
rect 4903 1257 4955 1263
rect 3323 1245 3329 1253
rect 4897 1245 4903 1253
rect 3323 1217 4903 1245
rect 3323 1210 3329 1217
rect 4897 1210 4903 1217
rect 3271 1199 3323 1205
rect 6535 1257 6587 1263
rect 4955 1245 4961 1253
rect 6529 1245 6535 1253
rect 4955 1217 6535 1245
rect 4955 1210 4961 1217
rect 6529 1210 6535 1217
rect 4903 1199 4955 1205
rect 8167 1257 8219 1263
rect 6587 1245 6593 1253
rect 8161 1245 8167 1253
rect 6587 1217 8167 1245
rect 6587 1210 6593 1217
rect 8161 1210 8167 1217
rect 6535 1199 6587 1205
rect 9799 1257 9851 1263
rect 8219 1245 8225 1253
rect 9793 1245 9799 1253
rect 8219 1217 9799 1245
rect 8219 1210 8225 1217
rect 9793 1210 9799 1217
rect 8167 1199 8219 1205
rect 11431 1257 11483 1263
rect 9851 1245 9857 1253
rect 11425 1245 11431 1253
rect 9851 1217 11431 1245
rect 9851 1210 9857 1217
rect 11425 1210 11431 1217
rect 9799 1199 9851 1205
rect 13063 1257 13115 1263
rect 11483 1245 11489 1253
rect 13057 1245 13063 1253
rect 11483 1217 13063 1245
rect 11483 1210 11489 1217
rect 13057 1210 13063 1217
rect 11431 1199 11483 1205
rect 14695 1257 14747 1263
rect 13115 1245 13121 1253
rect 14689 1245 14695 1253
rect 13115 1217 14695 1245
rect 13115 1210 13121 1217
rect 14689 1210 14695 1217
rect 13063 1199 13115 1205
rect 16327 1257 16379 1263
rect 14747 1245 14753 1253
rect 16321 1245 16327 1253
rect 14747 1217 16327 1245
rect 14747 1210 14753 1217
rect 16321 1210 16327 1217
rect 14695 1199 14747 1205
rect 17959 1257 18011 1263
rect 16379 1245 16385 1253
rect 17953 1245 17959 1253
rect 16379 1217 17959 1245
rect 16379 1210 16385 1217
rect 17953 1210 17959 1217
rect 16327 1199 16379 1205
rect 19591 1257 19643 1263
rect 18011 1245 18017 1253
rect 19585 1245 19591 1253
rect 18011 1217 19591 1245
rect 18011 1210 18017 1217
rect 19585 1210 19591 1217
rect 17959 1199 18011 1205
rect 21223 1257 21275 1263
rect 19643 1245 19649 1253
rect 21217 1245 21223 1253
rect 19643 1217 21223 1245
rect 19643 1210 19649 1217
rect 21217 1210 21223 1217
rect 19591 1199 19643 1205
rect 22855 1257 22907 1263
rect 21275 1245 21281 1253
rect 22849 1245 22855 1253
rect 21275 1217 22855 1245
rect 21275 1210 21281 1217
rect 22849 1210 22855 1217
rect 21223 1199 21275 1205
rect 24487 1257 24539 1263
rect 22907 1245 22913 1253
rect 24481 1245 24487 1253
rect 22907 1217 24487 1245
rect 22907 1210 22913 1217
rect 24481 1210 24487 1217
rect 22855 1199 22907 1205
rect 26119 1257 26171 1263
rect 24539 1245 24545 1253
rect 26113 1245 26119 1253
rect 24539 1217 26119 1245
rect 24539 1210 24545 1217
rect 26113 1210 26119 1217
rect 24487 1199 24539 1205
rect 27751 1257 27803 1263
rect 26171 1245 26177 1253
rect 27745 1245 27751 1253
rect 26171 1217 27751 1245
rect 26171 1210 26177 1217
rect 27745 1210 27751 1217
rect 26119 1199 26171 1205
rect 29383 1257 29435 1263
rect 27803 1245 27809 1253
rect 29377 1245 29383 1253
rect 27803 1217 29383 1245
rect 27803 1210 27809 1217
rect 29377 1210 29383 1217
rect 27751 1199 27803 1205
rect 31015 1257 31067 1263
rect 29435 1245 29441 1253
rect 31009 1245 31015 1253
rect 29435 1217 31015 1245
rect 29435 1210 29441 1217
rect 31009 1210 31015 1217
rect 29383 1199 29435 1205
rect 32647 1257 32699 1263
rect 31067 1245 31073 1253
rect 32641 1245 32647 1253
rect 31067 1217 32647 1245
rect 31067 1210 31073 1217
rect 32641 1210 32647 1217
rect 31015 1199 31067 1205
rect 34279 1257 34331 1263
rect 32699 1245 32705 1253
rect 34273 1245 34279 1253
rect 32699 1217 34279 1245
rect 32699 1210 32705 1217
rect 34273 1210 34279 1217
rect 32647 1199 32699 1205
rect 35911 1257 35963 1263
rect 34331 1245 34337 1253
rect 35905 1245 35911 1253
rect 34331 1217 35911 1245
rect 34331 1210 34337 1217
rect 35905 1210 35911 1217
rect 34279 1199 34331 1205
rect 37543 1257 37595 1263
rect 35963 1245 35969 1253
rect 37537 1245 37543 1253
rect 35963 1217 37543 1245
rect 35963 1210 35969 1217
rect 37537 1210 37543 1217
rect 35911 1199 35963 1205
rect 39175 1257 39227 1263
rect 37595 1245 37601 1253
rect 39169 1245 39175 1253
rect 37595 1217 39175 1245
rect 37595 1210 37601 1217
rect 39169 1210 39175 1217
rect 37543 1199 37595 1205
rect 40807 1257 40859 1263
rect 39227 1245 39233 1253
rect 40801 1245 40807 1253
rect 39227 1217 40807 1245
rect 39227 1210 39233 1217
rect 40801 1210 40807 1217
rect 39175 1199 39227 1205
rect 42439 1257 42491 1263
rect 40859 1245 40865 1253
rect 42433 1245 42439 1253
rect 40859 1217 42439 1245
rect 40859 1210 40865 1217
rect 42433 1210 42439 1217
rect 40807 1199 40859 1205
rect 44071 1257 44123 1263
rect 42491 1245 42497 1253
rect 44065 1245 44071 1253
rect 42491 1217 44071 1245
rect 42491 1210 42497 1217
rect 44065 1210 44071 1217
rect 42439 1199 42491 1205
rect 45703 1257 45755 1263
rect 44123 1245 44129 1253
rect 45697 1245 45703 1253
rect 44123 1217 45703 1245
rect 44123 1210 44129 1217
rect 45697 1210 45703 1217
rect 44071 1199 44123 1205
rect 47335 1257 47387 1263
rect 45755 1245 45761 1253
rect 47329 1245 47335 1253
rect 45755 1217 47335 1245
rect 45755 1210 45761 1217
rect 47329 1210 47335 1217
rect 45703 1199 45755 1205
rect 48967 1257 49019 1263
rect 47387 1245 47393 1253
rect 48961 1245 48967 1253
rect 47387 1217 48967 1245
rect 47387 1210 47393 1217
rect 48961 1210 48967 1217
rect 47335 1199 47387 1205
rect 50599 1257 50651 1263
rect 49019 1245 49025 1253
rect 50593 1245 50599 1253
rect 49019 1217 50599 1245
rect 49019 1210 49025 1217
rect 50593 1210 50599 1217
rect 48967 1199 49019 1205
rect 52231 1257 52283 1263
rect 50651 1245 50657 1253
rect 52225 1245 52231 1253
rect 50651 1217 52231 1245
rect 50651 1210 50657 1217
rect 52225 1210 52231 1217
rect 50599 1199 50651 1205
rect 52283 1210 52289 1253
rect 52231 1199 52283 1205
rect 7 1053 59 1059
rect 1 1006 7 1049
rect 1639 1053 1691 1059
rect 59 1041 65 1049
rect 1633 1041 1639 1049
rect 59 1013 1639 1041
rect 59 1006 65 1013
rect 1633 1006 1639 1013
rect 7 995 59 1001
rect 3271 1053 3323 1059
rect 1691 1041 1697 1049
rect 3265 1041 3271 1049
rect 1691 1013 3271 1041
rect 1691 1006 1697 1013
rect 3265 1006 3271 1013
rect 1639 995 1691 1001
rect 4903 1053 4955 1059
rect 3323 1041 3329 1049
rect 4897 1041 4903 1049
rect 3323 1013 4903 1041
rect 3323 1006 3329 1013
rect 4897 1006 4903 1013
rect 3271 995 3323 1001
rect 6535 1053 6587 1059
rect 4955 1041 4961 1049
rect 6529 1041 6535 1049
rect 4955 1013 6535 1041
rect 4955 1006 4961 1013
rect 6529 1006 6535 1013
rect 4903 995 4955 1001
rect 8167 1053 8219 1059
rect 6587 1041 6593 1049
rect 8161 1041 8167 1049
rect 6587 1013 8167 1041
rect 6587 1006 6593 1013
rect 8161 1006 8167 1013
rect 6535 995 6587 1001
rect 9799 1053 9851 1059
rect 8219 1041 8225 1049
rect 9793 1041 9799 1049
rect 8219 1013 9799 1041
rect 8219 1006 8225 1013
rect 9793 1006 9799 1013
rect 8167 995 8219 1001
rect 11431 1053 11483 1059
rect 9851 1041 9857 1049
rect 11425 1041 11431 1049
rect 9851 1013 11431 1041
rect 9851 1006 9857 1013
rect 11425 1006 11431 1013
rect 9799 995 9851 1001
rect 13063 1053 13115 1059
rect 11483 1041 11489 1049
rect 13057 1041 13063 1049
rect 11483 1013 13063 1041
rect 11483 1006 11489 1013
rect 13057 1006 13063 1013
rect 11431 995 11483 1001
rect 14695 1053 14747 1059
rect 13115 1041 13121 1049
rect 14689 1041 14695 1049
rect 13115 1013 14695 1041
rect 13115 1006 13121 1013
rect 14689 1006 14695 1013
rect 13063 995 13115 1001
rect 16327 1053 16379 1059
rect 14747 1041 14753 1049
rect 16321 1041 16327 1049
rect 14747 1013 16327 1041
rect 14747 1006 14753 1013
rect 16321 1006 16327 1013
rect 14695 995 14747 1001
rect 17959 1053 18011 1059
rect 16379 1041 16385 1049
rect 17953 1041 17959 1049
rect 16379 1013 17959 1041
rect 16379 1006 16385 1013
rect 17953 1006 17959 1013
rect 16327 995 16379 1001
rect 19591 1053 19643 1059
rect 18011 1041 18017 1049
rect 19585 1041 19591 1049
rect 18011 1013 19591 1041
rect 18011 1006 18017 1013
rect 19585 1006 19591 1013
rect 17959 995 18011 1001
rect 21223 1053 21275 1059
rect 19643 1041 19649 1049
rect 21217 1041 21223 1049
rect 19643 1013 21223 1041
rect 19643 1006 19649 1013
rect 21217 1006 21223 1013
rect 19591 995 19643 1001
rect 22855 1053 22907 1059
rect 21275 1041 21281 1049
rect 22849 1041 22855 1049
rect 21275 1013 22855 1041
rect 21275 1006 21281 1013
rect 22849 1006 22855 1013
rect 21223 995 21275 1001
rect 24487 1053 24539 1059
rect 22907 1041 22913 1049
rect 24481 1041 24487 1049
rect 22907 1013 24487 1041
rect 22907 1006 22913 1013
rect 24481 1006 24487 1013
rect 22855 995 22907 1001
rect 26119 1053 26171 1059
rect 24539 1041 24545 1049
rect 26113 1041 26119 1049
rect 24539 1013 26119 1041
rect 24539 1006 24545 1013
rect 26113 1006 26119 1013
rect 24487 995 24539 1001
rect 27751 1053 27803 1059
rect 26171 1041 26177 1049
rect 27745 1041 27751 1049
rect 26171 1013 27751 1041
rect 26171 1006 26177 1013
rect 27745 1006 27751 1013
rect 26119 995 26171 1001
rect 29383 1053 29435 1059
rect 27803 1041 27809 1049
rect 29377 1041 29383 1049
rect 27803 1013 29383 1041
rect 27803 1006 27809 1013
rect 29377 1006 29383 1013
rect 27751 995 27803 1001
rect 31015 1053 31067 1059
rect 29435 1041 29441 1049
rect 31009 1041 31015 1049
rect 29435 1013 31015 1041
rect 29435 1006 29441 1013
rect 31009 1006 31015 1013
rect 29383 995 29435 1001
rect 32647 1053 32699 1059
rect 31067 1041 31073 1049
rect 32641 1041 32647 1049
rect 31067 1013 32647 1041
rect 31067 1006 31073 1013
rect 32641 1006 32647 1013
rect 31015 995 31067 1001
rect 34279 1053 34331 1059
rect 32699 1041 32705 1049
rect 34273 1041 34279 1049
rect 32699 1013 34279 1041
rect 32699 1006 32705 1013
rect 34273 1006 34279 1013
rect 32647 995 32699 1001
rect 35911 1053 35963 1059
rect 34331 1041 34337 1049
rect 35905 1041 35911 1049
rect 34331 1013 35911 1041
rect 34331 1006 34337 1013
rect 35905 1006 35911 1013
rect 34279 995 34331 1001
rect 37543 1053 37595 1059
rect 35963 1041 35969 1049
rect 37537 1041 37543 1049
rect 35963 1013 37543 1041
rect 35963 1006 35969 1013
rect 37537 1006 37543 1013
rect 35911 995 35963 1001
rect 39175 1053 39227 1059
rect 37595 1041 37601 1049
rect 39169 1041 39175 1049
rect 37595 1013 39175 1041
rect 37595 1006 37601 1013
rect 39169 1006 39175 1013
rect 37543 995 37595 1001
rect 40807 1053 40859 1059
rect 39227 1041 39233 1049
rect 40801 1041 40807 1049
rect 39227 1013 40807 1041
rect 39227 1006 39233 1013
rect 40801 1006 40807 1013
rect 39175 995 39227 1001
rect 42439 1053 42491 1059
rect 40859 1041 40865 1049
rect 42433 1041 42439 1049
rect 40859 1013 42439 1041
rect 40859 1006 40865 1013
rect 42433 1006 42439 1013
rect 40807 995 40859 1001
rect 44071 1053 44123 1059
rect 42491 1041 42497 1049
rect 44065 1041 44071 1049
rect 42491 1013 44071 1041
rect 42491 1006 42497 1013
rect 44065 1006 44071 1013
rect 42439 995 42491 1001
rect 45703 1053 45755 1059
rect 44123 1041 44129 1049
rect 45697 1041 45703 1049
rect 44123 1013 45703 1041
rect 44123 1006 44129 1013
rect 45697 1006 45703 1013
rect 44071 995 44123 1001
rect 47335 1053 47387 1059
rect 45755 1041 45761 1049
rect 47329 1041 47335 1049
rect 45755 1013 47335 1041
rect 45755 1006 45761 1013
rect 47329 1006 47335 1013
rect 45703 995 45755 1001
rect 48967 1053 49019 1059
rect 47387 1041 47393 1049
rect 48961 1041 48967 1049
rect 47387 1013 48967 1041
rect 47387 1006 47393 1013
rect 48961 1006 48967 1013
rect 47335 995 47387 1001
rect 50599 1053 50651 1059
rect 49019 1041 49025 1049
rect 50593 1041 50599 1049
rect 49019 1013 50599 1041
rect 49019 1006 49025 1013
rect 50593 1006 50599 1013
rect 48967 995 49019 1001
rect 52231 1053 52283 1059
rect 50651 1041 50657 1049
rect 52225 1041 52231 1049
rect 50651 1013 52231 1041
rect 50651 1006 50657 1013
rect 52225 1006 52231 1013
rect 50599 995 50651 1001
rect 52283 1006 52289 1049
rect 52231 995 52283 1001
rect 212 847 218 899
rect 270 887 276 899
rect 416 887 422 899
rect 270 859 422 887
rect 270 847 276 859
rect 416 847 422 859
rect 474 887 480 899
rect 620 887 626 899
rect 474 859 626 887
rect 474 847 480 859
rect 620 847 626 859
rect 678 887 684 899
rect 824 887 830 899
rect 678 859 830 887
rect 678 847 684 859
rect 824 847 830 859
rect 882 887 888 899
rect 1028 887 1034 899
rect 882 859 1034 887
rect 882 847 888 859
rect 1028 847 1034 859
rect 1086 887 1092 899
rect 1232 887 1238 899
rect 1086 859 1238 887
rect 1086 847 1092 859
rect 1232 847 1238 859
rect 1290 887 1296 899
rect 1436 887 1442 899
rect 1290 859 1442 887
rect 1290 847 1296 859
rect 1436 847 1442 859
rect 1494 887 1500 899
rect 1640 887 1646 899
rect 1494 859 1646 887
rect 1494 847 1500 859
rect 1640 847 1646 859
rect 1698 887 1704 899
rect 1844 887 1850 899
rect 1698 859 1850 887
rect 1698 847 1704 859
rect 1844 847 1850 859
rect 1902 887 1908 899
rect 2048 887 2054 899
rect 1902 859 2054 887
rect 1902 847 1908 859
rect 2048 847 2054 859
rect 2106 887 2112 899
rect 2252 887 2258 899
rect 2106 859 2258 887
rect 2106 847 2112 859
rect 2252 847 2258 859
rect 2310 887 2316 899
rect 2456 887 2462 899
rect 2310 859 2462 887
rect 2310 847 2316 859
rect 2456 847 2462 859
rect 2514 887 2520 899
rect 2660 887 2666 899
rect 2514 859 2666 887
rect 2514 847 2520 859
rect 2660 847 2666 859
rect 2718 887 2724 899
rect 2864 887 2870 899
rect 2718 859 2870 887
rect 2718 847 2724 859
rect 2864 847 2870 859
rect 2922 887 2928 899
rect 3068 887 3074 899
rect 2922 859 3074 887
rect 2922 847 2928 859
rect 3068 847 3074 859
rect 3126 887 3132 899
rect 3272 887 3278 899
rect 3126 859 3278 887
rect 3126 847 3132 859
rect 3272 847 3278 859
rect 3330 887 3336 899
rect 3476 887 3482 899
rect 3330 859 3482 887
rect 3330 847 3336 859
rect 3476 847 3482 859
rect 3534 887 3540 899
rect 3680 887 3686 899
rect 3534 859 3686 887
rect 3534 847 3540 859
rect 3680 847 3686 859
rect 3738 887 3744 899
rect 3884 887 3890 899
rect 3738 859 3890 887
rect 3738 847 3744 859
rect 3884 847 3890 859
rect 3942 887 3948 899
rect 4088 887 4094 899
rect 3942 859 4094 887
rect 3942 847 3948 859
rect 4088 847 4094 859
rect 4146 887 4152 899
rect 4292 887 4298 899
rect 4146 859 4298 887
rect 4146 847 4152 859
rect 4292 847 4298 859
rect 4350 887 4356 899
rect 4496 887 4502 899
rect 4350 859 4502 887
rect 4350 847 4356 859
rect 4496 847 4502 859
rect 4554 887 4560 899
rect 4700 887 4706 899
rect 4554 859 4706 887
rect 4554 847 4560 859
rect 4700 847 4706 859
rect 4758 887 4764 899
rect 4904 887 4910 899
rect 4758 859 4910 887
rect 4758 847 4764 859
rect 4904 847 4910 859
rect 4962 887 4968 899
rect 5108 887 5114 899
rect 4962 859 5114 887
rect 4962 847 4968 859
rect 5108 847 5114 859
rect 5166 887 5172 899
rect 5312 887 5318 899
rect 5166 859 5318 887
rect 5166 847 5172 859
rect 5312 847 5318 859
rect 5370 887 5376 899
rect 5516 887 5522 899
rect 5370 859 5522 887
rect 5370 847 5376 859
rect 5516 847 5522 859
rect 5574 887 5580 899
rect 5720 887 5726 899
rect 5574 859 5726 887
rect 5574 847 5580 859
rect 5720 847 5726 859
rect 5778 887 5784 899
rect 5924 887 5930 899
rect 5778 859 5930 887
rect 5778 847 5784 859
rect 5924 847 5930 859
rect 5982 887 5988 899
rect 6128 887 6134 899
rect 5982 859 6134 887
rect 5982 847 5988 859
rect 6128 847 6134 859
rect 6186 887 6192 899
rect 6332 887 6338 899
rect 6186 859 6338 887
rect 6186 847 6192 859
rect 6332 847 6338 859
rect 6390 887 6396 899
rect 6536 887 6542 899
rect 6390 859 6542 887
rect 6390 847 6396 859
rect 6536 847 6542 859
rect 6594 887 6600 899
rect 6740 887 6746 899
rect 6594 859 6746 887
rect 6594 847 6600 859
rect 6740 847 6746 859
rect 6798 887 6804 899
rect 6944 887 6950 899
rect 6798 859 6950 887
rect 6798 847 6804 859
rect 6944 847 6950 859
rect 7002 887 7008 899
rect 7148 887 7154 899
rect 7002 859 7154 887
rect 7002 847 7008 859
rect 7148 847 7154 859
rect 7206 887 7212 899
rect 7352 887 7358 899
rect 7206 859 7358 887
rect 7206 847 7212 859
rect 7352 847 7358 859
rect 7410 887 7416 899
rect 7556 887 7562 899
rect 7410 859 7562 887
rect 7410 847 7416 859
rect 7556 847 7562 859
rect 7614 887 7620 899
rect 7760 887 7766 899
rect 7614 859 7766 887
rect 7614 847 7620 859
rect 7760 847 7766 859
rect 7818 887 7824 899
rect 7964 887 7970 899
rect 7818 859 7970 887
rect 7818 847 7824 859
rect 7964 847 7970 859
rect 8022 887 8028 899
rect 8168 887 8174 899
rect 8022 859 8174 887
rect 8022 847 8028 859
rect 8168 847 8174 859
rect 8226 887 8232 899
rect 8372 887 8378 899
rect 8226 859 8378 887
rect 8226 847 8232 859
rect 8372 847 8378 859
rect 8430 887 8436 899
rect 8576 887 8582 899
rect 8430 859 8582 887
rect 8430 847 8436 859
rect 8576 847 8582 859
rect 8634 887 8640 899
rect 8780 887 8786 899
rect 8634 859 8786 887
rect 8634 847 8640 859
rect 8780 847 8786 859
rect 8838 887 8844 899
rect 8984 887 8990 899
rect 8838 859 8990 887
rect 8838 847 8844 859
rect 8984 847 8990 859
rect 9042 887 9048 899
rect 9188 887 9194 899
rect 9042 859 9194 887
rect 9042 847 9048 859
rect 9188 847 9194 859
rect 9246 887 9252 899
rect 9392 887 9398 899
rect 9246 859 9398 887
rect 9246 847 9252 859
rect 9392 847 9398 859
rect 9450 887 9456 899
rect 9596 887 9602 899
rect 9450 859 9602 887
rect 9450 847 9456 859
rect 9596 847 9602 859
rect 9654 887 9660 899
rect 9800 887 9806 899
rect 9654 859 9806 887
rect 9654 847 9660 859
rect 9800 847 9806 859
rect 9858 887 9864 899
rect 10004 887 10010 899
rect 9858 859 10010 887
rect 9858 847 9864 859
rect 10004 847 10010 859
rect 10062 887 10068 899
rect 10208 887 10214 899
rect 10062 859 10214 887
rect 10062 847 10068 859
rect 10208 847 10214 859
rect 10266 887 10272 899
rect 10412 887 10418 899
rect 10266 859 10418 887
rect 10266 847 10272 859
rect 10412 847 10418 859
rect 10470 887 10476 899
rect 10616 887 10622 899
rect 10470 859 10622 887
rect 10470 847 10476 859
rect 10616 847 10622 859
rect 10674 887 10680 899
rect 10820 887 10826 899
rect 10674 859 10826 887
rect 10674 847 10680 859
rect 10820 847 10826 859
rect 10878 887 10884 899
rect 11024 887 11030 899
rect 10878 859 11030 887
rect 10878 847 10884 859
rect 11024 847 11030 859
rect 11082 887 11088 899
rect 11228 887 11234 899
rect 11082 859 11234 887
rect 11082 847 11088 859
rect 11228 847 11234 859
rect 11286 887 11292 899
rect 11432 887 11438 899
rect 11286 859 11438 887
rect 11286 847 11292 859
rect 11432 847 11438 859
rect 11490 887 11496 899
rect 11636 887 11642 899
rect 11490 859 11642 887
rect 11490 847 11496 859
rect 11636 847 11642 859
rect 11694 887 11700 899
rect 11840 887 11846 899
rect 11694 859 11846 887
rect 11694 847 11700 859
rect 11840 847 11846 859
rect 11898 887 11904 899
rect 12044 887 12050 899
rect 11898 859 12050 887
rect 11898 847 11904 859
rect 12044 847 12050 859
rect 12102 887 12108 899
rect 12248 887 12254 899
rect 12102 859 12254 887
rect 12102 847 12108 859
rect 12248 847 12254 859
rect 12306 887 12312 899
rect 12452 887 12458 899
rect 12306 859 12458 887
rect 12306 847 12312 859
rect 12452 847 12458 859
rect 12510 887 12516 899
rect 12656 887 12662 899
rect 12510 859 12662 887
rect 12510 847 12516 859
rect 12656 847 12662 859
rect 12714 887 12720 899
rect 12860 887 12866 899
rect 12714 859 12866 887
rect 12714 847 12720 859
rect 12860 847 12866 859
rect 12918 887 12924 899
rect 13064 887 13070 899
rect 12918 859 13070 887
rect 12918 847 12924 859
rect 13064 847 13070 859
rect 13122 887 13128 899
rect 13268 887 13274 899
rect 13122 859 13274 887
rect 13122 847 13128 859
rect 13268 847 13274 859
rect 13326 887 13332 899
rect 13472 887 13478 899
rect 13326 859 13478 887
rect 13326 847 13332 859
rect 13472 847 13478 859
rect 13530 887 13536 899
rect 13676 887 13682 899
rect 13530 859 13682 887
rect 13530 847 13536 859
rect 13676 847 13682 859
rect 13734 887 13740 899
rect 13880 887 13886 899
rect 13734 859 13886 887
rect 13734 847 13740 859
rect 13880 847 13886 859
rect 13938 887 13944 899
rect 14084 887 14090 899
rect 13938 859 14090 887
rect 13938 847 13944 859
rect 14084 847 14090 859
rect 14142 887 14148 899
rect 14288 887 14294 899
rect 14142 859 14294 887
rect 14142 847 14148 859
rect 14288 847 14294 859
rect 14346 887 14352 899
rect 14492 887 14498 899
rect 14346 859 14498 887
rect 14346 847 14352 859
rect 14492 847 14498 859
rect 14550 887 14556 899
rect 14696 887 14702 899
rect 14550 859 14702 887
rect 14550 847 14556 859
rect 14696 847 14702 859
rect 14754 887 14760 899
rect 14900 887 14906 899
rect 14754 859 14906 887
rect 14754 847 14760 859
rect 14900 847 14906 859
rect 14958 887 14964 899
rect 15104 887 15110 899
rect 14958 859 15110 887
rect 14958 847 14964 859
rect 15104 847 15110 859
rect 15162 887 15168 899
rect 15308 887 15314 899
rect 15162 859 15314 887
rect 15162 847 15168 859
rect 15308 847 15314 859
rect 15366 887 15372 899
rect 15512 887 15518 899
rect 15366 859 15518 887
rect 15366 847 15372 859
rect 15512 847 15518 859
rect 15570 887 15576 899
rect 15716 887 15722 899
rect 15570 859 15722 887
rect 15570 847 15576 859
rect 15716 847 15722 859
rect 15774 887 15780 899
rect 15920 887 15926 899
rect 15774 859 15926 887
rect 15774 847 15780 859
rect 15920 847 15926 859
rect 15978 887 15984 899
rect 16124 887 16130 899
rect 15978 859 16130 887
rect 15978 847 15984 859
rect 16124 847 16130 859
rect 16182 887 16188 899
rect 16328 887 16334 899
rect 16182 859 16334 887
rect 16182 847 16188 859
rect 16328 847 16334 859
rect 16386 887 16392 899
rect 16532 887 16538 899
rect 16386 859 16538 887
rect 16386 847 16392 859
rect 16532 847 16538 859
rect 16590 887 16596 899
rect 16736 887 16742 899
rect 16590 859 16742 887
rect 16590 847 16596 859
rect 16736 847 16742 859
rect 16794 887 16800 899
rect 16940 887 16946 899
rect 16794 859 16946 887
rect 16794 847 16800 859
rect 16940 847 16946 859
rect 16998 887 17004 899
rect 17144 887 17150 899
rect 16998 859 17150 887
rect 16998 847 17004 859
rect 17144 847 17150 859
rect 17202 887 17208 899
rect 17348 887 17354 899
rect 17202 859 17354 887
rect 17202 847 17208 859
rect 17348 847 17354 859
rect 17406 887 17412 899
rect 17552 887 17558 899
rect 17406 859 17558 887
rect 17406 847 17412 859
rect 17552 847 17558 859
rect 17610 887 17616 899
rect 17756 887 17762 899
rect 17610 859 17762 887
rect 17610 847 17616 859
rect 17756 847 17762 859
rect 17814 887 17820 899
rect 17960 887 17966 899
rect 17814 859 17966 887
rect 17814 847 17820 859
rect 17960 847 17966 859
rect 18018 887 18024 899
rect 18164 887 18170 899
rect 18018 859 18170 887
rect 18018 847 18024 859
rect 18164 847 18170 859
rect 18222 887 18228 899
rect 18368 887 18374 899
rect 18222 859 18374 887
rect 18222 847 18228 859
rect 18368 847 18374 859
rect 18426 887 18432 899
rect 18572 887 18578 899
rect 18426 859 18578 887
rect 18426 847 18432 859
rect 18572 847 18578 859
rect 18630 887 18636 899
rect 18776 887 18782 899
rect 18630 859 18782 887
rect 18630 847 18636 859
rect 18776 847 18782 859
rect 18834 887 18840 899
rect 18980 887 18986 899
rect 18834 859 18986 887
rect 18834 847 18840 859
rect 18980 847 18986 859
rect 19038 887 19044 899
rect 19184 887 19190 899
rect 19038 859 19190 887
rect 19038 847 19044 859
rect 19184 847 19190 859
rect 19242 887 19248 899
rect 19388 887 19394 899
rect 19242 859 19394 887
rect 19242 847 19248 859
rect 19388 847 19394 859
rect 19446 887 19452 899
rect 19592 887 19598 899
rect 19446 859 19598 887
rect 19446 847 19452 859
rect 19592 847 19598 859
rect 19650 887 19656 899
rect 19796 887 19802 899
rect 19650 859 19802 887
rect 19650 847 19656 859
rect 19796 847 19802 859
rect 19854 887 19860 899
rect 20000 887 20006 899
rect 19854 859 20006 887
rect 19854 847 19860 859
rect 20000 847 20006 859
rect 20058 887 20064 899
rect 20204 887 20210 899
rect 20058 859 20210 887
rect 20058 847 20064 859
rect 20204 847 20210 859
rect 20262 887 20268 899
rect 20408 887 20414 899
rect 20262 859 20414 887
rect 20262 847 20268 859
rect 20408 847 20414 859
rect 20466 887 20472 899
rect 20612 887 20618 899
rect 20466 859 20618 887
rect 20466 847 20472 859
rect 20612 847 20618 859
rect 20670 887 20676 899
rect 20816 887 20822 899
rect 20670 859 20822 887
rect 20670 847 20676 859
rect 20816 847 20822 859
rect 20874 887 20880 899
rect 21020 887 21026 899
rect 20874 859 21026 887
rect 20874 847 20880 859
rect 21020 847 21026 859
rect 21078 887 21084 899
rect 21224 887 21230 899
rect 21078 859 21230 887
rect 21078 847 21084 859
rect 21224 847 21230 859
rect 21282 887 21288 899
rect 21428 887 21434 899
rect 21282 859 21434 887
rect 21282 847 21288 859
rect 21428 847 21434 859
rect 21486 887 21492 899
rect 21632 887 21638 899
rect 21486 859 21638 887
rect 21486 847 21492 859
rect 21632 847 21638 859
rect 21690 887 21696 899
rect 21836 887 21842 899
rect 21690 859 21842 887
rect 21690 847 21696 859
rect 21836 847 21842 859
rect 21894 887 21900 899
rect 22040 887 22046 899
rect 21894 859 22046 887
rect 21894 847 21900 859
rect 22040 847 22046 859
rect 22098 887 22104 899
rect 22244 887 22250 899
rect 22098 859 22250 887
rect 22098 847 22104 859
rect 22244 847 22250 859
rect 22302 887 22308 899
rect 22448 887 22454 899
rect 22302 859 22454 887
rect 22302 847 22308 859
rect 22448 847 22454 859
rect 22506 887 22512 899
rect 22652 887 22658 899
rect 22506 859 22658 887
rect 22506 847 22512 859
rect 22652 847 22658 859
rect 22710 887 22716 899
rect 22856 887 22862 899
rect 22710 859 22862 887
rect 22710 847 22716 859
rect 22856 847 22862 859
rect 22914 887 22920 899
rect 23060 887 23066 899
rect 22914 859 23066 887
rect 22914 847 22920 859
rect 23060 847 23066 859
rect 23118 887 23124 899
rect 23264 887 23270 899
rect 23118 859 23270 887
rect 23118 847 23124 859
rect 23264 847 23270 859
rect 23322 887 23328 899
rect 23468 887 23474 899
rect 23322 859 23474 887
rect 23322 847 23328 859
rect 23468 847 23474 859
rect 23526 887 23532 899
rect 23672 887 23678 899
rect 23526 859 23678 887
rect 23526 847 23532 859
rect 23672 847 23678 859
rect 23730 887 23736 899
rect 23876 887 23882 899
rect 23730 859 23882 887
rect 23730 847 23736 859
rect 23876 847 23882 859
rect 23934 887 23940 899
rect 24080 887 24086 899
rect 23934 859 24086 887
rect 23934 847 23940 859
rect 24080 847 24086 859
rect 24138 887 24144 899
rect 24284 887 24290 899
rect 24138 859 24290 887
rect 24138 847 24144 859
rect 24284 847 24290 859
rect 24342 887 24348 899
rect 24488 887 24494 899
rect 24342 859 24494 887
rect 24342 847 24348 859
rect 24488 847 24494 859
rect 24546 887 24552 899
rect 24692 887 24698 899
rect 24546 859 24698 887
rect 24546 847 24552 859
rect 24692 847 24698 859
rect 24750 887 24756 899
rect 24896 887 24902 899
rect 24750 859 24902 887
rect 24750 847 24756 859
rect 24896 847 24902 859
rect 24954 887 24960 899
rect 25100 887 25106 899
rect 24954 859 25106 887
rect 24954 847 24960 859
rect 25100 847 25106 859
rect 25158 887 25164 899
rect 25304 887 25310 899
rect 25158 859 25310 887
rect 25158 847 25164 859
rect 25304 847 25310 859
rect 25362 887 25368 899
rect 25508 887 25514 899
rect 25362 859 25514 887
rect 25362 847 25368 859
rect 25508 847 25514 859
rect 25566 887 25572 899
rect 25712 887 25718 899
rect 25566 859 25718 887
rect 25566 847 25572 859
rect 25712 847 25718 859
rect 25770 887 25776 899
rect 25916 887 25922 899
rect 25770 859 25922 887
rect 25770 847 25776 859
rect 25916 847 25922 859
rect 25974 887 25980 899
rect 26120 887 26126 899
rect 25974 859 26126 887
rect 25974 847 25980 859
rect 26120 847 26126 859
rect 26178 887 26184 899
rect 26324 887 26330 899
rect 26178 859 26330 887
rect 26178 847 26184 859
rect 26324 847 26330 859
rect 26382 887 26388 899
rect 26528 887 26534 899
rect 26382 859 26534 887
rect 26382 847 26388 859
rect 26528 847 26534 859
rect 26586 887 26592 899
rect 26732 887 26738 899
rect 26586 859 26738 887
rect 26586 847 26592 859
rect 26732 847 26738 859
rect 26790 887 26796 899
rect 26936 887 26942 899
rect 26790 859 26942 887
rect 26790 847 26796 859
rect 26936 847 26942 859
rect 26994 887 27000 899
rect 27140 887 27146 899
rect 26994 859 27146 887
rect 26994 847 27000 859
rect 27140 847 27146 859
rect 27198 887 27204 899
rect 27344 887 27350 899
rect 27198 859 27350 887
rect 27198 847 27204 859
rect 27344 847 27350 859
rect 27402 887 27408 899
rect 27548 887 27554 899
rect 27402 859 27554 887
rect 27402 847 27408 859
rect 27548 847 27554 859
rect 27606 887 27612 899
rect 27752 887 27758 899
rect 27606 859 27758 887
rect 27606 847 27612 859
rect 27752 847 27758 859
rect 27810 887 27816 899
rect 27956 887 27962 899
rect 27810 859 27962 887
rect 27810 847 27816 859
rect 27956 847 27962 859
rect 28014 887 28020 899
rect 28160 887 28166 899
rect 28014 859 28166 887
rect 28014 847 28020 859
rect 28160 847 28166 859
rect 28218 887 28224 899
rect 28364 887 28370 899
rect 28218 859 28370 887
rect 28218 847 28224 859
rect 28364 847 28370 859
rect 28422 887 28428 899
rect 28568 887 28574 899
rect 28422 859 28574 887
rect 28422 847 28428 859
rect 28568 847 28574 859
rect 28626 887 28632 899
rect 28772 887 28778 899
rect 28626 859 28778 887
rect 28626 847 28632 859
rect 28772 847 28778 859
rect 28830 887 28836 899
rect 28976 887 28982 899
rect 28830 859 28982 887
rect 28830 847 28836 859
rect 28976 847 28982 859
rect 29034 887 29040 899
rect 29180 887 29186 899
rect 29034 859 29186 887
rect 29034 847 29040 859
rect 29180 847 29186 859
rect 29238 887 29244 899
rect 29384 887 29390 899
rect 29238 859 29390 887
rect 29238 847 29244 859
rect 29384 847 29390 859
rect 29442 887 29448 899
rect 29588 887 29594 899
rect 29442 859 29594 887
rect 29442 847 29448 859
rect 29588 847 29594 859
rect 29646 887 29652 899
rect 29792 887 29798 899
rect 29646 859 29798 887
rect 29646 847 29652 859
rect 29792 847 29798 859
rect 29850 887 29856 899
rect 29996 887 30002 899
rect 29850 859 30002 887
rect 29850 847 29856 859
rect 29996 847 30002 859
rect 30054 887 30060 899
rect 30200 887 30206 899
rect 30054 859 30206 887
rect 30054 847 30060 859
rect 30200 847 30206 859
rect 30258 887 30264 899
rect 30404 887 30410 899
rect 30258 859 30410 887
rect 30258 847 30264 859
rect 30404 847 30410 859
rect 30462 887 30468 899
rect 30608 887 30614 899
rect 30462 859 30614 887
rect 30462 847 30468 859
rect 30608 847 30614 859
rect 30666 887 30672 899
rect 30812 887 30818 899
rect 30666 859 30818 887
rect 30666 847 30672 859
rect 30812 847 30818 859
rect 30870 887 30876 899
rect 31016 887 31022 899
rect 30870 859 31022 887
rect 30870 847 30876 859
rect 31016 847 31022 859
rect 31074 887 31080 899
rect 31220 887 31226 899
rect 31074 859 31226 887
rect 31074 847 31080 859
rect 31220 847 31226 859
rect 31278 887 31284 899
rect 31424 887 31430 899
rect 31278 859 31430 887
rect 31278 847 31284 859
rect 31424 847 31430 859
rect 31482 887 31488 899
rect 31628 887 31634 899
rect 31482 859 31634 887
rect 31482 847 31488 859
rect 31628 847 31634 859
rect 31686 887 31692 899
rect 31832 887 31838 899
rect 31686 859 31838 887
rect 31686 847 31692 859
rect 31832 847 31838 859
rect 31890 887 31896 899
rect 32036 887 32042 899
rect 31890 859 32042 887
rect 31890 847 31896 859
rect 32036 847 32042 859
rect 32094 887 32100 899
rect 32240 887 32246 899
rect 32094 859 32246 887
rect 32094 847 32100 859
rect 32240 847 32246 859
rect 32298 887 32304 899
rect 32444 887 32450 899
rect 32298 859 32450 887
rect 32298 847 32304 859
rect 32444 847 32450 859
rect 32502 887 32508 899
rect 32648 887 32654 899
rect 32502 859 32654 887
rect 32502 847 32508 859
rect 32648 847 32654 859
rect 32706 887 32712 899
rect 32852 887 32858 899
rect 32706 859 32858 887
rect 32706 847 32712 859
rect 32852 847 32858 859
rect 32910 887 32916 899
rect 33056 887 33062 899
rect 32910 859 33062 887
rect 32910 847 32916 859
rect 33056 847 33062 859
rect 33114 887 33120 899
rect 33260 887 33266 899
rect 33114 859 33266 887
rect 33114 847 33120 859
rect 33260 847 33266 859
rect 33318 887 33324 899
rect 33464 887 33470 899
rect 33318 859 33470 887
rect 33318 847 33324 859
rect 33464 847 33470 859
rect 33522 887 33528 899
rect 33668 887 33674 899
rect 33522 859 33674 887
rect 33522 847 33528 859
rect 33668 847 33674 859
rect 33726 887 33732 899
rect 33872 887 33878 899
rect 33726 859 33878 887
rect 33726 847 33732 859
rect 33872 847 33878 859
rect 33930 887 33936 899
rect 34076 887 34082 899
rect 33930 859 34082 887
rect 33930 847 33936 859
rect 34076 847 34082 859
rect 34134 887 34140 899
rect 34280 887 34286 899
rect 34134 859 34286 887
rect 34134 847 34140 859
rect 34280 847 34286 859
rect 34338 887 34344 899
rect 34484 887 34490 899
rect 34338 859 34490 887
rect 34338 847 34344 859
rect 34484 847 34490 859
rect 34542 887 34548 899
rect 34688 887 34694 899
rect 34542 859 34694 887
rect 34542 847 34548 859
rect 34688 847 34694 859
rect 34746 887 34752 899
rect 34892 887 34898 899
rect 34746 859 34898 887
rect 34746 847 34752 859
rect 34892 847 34898 859
rect 34950 887 34956 899
rect 35096 887 35102 899
rect 34950 859 35102 887
rect 34950 847 34956 859
rect 35096 847 35102 859
rect 35154 887 35160 899
rect 35300 887 35306 899
rect 35154 859 35306 887
rect 35154 847 35160 859
rect 35300 847 35306 859
rect 35358 887 35364 899
rect 35504 887 35510 899
rect 35358 859 35510 887
rect 35358 847 35364 859
rect 35504 847 35510 859
rect 35562 887 35568 899
rect 35708 887 35714 899
rect 35562 859 35714 887
rect 35562 847 35568 859
rect 35708 847 35714 859
rect 35766 887 35772 899
rect 35912 887 35918 899
rect 35766 859 35918 887
rect 35766 847 35772 859
rect 35912 847 35918 859
rect 35970 887 35976 899
rect 36116 887 36122 899
rect 35970 859 36122 887
rect 35970 847 35976 859
rect 36116 847 36122 859
rect 36174 887 36180 899
rect 36320 887 36326 899
rect 36174 859 36326 887
rect 36174 847 36180 859
rect 36320 847 36326 859
rect 36378 887 36384 899
rect 36524 887 36530 899
rect 36378 859 36530 887
rect 36378 847 36384 859
rect 36524 847 36530 859
rect 36582 887 36588 899
rect 36728 887 36734 899
rect 36582 859 36734 887
rect 36582 847 36588 859
rect 36728 847 36734 859
rect 36786 887 36792 899
rect 36932 887 36938 899
rect 36786 859 36938 887
rect 36786 847 36792 859
rect 36932 847 36938 859
rect 36990 887 36996 899
rect 37136 887 37142 899
rect 36990 859 37142 887
rect 36990 847 36996 859
rect 37136 847 37142 859
rect 37194 887 37200 899
rect 37340 887 37346 899
rect 37194 859 37346 887
rect 37194 847 37200 859
rect 37340 847 37346 859
rect 37398 887 37404 899
rect 37544 887 37550 899
rect 37398 859 37550 887
rect 37398 847 37404 859
rect 37544 847 37550 859
rect 37602 887 37608 899
rect 37748 887 37754 899
rect 37602 859 37754 887
rect 37602 847 37608 859
rect 37748 847 37754 859
rect 37806 887 37812 899
rect 37952 887 37958 899
rect 37806 859 37958 887
rect 37806 847 37812 859
rect 37952 847 37958 859
rect 38010 887 38016 899
rect 38156 887 38162 899
rect 38010 859 38162 887
rect 38010 847 38016 859
rect 38156 847 38162 859
rect 38214 887 38220 899
rect 38360 887 38366 899
rect 38214 859 38366 887
rect 38214 847 38220 859
rect 38360 847 38366 859
rect 38418 887 38424 899
rect 38564 887 38570 899
rect 38418 859 38570 887
rect 38418 847 38424 859
rect 38564 847 38570 859
rect 38622 887 38628 899
rect 38768 887 38774 899
rect 38622 859 38774 887
rect 38622 847 38628 859
rect 38768 847 38774 859
rect 38826 887 38832 899
rect 38972 887 38978 899
rect 38826 859 38978 887
rect 38826 847 38832 859
rect 38972 847 38978 859
rect 39030 887 39036 899
rect 39176 887 39182 899
rect 39030 859 39182 887
rect 39030 847 39036 859
rect 39176 847 39182 859
rect 39234 887 39240 899
rect 39380 887 39386 899
rect 39234 859 39386 887
rect 39234 847 39240 859
rect 39380 847 39386 859
rect 39438 887 39444 899
rect 39584 887 39590 899
rect 39438 859 39590 887
rect 39438 847 39444 859
rect 39584 847 39590 859
rect 39642 887 39648 899
rect 39788 887 39794 899
rect 39642 859 39794 887
rect 39642 847 39648 859
rect 39788 847 39794 859
rect 39846 887 39852 899
rect 39992 887 39998 899
rect 39846 859 39998 887
rect 39846 847 39852 859
rect 39992 847 39998 859
rect 40050 887 40056 899
rect 40196 887 40202 899
rect 40050 859 40202 887
rect 40050 847 40056 859
rect 40196 847 40202 859
rect 40254 887 40260 899
rect 40400 887 40406 899
rect 40254 859 40406 887
rect 40254 847 40260 859
rect 40400 847 40406 859
rect 40458 887 40464 899
rect 40604 887 40610 899
rect 40458 859 40610 887
rect 40458 847 40464 859
rect 40604 847 40610 859
rect 40662 887 40668 899
rect 40808 887 40814 899
rect 40662 859 40814 887
rect 40662 847 40668 859
rect 40808 847 40814 859
rect 40866 887 40872 899
rect 41012 887 41018 899
rect 40866 859 41018 887
rect 40866 847 40872 859
rect 41012 847 41018 859
rect 41070 887 41076 899
rect 41216 887 41222 899
rect 41070 859 41222 887
rect 41070 847 41076 859
rect 41216 847 41222 859
rect 41274 887 41280 899
rect 41420 887 41426 899
rect 41274 859 41426 887
rect 41274 847 41280 859
rect 41420 847 41426 859
rect 41478 887 41484 899
rect 41624 887 41630 899
rect 41478 859 41630 887
rect 41478 847 41484 859
rect 41624 847 41630 859
rect 41682 887 41688 899
rect 41828 887 41834 899
rect 41682 859 41834 887
rect 41682 847 41688 859
rect 41828 847 41834 859
rect 41886 887 41892 899
rect 42032 887 42038 899
rect 41886 859 42038 887
rect 41886 847 41892 859
rect 42032 847 42038 859
rect 42090 887 42096 899
rect 42236 887 42242 899
rect 42090 859 42242 887
rect 42090 847 42096 859
rect 42236 847 42242 859
rect 42294 887 42300 899
rect 42440 887 42446 899
rect 42294 859 42446 887
rect 42294 847 42300 859
rect 42440 847 42446 859
rect 42498 887 42504 899
rect 42644 887 42650 899
rect 42498 859 42650 887
rect 42498 847 42504 859
rect 42644 847 42650 859
rect 42702 887 42708 899
rect 42848 887 42854 899
rect 42702 859 42854 887
rect 42702 847 42708 859
rect 42848 847 42854 859
rect 42906 887 42912 899
rect 43052 887 43058 899
rect 42906 859 43058 887
rect 42906 847 42912 859
rect 43052 847 43058 859
rect 43110 887 43116 899
rect 43256 887 43262 899
rect 43110 859 43262 887
rect 43110 847 43116 859
rect 43256 847 43262 859
rect 43314 887 43320 899
rect 43460 887 43466 899
rect 43314 859 43466 887
rect 43314 847 43320 859
rect 43460 847 43466 859
rect 43518 887 43524 899
rect 43664 887 43670 899
rect 43518 859 43670 887
rect 43518 847 43524 859
rect 43664 847 43670 859
rect 43722 887 43728 899
rect 43868 887 43874 899
rect 43722 859 43874 887
rect 43722 847 43728 859
rect 43868 847 43874 859
rect 43926 887 43932 899
rect 44072 887 44078 899
rect 43926 859 44078 887
rect 43926 847 43932 859
rect 44072 847 44078 859
rect 44130 887 44136 899
rect 44276 887 44282 899
rect 44130 859 44282 887
rect 44130 847 44136 859
rect 44276 847 44282 859
rect 44334 887 44340 899
rect 44480 887 44486 899
rect 44334 859 44486 887
rect 44334 847 44340 859
rect 44480 847 44486 859
rect 44538 887 44544 899
rect 44684 887 44690 899
rect 44538 859 44690 887
rect 44538 847 44544 859
rect 44684 847 44690 859
rect 44742 887 44748 899
rect 44888 887 44894 899
rect 44742 859 44894 887
rect 44742 847 44748 859
rect 44888 847 44894 859
rect 44946 887 44952 899
rect 45092 887 45098 899
rect 44946 859 45098 887
rect 44946 847 44952 859
rect 45092 847 45098 859
rect 45150 887 45156 899
rect 45296 887 45302 899
rect 45150 859 45302 887
rect 45150 847 45156 859
rect 45296 847 45302 859
rect 45354 887 45360 899
rect 45500 887 45506 899
rect 45354 859 45506 887
rect 45354 847 45360 859
rect 45500 847 45506 859
rect 45558 887 45564 899
rect 45704 887 45710 899
rect 45558 859 45710 887
rect 45558 847 45564 859
rect 45704 847 45710 859
rect 45762 887 45768 899
rect 45908 887 45914 899
rect 45762 859 45914 887
rect 45762 847 45768 859
rect 45908 847 45914 859
rect 45966 887 45972 899
rect 46112 887 46118 899
rect 45966 859 46118 887
rect 45966 847 45972 859
rect 46112 847 46118 859
rect 46170 887 46176 899
rect 46316 887 46322 899
rect 46170 859 46322 887
rect 46170 847 46176 859
rect 46316 847 46322 859
rect 46374 887 46380 899
rect 46520 887 46526 899
rect 46374 859 46526 887
rect 46374 847 46380 859
rect 46520 847 46526 859
rect 46578 887 46584 899
rect 46724 887 46730 899
rect 46578 859 46730 887
rect 46578 847 46584 859
rect 46724 847 46730 859
rect 46782 887 46788 899
rect 46928 887 46934 899
rect 46782 859 46934 887
rect 46782 847 46788 859
rect 46928 847 46934 859
rect 46986 887 46992 899
rect 47132 887 47138 899
rect 46986 859 47138 887
rect 46986 847 46992 859
rect 47132 847 47138 859
rect 47190 887 47196 899
rect 47336 887 47342 899
rect 47190 859 47342 887
rect 47190 847 47196 859
rect 47336 847 47342 859
rect 47394 887 47400 899
rect 47540 887 47546 899
rect 47394 859 47546 887
rect 47394 847 47400 859
rect 47540 847 47546 859
rect 47598 887 47604 899
rect 47744 887 47750 899
rect 47598 859 47750 887
rect 47598 847 47604 859
rect 47744 847 47750 859
rect 47802 887 47808 899
rect 47948 887 47954 899
rect 47802 859 47954 887
rect 47802 847 47808 859
rect 47948 847 47954 859
rect 48006 887 48012 899
rect 48152 887 48158 899
rect 48006 859 48158 887
rect 48006 847 48012 859
rect 48152 847 48158 859
rect 48210 887 48216 899
rect 48356 887 48362 899
rect 48210 859 48362 887
rect 48210 847 48216 859
rect 48356 847 48362 859
rect 48414 887 48420 899
rect 48560 887 48566 899
rect 48414 859 48566 887
rect 48414 847 48420 859
rect 48560 847 48566 859
rect 48618 887 48624 899
rect 48764 887 48770 899
rect 48618 859 48770 887
rect 48618 847 48624 859
rect 48764 847 48770 859
rect 48822 887 48828 899
rect 48968 887 48974 899
rect 48822 859 48974 887
rect 48822 847 48828 859
rect 48968 847 48974 859
rect 49026 887 49032 899
rect 49172 887 49178 899
rect 49026 859 49178 887
rect 49026 847 49032 859
rect 49172 847 49178 859
rect 49230 887 49236 899
rect 49376 887 49382 899
rect 49230 859 49382 887
rect 49230 847 49236 859
rect 49376 847 49382 859
rect 49434 887 49440 899
rect 49580 887 49586 899
rect 49434 859 49586 887
rect 49434 847 49440 859
rect 49580 847 49586 859
rect 49638 887 49644 899
rect 49784 887 49790 899
rect 49638 859 49790 887
rect 49638 847 49644 859
rect 49784 847 49790 859
rect 49842 887 49848 899
rect 49988 887 49994 899
rect 49842 859 49994 887
rect 49842 847 49848 859
rect 49988 847 49994 859
rect 50046 887 50052 899
rect 50192 887 50198 899
rect 50046 859 50198 887
rect 50046 847 50052 859
rect 50192 847 50198 859
rect 50250 887 50256 899
rect 50396 887 50402 899
rect 50250 859 50402 887
rect 50250 847 50256 859
rect 50396 847 50402 859
rect 50454 887 50460 899
rect 50600 887 50606 899
rect 50454 859 50606 887
rect 50454 847 50460 859
rect 50600 847 50606 859
rect 50658 887 50664 899
rect 50804 887 50810 899
rect 50658 859 50810 887
rect 50658 847 50664 859
rect 50804 847 50810 859
rect 50862 887 50868 899
rect 51008 887 51014 899
rect 50862 859 51014 887
rect 50862 847 50868 859
rect 51008 847 51014 859
rect 51066 887 51072 899
rect 51212 887 51218 899
rect 51066 859 51218 887
rect 51066 847 51072 859
rect 51212 847 51218 859
rect 51270 887 51276 899
rect 51416 887 51422 899
rect 51270 859 51422 887
rect 51270 847 51276 859
rect 51416 847 51422 859
rect 51474 887 51480 899
rect 51620 887 51626 899
rect 51474 859 51626 887
rect 51474 847 51480 859
rect 51620 847 51626 859
rect 51678 887 51684 899
rect 51824 887 51830 899
rect 51678 859 51830 887
rect 51678 847 51684 859
rect 51824 847 51830 859
rect 51882 887 51888 899
rect 52028 887 52034 899
rect 51882 859 52034 887
rect 51882 847 51888 859
rect 52028 847 52034 859
rect 52086 887 52092 899
rect 52246 887 52252 899
rect 52086 859 52252 887
rect 52086 847 52092 859
rect 52246 847 52252 859
rect 52304 847 52310 899
rect 61 368 89 396
rect 12 -32 40 32
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_0
timestamp 1581449086
transform 1 0 52020 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1
timestamp 1581449086
transform 1 0 51816 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_2
timestamp 1581449086
transform 1 0 51612 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_3
timestamp 1581449086
transform 1 0 51408 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_4
timestamp 1581449086
transform 1 0 51204 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_5
timestamp 1581449086
transform 1 0 51000 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_6
timestamp 1581449086
transform 1 0 50796 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_7
timestamp 1581449086
transform 1 0 50592 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_8
timestamp 1581449086
transform 1 0 50388 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_9
timestamp 1581449086
transform 1 0 50184 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_10
timestamp 1581449086
transform 1 0 49980 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_11
timestamp 1581449086
transform 1 0 49776 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_12
timestamp 1581449086
transform 1 0 49572 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_13
timestamp 1581449086
transform 1 0 49368 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_14
timestamp 1581449086
transform 1 0 49164 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_15
timestamp 1581449086
transform 1 0 48960 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_16
timestamp 1581449086
transform 1 0 48756 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_17
timestamp 1581449086
transform 1 0 48552 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_18
timestamp 1581449086
transform 1 0 48348 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_19
timestamp 1581449086
transform 1 0 48144 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_20
timestamp 1581449086
transform 1 0 47940 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_21
timestamp 1581449086
transform 1 0 47736 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_22
timestamp 1581449086
transform 1 0 47532 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_23
timestamp 1581449086
transform 1 0 47328 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_24
timestamp 1581449086
transform 1 0 47124 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_25
timestamp 1581449086
transform 1 0 46920 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_26
timestamp 1581449086
transform 1 0 46716 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_27
timestamp 1581449086
transform 1 0 46512 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_28
timestamp 1581449086
transform 1 0 46308 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_29
timestamp 1581449086
transform 1 0 46104 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_30
timestamp 1581449086
transform 1 0 45900 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_31
timestamp 1581449086
transform 1 0 45696 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_32
timestamp 1581449086
transform 1 0 45492 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_33
timestamp 1581449086
transform 1 0 45288 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_34
timestamp 1581449086
transform 1 0 45084 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_35
timestamp 1581449086
transform 1 0 44880 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_36
timestamp 1581449086
transform 1 0 44676 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_37
timestamp 1581449086
transform 1 0 44472 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_38
timestamp 1581449086
transform 1 0 44268 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_39
timestamp 1581449086
transform 1 0 44064 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_40
timestamp 1581449086
transform 1 0 43860 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_41
timestamp 1581449086
transform 1 0 43656 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_42
timestamp 1581449086
transform 1 0 43452 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_43
timestamp 1581449086
transform 1 0 43248 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_44
timestamp 1581449086
transform 1 0 43044 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_45
timestamp 1581449086
transform 1 0 42840 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_46
timestamp 1581449086
transform 1 0 42636 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_47
timestamp 1581449086
transform 1 0 42432 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_48
timestamp 1581449086
transform 1 0 42228 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_49
timestamp 1581449086
transform 1 0 42024 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_50
timestamp 1581449086
transform 1 0 41820 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_51
timestamp 1581449086
transform 1 0 41616 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_52
timestamp 1581449086
transform 1 0 41412 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_53
timestamp 1581449086
transform 1 0 41208 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_54
timestamp 1581449086
transform 1 0 41004 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_55
timestamp 1581449086
transform 1 0 40800 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_56
timestamp 1581449086
transform 1 0 40596 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_57
timestamp 1581449086
transform 1 0 40392 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_58
timestamp 1581449086
transform 1 0 40188 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_59
timestamp 1581449086
transform 1 0 39984 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_60
timestamp 1581449086
transform 1 0 39780 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_61
timestamp 1581449086
transform 1 0 39576 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_62
timestamp 1581449086
transform 1 0 39372 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_63
timestamp 1581449086
transform 1 0 39168 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_64
timestamp 1581449086
transform 1 0 38964 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_65
timestamp 1581449086
transform 1 0 38760 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_66
timestamp 1581449086
transform 1 0 38556 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_67
timestamp 1581449086
transform 1 0 38352 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_68
timestamp 1581449086
transform 1 0 38148 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_69
timestamp 1581449086
transform 1 0 37944 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_70
timestamp 1581449086
transform 1 0 37740 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_71
timestamp 1581449086
transform 1 0 37536 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_72
timestamp 1581449086
transform 1 0 37332 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_73
timestamp 1581449086
transform 1 0 37128 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_74
timestamp 1581449086
transform 1 0 36924 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_75
timestamp 1581449086
transform 1 0 36720 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_76
timestamp 1581449086
transform 1 0 36516 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_77
timestamp 1581449086
transform 1 0 36312 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_78
timestamp 1581449086
transform 1 0 36108 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_79
timestamp 1581449086
transform 1 0 35904 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_80
timestamp 1581449086
transform 1 0 35700 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_81
timestamp 1581449086
transform 1 0 35496 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_82
timestamp 1581449086
transform 1 0 35292 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_83
timestamp 1581449086
transform 1 0 35088 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_84
timestamp 1581449086
transform 1 0 34884 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_85
timestamp 1581449086
transform 1 0 34680 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_86
timestamp 1581449086
transform 1 0 34476 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_87
timestamp 1581449086
transform 1 0 34272 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_88
timestamp 1581449086
transform 1 0 34068 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_89
timestamp 1581449086
transform 1 0 33864 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_90
timestamp 1581449086
transform 1 0 33660 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_91
timestamp 1581449086
transform 1 0 33456 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_92
timestamp 1581449086
transform 1 0 33252 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_93
timestamp 1581449086
transform 1 0 33048 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_94
timestamp 1581449086
transform 1 0 32844 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_95
timestamp 1581449086
transform 1 0 32640 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_96
timestamp 1581449086
transform 1 0 32436 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_97
timestamp 1581449086
transform 1 0 32232 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_98
timestamp 1581449086
transform 1 0 32028 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_99
timestamp 1581449086
transform 1 0 31824 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_100
timestamp 1581449086
transform 1 0 31620 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_101
timestamp 1581449086
transform 1 0 31416 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_102
timestamp 1581449086
transform 1 0 31212 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_103
timestamp 1581449086
transform 1 0 31008 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_104
timestamp 1581449086
transform 1 0 30804 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_105
timestamp 1581449086
transform 1 0 30600 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_106
timestamp 1581449086
transform 1 0 30396 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_107
timestamp 1581449086
transform 1 0 30192 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_108
timestamp 1581449086
transform 1 0 29988 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_109
timestamp 1581449086
transform 1 0 29784 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_110
timestamp 1581449086
transform 1 0 29580 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_111
timestamp 1581449086
transform 1 0 29376 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_112
timestamp 1581449086
transform 1 0 29172 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_113
timestamp 1581449086
transform 1 0 28968 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_114
timestamp 1581449086
transform 1 0 28764 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_115
timestamp 1581449086
transform 1 0 28560 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_116
timestamp 1581449086
transform 1 0 28356 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_117
timestamp 1581449086
transform 1 0 28152 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_118
timestamp 1581449086
transform 1 0 27948 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_119
timestamp 1581449086
transform 1 0 27744 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_120
timestamp 1581449086
transform 1 0 27540 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_121
timestamp 1581449086
transform 1 0 27336 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_122
timestamp 1581449086
transform 1 0 27132 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_123
timestamp 1581449086
transform 1 0 26928 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_124
timestamp 1581449086
transform 1 0 26724 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_125
timestamp 1581449086
transform 1 0 26520 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_126
timestamp 1581449086
transform 1 0 26316 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_127
timestamp 1581449086
transform 1 0 26112 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_128
timestamp 1581449086
transform 1 0 25908 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_129
timestamp 1581449086
transform 1 0 25704 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_130
timestamp 1581449086
transform 1 0 25500 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_131
timestamp 1581449086
transform 1 0 25296 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_132
timestamp 1581449086
transform 1 0 25092 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_133
timestamp 1581449086
transform 1 0 24888 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_134
timestamp 1581449086
transform 1 0 24684 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_135
timestamp 1581449086
transform 1 0 24480 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_136
timestamp 1581449086
transform 1 0 24276 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_137
timestamp 1581449086
transform 1 0 24072 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_138
timestamp 1581449086
transform 1 0 23868 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_139
timestamp 1581449086
transform 1 0 23664 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_140
timestamp 1581449086
transform 1 0 23460 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_141
timestamp 1581449086
transform 1 0 23256 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_142
timestamp 1581449086
transform 1 0 23052 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_143
timestamp 1581449086
transform 1 0 22848 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_144
timestamp 1581449086
transform 1 0 22644 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_145
timestamp 1581449086
transform 1 0 22440 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_146
timestamp 1581449086
transform 1 0 22236 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_147
timestamp 1581449086
transform 1 0 22032 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_148
timestamp 1581449086
transform 1 0 21828 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_149
timestamp 1581449086
transform 1 0 21624 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_150
timestamp 1581449086
transform 1 0 21420 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_151
timestamp 1581449086
transform 1 0 21216 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_152
timestamp 1581449086
transform 1 0 21012 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_153
timestamp 1581449086
transform 1 0 20808 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_154
timestamp 1581449086
transform 1 0 20604 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_155
timestamp 1581449086
transform 1 0 20400 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_156
timestamp 1581449086
transform 1 0 20196 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_157
timestamp 1581449086
transform 1 0 19992 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_158
timestamp 1581449086
transform 1 0 19788 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_159
timestamp 1581449086
transform 1 0 19584 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_160
timestamp 1581449086
transform 1 0 19380 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_161
timestamp 1581449086
transform 1 0 19176 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_162
timestamp 1581449086
transform 1 0 18972 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_163
timestamp 1581449086
transform 1 0 18768 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_164
timestamp 1581449086
transform 1 0 18564 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_165
timestamp 1581449086
transform 1 0 18360 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_166
timestamp 1581449086
transform 1 0 18156 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_167
timestamp 1581449086
transform 1 0 17952 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_168
timestamp 1581449086
transform 1 0 17748 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_169
timestamp 1581449086
transform 1 0 17544 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_170
timestamp 1581449086
transform 1 0 17340 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_171
timestamp 1581449086
transform 1 0 17136 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_172
timestamp 1581449086
transform 1 0 16932 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_173
timestamp 1581449086
transform 1 0 16728 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_174
timestamp 1581449086
transform 1 0 16524 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_175
timestamp 1581449086
transform 1 0 16320 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_176
timestamp 1581449086
transform 1 0 16116 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_177
timestamp 1581449086
transform 1 0 15912 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_178
timestamp 1581449086
transform 1 0 15708 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_179
timestamp 1581449086
transform 1 0 15504 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_180
timestamp 1581449086
transform 1 0 15300 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_181
timestamp 1581449086
transform 1 0 15096 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_182
timestamp 1581449086
transform 1 0 14892 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_183
timestamp 1581449086
transform 1 0 14688 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_184
timestamp 1581449086
transform 1 0 14484 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_185
timestamp 1581449086
transform 1 0 14280 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_186
timestamp 1581449086
transform 1 0 14076 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_187
timestamp 1581449086
transform 1 0 13872 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_188
timestamp 1581449086
transform 1 0 13668 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_189
timestamp 1581449086
transform 1 0 13464 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_190
timestamp 1581449086
transform 1 0 13260 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_191
timestamp 1581449086
transform 1 0 13056 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_192
timestamp 1581449086
transform 1 0 12852 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_193
timestamp 1581449086
transform 1 0 12648 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_194
timestamp 1581449086
transform 1 0 12444 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_195
timestamp 1581449086
transform 1 0 12240 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_196
timestamp 1581449086
transform 1 0 12036 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_197
timestamp 1581449086
transform 1 0 11832 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_198
timestamp 1581449086
transform 1 0 11628 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_199
timestamp 1581449086
transform 1 0 11424 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_200
timestamp 1581449086
transform 1 0 11220 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_201
timestamp 1581449086
transform 1 0 11016 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_202
timestamp 1581449086
transform 1 0 10812 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_203
timestamp 1581449086
transform 1 0 10608 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_204
timestamp 1581449086
transform 1 0 10404 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_205
timestamp 1581449086
transform 1 0 10200 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_206
timestamp 1581449086
transform 1 0 9996 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_207
timestamp 1581449086
transform 1 0 9792 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_208
timestamp 1581449086
transform 1 0 9588 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_209
timestamp 1581449086
transform 1 0 9384 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_210
timestamp 1581449086
transform 1 0 9180 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_211
timestamp 1581449086
transform 1 0 8976 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_212
timestamp 1581449086
transform 1 0 8772 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_213
timestamp 1581449086
transform 1 0 8568 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_214
timestamp 1581449086
transform 1 0 8364 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_215
timestamp 1581449086
transform 1 0 8160 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_216
timestamp 1581449086
transform 1 0 7956 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_217
timestamp 1581449086
transform 1 0 7752 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_218
timestamp 1581449086
transform 1 0 7548 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_219
timestamp 1581449086
transform 1 0 7344 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_220
timestamp 1581449086
transform 1 0 7140 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_221
timestamp 1581449086
transform 1 0 6936 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_222
timestamp 1581449086
transform 1 0 6732 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_223
timestamp 1581449086
transform 1 0 6528 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_224
timestamp 1581449086
transform 1 0 6324 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_225
timestamp 1581449086
transform 1 0 6120 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_226
timestamp 1581449086
transform 1 0 5916 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_227
timestamp 1581449086
transform 1 0 5712 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_228
timestamp 1581449086
transform 1 0 5508 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_229
timestamp 1581449086
transform 1 0 5304 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_230
timestamp 1581449086
transform 1 0 5100 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_231
timestamp 1581449086
transform 1 0 4896 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_232
timestamp 1581449086
transform 1 0 4692 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_233
timestamp 1581449086
transform 1 0 4488 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_234
timestamp 1581449086
transform 1 0 4284 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_235
timestamp 1581449086
transform 1 0 4080 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_236
timestamp 1581449086
transform 1 0 3876 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_237
timestamp 1581449086
transform 1 0 3672 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_238
timestamp 1581449086
transform 1 0 3468 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_239
timestamp 1581449086
transform 1 0 3264 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_240
timestamp 1581449086
transform 1 0 3060 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_241
timestamp 1581449086
transform 1 0 2856 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_242
timestamp 1581449086
transform 1 0 2652 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_243
timestamp 1581449086
transform 1 0 2448 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_244
timestamp 1581449086
transform 1 0 2244 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_245
timestamp 1581449086
transform 1 0 2040 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_246
timestamp 1581449086
transform 1 0 1836 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_247
timestamp 1581449086
transform 1 0 1632 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_248
timestamp 1581449086
transform 1 0 1428 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_249
timestamp 1581449086
transform 1 0 1224 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_250
timestamp 1581449086
transform 1 0 1020 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_251
timestamp 1581449086
transform 1 0 816 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_252
timestamp 1581449086
transform 1 0 612 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_253
timestamp 1581449086
transform 1 0 408 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_254
timestamp 1581449086
transform 1 0 204 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_255
timestamp 1581449086
transform 1 0 0 0 1 2609
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_256
timestamp 1581449086
transform 1 0 51816 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_257
timestamp 1581449086
transform 1 0 51612 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_258
timestamp 1581449086
transform 1 0 50796 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_259
timestamp 1581449086
transform 1 0 50388 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_260
timestamp 1581449086
transform 1 0 50184 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_261
timestamp 1581449086
transform 1 0 49980 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_262
timestamp 1581449086
transform 1 0 49776 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_263
timestamp 1581449086
transform 1 0 49164 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_264
timestamp 1581449086
transform 1 0 48960 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_265
timestamp 1581449086
transform 1 0 48552 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_266
timestamp 1581449086
transform 1 0 47736 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_267
timestamp 1581449086
transform 1 0 47532 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_268
timestamp 1581449086
transform 1 0 47328 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_269
timestamp 1581449086
transform 1 0 46716 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_270
timestamp 1581449086
transform 1 0 46512 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_271
timestamp 1581449086
transform 1 0 46308 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_272
timestamp 1581449086
transform 1 0 45900 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_273
timestamp 1581449086
transform 1 0 45696 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_274
timestamp 1581449086
transform 1 0 45492 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_275
timestamp 1581449086
transform 1 0 45288 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_276
timestamp 1581449086
transform 1 0 44880 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_277
timestamp 1581449086
transform 1 0 44472 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_278
timestamp 1581449086
transform 1 0 43860 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_279
timestamp 1581449086
transform 1 0 43656 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_280
timestamp 1581449086
transform 1 0 43452 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_281
timestamp 1581449086
transform 1 0 43248 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_282
timestamp 1581449086
transform 1 0 42636 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_283
timestamp 1581449086
transform 1 0 42432 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_284
timestamp 1581449086
transform 1 0 42228 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_285
timestamp 1581449086
transform 1 0 42024 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_286
timestamp 1581449086
transform 1 0 41820 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_287
timestamp 1581449086
transform 1 0 41616 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_288
timestamp 1581449086
transform 1 0 41004 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_289
timestamp 1581449086
transform 1 0 40800 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_290
timestamp 1581449086
transform 1 0 40596 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_291
timestamp 1581449086
transform 1 0 40392 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_292
timestamp 1581449086
transform 1 0 40188 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_293
timestamp 1581449086
transform 1 0 39984 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_294
timestamp 1581449086
transform 1 0 39168 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_295
timestamp 1581449086
transform 1 0 38760 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_296
timestamp 1581449086
transform 1 0 38352 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_297
timestamp 1581449086
transform 1 0 37740 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_298
timestamp 1581449086
transform 1 0 37128 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_299
timestamp 1581449086
transform 1 0 36720 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_300
timestamp 1581449086
transform 1 0 36516 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_301
timestamp 1581449086
transform 1 0 36108 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_302
timestamp 1581449086
transform 1 0 35904 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_303
timestamp 1581449086
transform 1 0 35292 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_304
timestamp 1581449086
transform 1 0 35088 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_305
timestamp 1581449086
transform 1 0 34068 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_306
timestamp 1581449086
transform 1 0 33660 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_307
timestamp 1581449086
transform 1 0 33456 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_308
timestamp 1581449086
transform 1 0 33048 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_309
timestamp 1581449086
transform 1 0 32436 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_310
timestamp 1581449086
transform 1 0 31824 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_311
timestamp 1581449086
transform 1 0 31416 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_312
timestamp 1581449086
transform 1 0 30804 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_313
timestamp 1581449086
transform 1 0 30600 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_314
timestamp 1581449086
transform 1 0 30396 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_315
timestamp 1581449086
transform 1 0 30192 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_316
timestamp 1581449086
transform 1 0 29784 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_317
timestamp 1581449086
transform 1 0 29580 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_318
timestamp 1581449086
transform 1 0 29172 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_319
timestamp 1581449086
transform 1 0 28764 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_320
timestamp 1581449086
transform 1 0 28560 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_321
timestamp 1581449086
transform 1 0 28152 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_322
timestamp 1581449086
transform 1 0 27948 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_323
timestamp 1581449086
transform 1 0 27336 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_324
timestamp 1581449086
transform 1 0 26928 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_325
timestamp 1581449086
transform 1 0 26112 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_326
timestamp 1581449086
transform 1 0 25908 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_327
timestamp 1581449086
transform 1 0 25704 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_328
timestamp 1581449086
transform 1 0 25092 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_329
timestamp 1581449086
transform 1 0 24684 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_330
timestamp 1581449086
transform 1 0 24480 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_331
timestamp 1581449086
transform 1 0 23664 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_332
timestamp 1581449086
transform 1 0 23460 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_333
timestamp 1581449086
transform 1 0 22848 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_334
timestamp 1581449086
transform 1 0 22032 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_335
timestamp 1581449086
transform 1 0 21828 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_336
timestamp 1581449086
transform 1 0 21420 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_337
timestamp 1581449086
transform 1 0 21216 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_338
timestamp 1581449086
transform 1 0 20808 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_339
timestamp 1581449086
transform 1 0 20400 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_340
timestamp 1581449086
transform 1 0 19992 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_341
timestamp 1581449086
transform 1 0 19584 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_342
timestamp 1581449086
transform 1 0 19380 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_343
timestamp 1581449086
transform 1 0 19176 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_344
timestamp 1581449086
transform 1 0 18972 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_345
timestamp 1581449086
transform 1 0 18768 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_346
timestamp 1581449086
transform 1 0 17748 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_347
timestamp 1581449086
transform 1 0 17544 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_348
timestamp 1581449086
transform 1 0 17136 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_349
timestamp 1581449086
transform 1 0 16524 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_350
timestamp 1581449086
transform 1 0 16116 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_351
timestamp 1581449086
transform 1 0 15912 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_352
timestamp 1581449086
transform 1 0 15708 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_353
timestamp 1581449086
transform 1 0 15300 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_354
timestamp 1581449086
transform 1 0 15096 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_355
timestamp 1581449086
transform 1 0 14280 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_356
timestamp 1581449086
transform 1 0 13872 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_357
timestamp 1581449086
transform 1 0 13668 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_358
timestamp 1581449086
transform 1 0 13464 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_359
timestamp 1581449086
transform 1 0 13260 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_360
timestamp 1581449086
transform 1 0 13056 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_361
timestamp 1581449086
transform 1 0 11220 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_362
timestamp 1581449086
transform 1 0 11016 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_363
timestamp 1581449086
transform 1 0 9588 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_364
timestamp 1581449086
transform 1 0 9384 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_365
timestamp 1581449086
transform 1 0 9180 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_366
timestamp 1581449086
transform 1 0 8772 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_367
timestamp 1581449086
transform 1 0 8568 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_368
timestamp 1581449086
transform 1 0 8160 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_369
timestamp 1581449086
transform 1 0 7752 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_370
timestamp 1581449086
transform 1 0 7140 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_371
timestamp 1581449086
transform 1 0 6732 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_372
timestamp 1581449086
transform 1 0 6120 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_373
timestamp 1581449086
transform 1 0 5712 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_374
timestamp 1581449086
transform 1 0 5100 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_375
timestamp 1581449086
transform 1 0 4896 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_376
timestamp 1581449086
transform 1 0 4488 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_377
timestamp 1581449086
transform 1 0 4284 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_378
timestamp 1581449086
transform 1 0 3468 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_379
timestamp 1581449086
transform 1 0 3264 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_380
timestamp 1581449086
transform 1 0 3060 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_381
timestamp 1581449086
transform 1 0 1836 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_382
timestamp 1581449086
transform 1 0 1632 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_383
timestamp 1581449086
transform 1 0 1428 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_384
timestamp 1581449086
transform 1 0 1224 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_385
timestamp 1581449086
transform 1 0 1020 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_386
timestamp 1581449086
transform 1 0 816 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_387
timestamp 1581449086
transform 1 0 612 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_388
timestamp 1581449086
transform 1 0 408 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_389
timestamp 1581449086
transform 1 0 52020 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_390
timestamp 1581449086
transform 1 0 51816 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_391
timestamp 1581449086
transform 1 0 51408 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_392
timestamp 1581449086
transform 1 0 51204 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_393
timestamp 1581449086
transform 1 0 50388 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_394
timestamp 1581449086
transform 1 0 50184 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_395
timestamp 1581449086
transform 1 0 49980 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_396
timestamp 1581449086
transform 1 0 49776 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_397
timestamp 1581449086
transform 1 0 48960 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_398
timestamp 1581449086
transform 1 0 48552 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_399
timestamp 1581449086
transform 1 0 47940 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_400
timestamp 1581449086
transform 1 0 47736 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_401
timestamp 1581449086
transform 1 0 47328 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_402
timestamp 1581449086
transform 1 0 46920 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_403
timestamp 1581449086
transform 1 0 46716 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_404
timestamp 1581449086
transform 1 0 46104 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_405
timestamp 1581449086
transform 1 0 45900 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_406
timestamp 1581449086
transform 1 0 45492 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_407
timestamp 1581449086
transform 1 0 44880 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_408
timestamp 1581449086
transform 1 0 44676 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_409
timestamp 1581449086
transform 1 0 44064 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_410
timestamp 1581449086
transform 1 0 43860 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_411
timestamp 1581449086
transform 1 0 43248 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_412
timestamp 1581449086
transform 1 0 43044 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_413
timestamp 1581449086
transform 1 0 42228 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_414
timestamp 1581449086
transform 1 0 42024 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_415
timestamp 1581449086
transform 1 0 41820 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_416
timestamp 1581449086
transform 1 0 41208 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_417
timestamp 1581449086
transform 1 0 40596 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_418
timestamp 1581449086
transform 1 0 39984 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_419
timestamp 1581449086
transform 1 0 39780 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_420
timestamp 1581449086
transform 1 0 38964 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_421
timestamp 1581449086
transform 1 0 37944 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_422
timestamp 1581449086
transform 1 0 37536 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_423
timestamp 1581449086
transform 1 0 37332 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_424
timestamp 1581449086
transform 1 0 37128 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_425
timestamp 1581449086
transform 1 0 36924 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_426
timestamp 1581449086
transform 1 0 36312 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_427
timestamp 1581449086
transform 1 0 35700 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_428
timestamp 1581449086
transform 1 0 35088 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_429
timestamp 1581449086
transform 1 0 34884 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_430
timestamp 1581449086
transform 1 0 34680 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_431
timestamp 1581449086
transform 1 0 34476 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_432
timestamp 1581449086
transform 1 0 34068 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_433
timestamp 1581449086
transform 1 0 33864 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_434
timestamp 1581449086
transform 1 0 33660 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_435
timestamp 1581449086
transform 1 0 33456 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_436
timestamp 1581449086
transform 1 0 33252 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_437
timestamp 1581449086
transform 1 0 32844 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_438
timestamp 1581449086
transform 1 0 31620 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_439
timestamp 1581449086
transform 1 0 31416 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_440
timestamp 1581449086
transform 1 0 30804 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_441
timestamp 1581449086
transform 1 0 30396 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_442
timestamp 1581449086
transform 1 0 29988 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_443
timestamp 1581449086
transform 1 0 29784 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_444
timestamp 1581449086
transform 1 0 29580 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_445
timestamp 1581449086
transform 1 0 29172 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_446
timestamp 1581449086
transform 1 0 28968 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_447
timestamp 1581449086
transform 1 0 28152 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_448
timestamp 1581449086
transform 1 0 27948 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_449
timestamp 1581449086
transform 1 0 27744 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_450
timestamp 1581449086
transform 1 0 27336 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_451
timestamp 1581449086
transform 1 0 27132 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_452
timestamp 1581449086
transform 1 0 26724 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_453
timestamp 1581449086
transform 1 0 26112 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_454
timestamp 1581449086
transform 1 0 24684 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_455
timestamp 1581449086
transform 1 0 24276 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_456
timestamp 1581449086
transform 1 0 23052 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_457
timestamp 1581449086
transform 1 0 22644 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_458
timestamp 1581449086
transform 1 0 22440 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_459
timestamp 1581449086
transform 1 0 22032 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_460
timestamp 1581449086
transform 1 0 21420 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_461
timestamp 1581449086
transform 1 0 21216 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_462
timestamp 1581449086
transform 1 0 21012 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_463
timestamp 1581449086
transform 1 0 20808 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_464
timestamp 1581449086
transform 1 0 20604 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_465
timestamp 1581449086
transform 1 0 20400 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_466
timestamp 1581449086
transform 1 0 19992 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_467
timestamp 1581449086
transform 1 0 19176 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_468
timestamp 1581449086
transform 1 0 18972 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_469
timestamp 1581449086
transform 1 0 18768 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_470
timestamp 1581449086
transform 1 0 18564 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_471
timestamp 1581449086
transform 1 0 18156 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_472
timestamp 1581449086
transform 1 0 17748 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_473
timestamp 1581449086
transform 1 0 16932 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_474
timestamp 1581449086
transform 1 0 16524 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_475
timestamp 1581449086
transform 1 0 16320 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_476
timestamp 1581449086
transform 1 0 15708 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_477
timestamp 1581449086
transform 1 0 15096 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_478
timestamp 1581449086
transform 1 0 14280 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_479
timestamp 1581449086
transform 1 0 14076 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_480
timestamp 1581449086
transform 1 0 13668 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_481
timestamp 1581449086
transform 1 0 13056 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_482
timestamp 1581449086
transform 1 0 12648 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_483
timestamp 1581449086
transform 1 0 12240 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_484
timestamp 1581449086
transform 1 0 11832 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_485
timestamp 1581449086
transform 1 0 11424 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_486
timestamp 1581449086
transform 1 0 11016 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_487
timestamp 1581449086
transform 1 0 10812 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_488
timestamp 1581449086
transform 1 0 10200 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_489
timestamp 1581449086
transform 1 0 9996 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_490
timestamp 1581449086
transform 1 0 9180 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_491
timestamp 1581449086
transform 1 0 8772 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_492
timestamp 1581449086
transform 1 0 8568 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_493
timestamp 1581449086
transform 1 0 8364 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_494
timestamp 1581449086
transform 1 0 7956 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_495
timestamp 1581449086
transform 1 0 7752 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_496
timestamp 1581449086
transform 1 0 7548 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_497
timestamp 1581449086
transform 1 0 7344 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_498
timestamp 1581449086
transform 1 0 6732 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_499
timestamp 1581449086
transform 1 0 6528 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_500
timestamp 1581449086
transform 1 0 6120 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_501
timestamp 1581449086
transform 1 0 5712 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_502
timestamp 1581449086
transform 1 0 5508 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_503
timestamp 1581449086
transform 1 0 5100 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_504
timestamp 1581449086
transform 1 0 4896 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_505
timestamp 1581449086
transform 1 0 4692 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_506
timestamp 1581449086
transform 1 0 4080 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_507
timestamp 1581449086
transform 1 0 3876 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_508
timestamp 1581449086
transform 1 0 3672 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_509
timestamp 1581449086
transform 1 0 3060 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_510
timestamp 1581449086
transform 1 0 2856 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_511
timestamp 1581449086
transform 1 0 2652 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_512
timestamp 1581449086
transform 1 0 51816 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_513
timestamp 1581449086
transform 1 0 51408 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_514
timestamp 1581449086
transform 1 0 51204 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_515
timestamp 1581449086
transform 1 0 50796 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_516
timestamp 1581449086
transform 1 0 50592 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_517
timestamp 1581449086
transform 1 0 49572 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_518
timestamp 1581449086
transform 1 0 49164 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_519
timestamp 1581449086
transform 1 0 48552 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_520
timestamp 1581449086
transform 1 0 48348 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_521
timestamp 1581449086
transform 1 0 46512 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_522
timestamp 1581449086
transform 1 0 45900 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_523
timestamp 1581449086
transform 1 0 45492 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_524
timestamp 1581449086
transform 1 0 44880 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_525
timestamp 1581449086
transform 1 0 44472 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_526
timestamp 1581449086
transform 1 0 43860 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_527
timestamp 1581449086
transform 1 0 43452 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_528
timestamp 1581449086
transform 1 0 43044 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_529
timestamp 1581449086
transform 1 0 42840 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_530
timestamp 1581449086
transform 1 0 42432 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_531
timestamp 1581449086
transform 1 0 42228 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_532
timestamp 1581449086
transform 1 0 41208 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_533
timestamp 1581449086
transform 1 0 41004 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_534
timestamp 1581449086
transform 1 0 40392 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_535
timestamp 1581449086
transform 1 0 39780 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_536
timestamp 1581449086
transform 1 0 39168 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_537
timestamp 1581449086
transform 1 0 38760 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_538
timestamp 1581449086
transform 1 0 38148 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_539
timestamp 1581449086
transform 1 0 37944 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_540
timestamp 1581449086
transform 1 0 36924 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_541
timestamp 1581449086
transform 1 0 36312 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_542
timestamp 1581449086
transform 1 0 36108 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_543
timestamp 1581449086
transform 1 0 35496 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_544
timestamp 1581449086
transform 1 0 35292 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_545
timestamp 1581449086
transform 1 0 34476 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_546
timestamp 1581449086
transform 1 0 33456 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_547
timestamp 1581449086
transform 1 0 33048 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_548
timestamp 1581449086
transform 1 0 32640 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_549
timestamp 1581449086
transform 1 0 32232 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_550
timestamp 1581449086
transform 1 0 31620 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_551
timestamp 1581449086
transform 1 0 30804 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_552
timestamp 1581449086
transform 1 0 30600 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_553
timestamp 1581449086
transform 1 0 30192 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_554
timestamp 1581449086
transform 1 0 29580 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_555
timestamp 1581449086
transform 1 0 29376 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_556
timestamp 1581449086
transform 1 0 28560 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_557
timestamp 1581449086
transform 1 0 28356 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_558
timestamp 1581449086
transform 1 0 27948 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_559
timestamp 1581449086
transform 1 0 27744 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_560
timestamp 1581449086
transform 1 0 27540 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_561
timestamp 1581449086
transform 1 0 26928 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_562
timestamp 1581449086
transform 1 0 26520 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_563
timestamp 1581449086
transform 1 0 26112 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_564
timestamp 1581449086
transform 1 0 25500 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_565
timestamp 1581449086
transform 1 0 24888 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_566
timestamp 1581449086
transform 1 0 24480 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_567
timestamp 1581449086
transform 1 0 24276 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_568
timestamp 1581449086
transform 1 0 24072 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_569
timestamp 1581449086
transform 1 0 23664 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_570
timestamp 1581449086
transform 1 0 23256 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_571
timestamp 1581449086
transform 1 0 23052 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_572
timestamp 1581449086
transform 1 0 22848 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_573
timestamp 1581449086
transform 1 0 22440 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_574
timestamp 1581449086
transform 1 0 21828 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_575
timestamp 1581449086
transform 1 0 21216 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_576
timestamp 1581449086
transform 1 0 21012 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_577
timestamp 1581449086
transform 1 0 20808 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_578
timestamp 1581449086
transform 1 0 20604 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_579
timestamp 1581449086
transform 1 0 20196 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_580
timestamp 1581449086
transform 1 0 19992 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_581
timestamp 1581449086
transform 1 0 19788 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_582
timestamp 1581449086
transform 1 0 19584 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_583
timestamp 1581449086
transform 1 0 18972 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_584
timestamp 1581449086
transform 1 0 18768 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_585
timestamp 1581449086
transform 1 0 18156 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_586
timestamp 1581449086
transform 1 0 17952 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_587
timestamp 1581449086
transform 1 0 17748 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_588
timestamp 1581449086
transform 1 0 16932 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_589
timestamp 1581449086
transform 1 0 16320 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_590
timestamp 1581449086
transform 1 0 16116 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_591
timestamp 1581449086
transform 1 0 15300 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_592
timestamp 1581449086
transform 1 0 15096 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_593
timestamp 1581449086
transform 1 0 14076 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_594
timestamp 1581449086
transform 1 0 13872 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_595
timestamp 1581449086
transform 1 0 13056 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_596
timestamp 1581449086
transform 1 0 12240 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_597
timestamp 1581449086
transform 1 0 12036 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_598
timestamp 1581449086
transform 1 0 10812 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_599
timestamp 1581449086
transform 1 0 10404 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_600
timestamp 1581449086
transform 1 0 10200 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_601
timestamp 1581449086
transform 1 0 9792 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_602
timestamp 1581449086
transform 1 0 9384 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_603
timestamp 1581449086
transform 1 0 9180 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_604
timestamp 1581449086
transform 1 0 8772 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_605
timestamp 1581449086
transform 1 0 6732 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_606
timestamp 1581449086
transform 1 0 6324 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_607
timestamp 1581449086
transform 1 0 6120 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_608
timestamp 1581449086
transform 1 0 5916 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_609
timestamp 1581449086
transform 1 0 5712 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_610
timestamp 1581449086
transform 1 0 4488 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_611
timestamp 1581449086
transform 1 0 3468 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_612
timestamp 1581449086
transform 1 0 3264 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_613
timestamp 1581449086
transform 1 0 2856 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_614
timestamp 1581449086
transform 1 0 2652 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_615
timestamp 1581449086
transform 1 0 2448 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_616
timestamp 1581449086
transform 1 0 2244 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_617
timestamp 1581449086
transform 1 0 2040 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_618
timestamp 1581449086
transform 1 0 1224 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_619
timestamp 1581449086
transform 1 0 1020 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_620
timestamp 1581449086
transform 1 0 816 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_621
timestamp 1581449086
transform 1 0 612 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_622
timestamp 1581449086
transform 1 0 408 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_623
timestamp 1581449086
transform 1 0 204 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_624
timestamp 1581449086
transform 1 0 0 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_625
timestamp 1581449086
transform 1 0 52020 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_626
timestamp 1581449086
transform 1 0 51612 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_627
timestamp 1581449086
transform 1 0 51204 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_628
timestamp 1581449086
transform 1 0 50592 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_629
timestamp 1581449086
transform 1 0 50184 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_630
timestamp 1581449086
transform 1 0 49980 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_631
timestamp 1581449086
transform 1 0 49572 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_632
timestamp 1581449086
transform 1 0 48756 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_633
timestamp 1581449086
transform 1 0 48552 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_634
timestamp 1581449086
transform 1 0 48144 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_635
timestamp 1581449086
transform 1 0 47736 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_636
timestamp 1581449086
transform 1 0 47328 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_637
timestamp 1581449086
transform 1 0 46920 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_638
timestamp 1581449086
transform 1 0 46716 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_639
timestamp 1581449086
transform 1 0 46104 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_640
timestamp 1581449086
transform 1 0 45900 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_641
timestamp 1581449086
transform 1 0 45084 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_642
timestamp 1581449086
transform 1 0 44880 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_643
timestamp 1581449086
transform 1 0 44676 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_644
timestamp 1581449086
transform 1 0 44472 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_645
timestamp 1581449086
transform 1 0 44268 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_646
timestamp 1581449086
transform 1 0 43656 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_647
timestamp 1581449086
transform 1 0 43452 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_648
timestamp 1581449086
transform 1 0 42840 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_649
timestamp 1581449086
transform 1 0 42636 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_650
timestamp 1581449086
transform 1 0 41616 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_651
timestamp 1581449086
transform 1 0 41208 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_652
timestamp 1581449086
transform 1 0 40596 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_653
timestamp 1581449086
transform 1 0 40188 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_654
timestamp 1581449086
transform 1 0 39576 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_655
timestamp 1581449086
transform 1 0 39168 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_656
timestamp 1581449086
transform 1 0 38760 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_657
timestamp 1581449086
transform 1 0 38352 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_658
timestamp 1581449086
transform 1 0 38148 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_659
timestamp 1581449086
transform 1 0 37944 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_660
timestamp 1581449086
transform 1 0 37740 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_661
timestamp 1581449086
transform 1 0 36924 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_662
timestamp 1581449086
transform 1 0 36720 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_663
timestamp 1581449086
transform 1 0 35904 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_664
timestamp 1581449086
transform 1 0 35700 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_665
timestamp 1581449086
transform 1 0 34884 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_666
timestamp 1581449086
transform 1 0 34680 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_667
timestamp 1581449086
transform 1 0 34068 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_668
timestamp 1581449086
transform 1 0 33864 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_669
timestamp 1581449086
transform 1 0 33660 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_670
timestamp 1581449086
transform 1 0 33252 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_671
timestamp 1581449086
transform 1 0 33048 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_672
timestamp 1581449086
transform 1 0 32640 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_673
timestamp 1581449086
transform 1 0 31824 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_674
timestamp 1581449086
transform 1 0 30804 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_675
timestamp 1581449086
transform 1 0 30192 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_676
timestamp 1581449086
transform 1 0 29784 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_677
timestamp 1581449086
transform 1 0 29580 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_678
timestamp 1581449086
transform 1 0 28968 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_679
timestamp 1581449086
transform 1 0 28560 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_680
timestamp 1581449086
transform 1 0 28152 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_681
timestamp 1581449086
transform 1 0 27336 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_682
timestamp 1581449086
transform 1 0 24684 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_683
timestamp 1581449086
transform 1 0 24480 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_684
timestamp 1581449086
transform 1 0 24276 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_685
timestamp 1581449086
transform 1 0 24072 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_686
timestamp 1581449086
transform 1 0 23868 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_687
timestamp 1581449086
transform 1 0 23664 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_688
timestamp 1581449086
transform 1 0 23052 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_689
timestamp 1581449086
transform 1 0 22848 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_690
timestamp 1581449086
transform 1 0 21624 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_691
timestamp 1581449086
transform 1 0 21216 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_692
timestamp 1581449086
transform 1 0 20604 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_693
timestamp 1581449086
transform 1 0 20400 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_694
timestamp 1581449086
transform 1 0 20196 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_695
timestamp 1581449086
transform 1 0 19992 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_696
timestamp 1581449086
transform 1 0 19788 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_697
timestamp 1581449086
transform 1 0 19380 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_698
timestamp 1581449086
transform 1 0 18564 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_699
timestamp 1581449086
transform 1 0 18156 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_700
timestamp 1581449086
transform 1 0 17952 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_701
timestamp 1581449086
transform 1 0 17748 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_702
timestamp 1581449086
transform 1 0 17340 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_703
timestamp 1581449086
transform 1 0 16932 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_704
timestamp 1581449086
transform 1 0 16728 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_705
timestamp 1581449086
transform 1 0 16320 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_706
timestamp 1581449086
transform 1 0 16116 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_707
timestamp 1581449086
transform 1 0 15912 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_708
timestamp 1581449086
transform 1 0 15708 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_709
timestamp 1581449086
transform 1 0 14280 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_710
timestamp 1581449086
transform 1 0 13056 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_711
timestamp 1581449086
transform 1 0 12648 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_712
timestamp 1581449086
transform 1 0 12240 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_713
timestamp 1581449086
transform 1 0 12036 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_714
timestamp 1581449086
transform 1 0 11832 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_715
timestamp 1581449086
transform 1 0 11424 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_716
timestamp 1581449086
transform 1 0 11220 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_717
timestamp 1581449086
transform 1 0 10812 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_718
timestamp 1581449086
transform 1 0 10404 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_719
timestamp 1581449086
transform 1 0 9996 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_720
timestamp 1581449086
transform 1 0 9792 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_721
timestamp 1581449086
transform 1 0 9180 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_722
timestamp 1581449086
transform 1 0 8976 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_723
timestamp 1581449086
transform 1 0 8568 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_724
timestamp 1581449086
transform 1 0 8364 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_725
timestamp 1581449086
transform 1 0 8160 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_726
timestamp 1581449086
transform 1 0 6936 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_727
timestamp 1581449086
transform 1 0 6732 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_728
timestamp 1581449086
transform 1 0 6324 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_729
timestamp 1581449086
transform 1 0 5916 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_730
timestamp 1581449086
transform 1 0 5508 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_731
timestamp 1581449086
transform 1 0 4284 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_732
timestamp 1581449086
transform 1 0 4080 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_733
timestamp 1581449086
transform 1 0 3468 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_734
timestamp 1581449086
transform 1 0 3264 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_735
timestamp 1581449086
transform 1 0 2652 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_736
timestamp 1581449086
transform 1 0 2448 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_737
timestamp 1581449086
transform 1 0 2244 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_738
timestamp 1581449086
transform 1 0 2040 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_739
timestamp 1581449086
transform 1 0 1428 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_740
timestamp 1581449086
transform 1 0 1224 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_741
timestamp 1581449086
transform 1 0 52020 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_742
timestamp 1581449086
transform 1 0 51816 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_743
timestamp 1581449086
transform 1 0 51612 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_744
timestamp 1581449086
transform 1 0 51408 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_745
timestamp 1581449086
transform 1 0 51204 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_746
timestamp 1581449086
transform 1 0 50796 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_747
timestamp 1581449086
transform 1 0 50388 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_748
timestamp 1581449086
transform 1 0 49980 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_749
timestamp 1581449086
transform 1 0 49776 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_750
timestamp 1581449086
transform 1 0 49572 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_751
timestamp 1581449086
transform 1 0 48960 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_752
timestamp 1581449086
transform 1 0 48756 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_753
timestamp 1581449086
transform 1 0 48348 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_754
timestamp 1581449086
transform 1 0 47940 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_755
timestamp 1581449086
transform 1 0 47532 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_756
timestamp 1581449086
transform 1 0 46104 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_757
timestamp 1581449086
transform 1 0 45900 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_758
timestamp 1581449086
transform 1 0 45288 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_759
timestamp 1581449086
transform 1 0 44880 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_760
timestamp 1581449086
transform 1 0 44064 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_761
timestamp 1581449086
transform 1 0 43860 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_762
timestamp 1581449086
transform 1 0 43248 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_763
timestamp 1581449086
transform 1 0 42636 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_764
timestamp 1581449086
transform 1 0 42228 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_765
timestamp 1581449086
transform 1 0 42024 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_766
timestamp 1581449086
transform 1 0 41820 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_767
timestamp 1581449086
transform 1 0 41616 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_768
timestamp 1581449086
transform 1 0 41412 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_769
timestamp 1581449086
transform 1 0 41208 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_770
timestamp 1581449086
transform 1 0 41004 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_771
timestamp 1581449086
transform 1 0 40800 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_772
timestamp 1581449086
transform 1 0 39984 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_773
timestamp 1581449086
transform 1 0 39780 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_774
timestamp 1581449086
transform 1 0 39576 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_775
timestamp 1581449086
transform 1 0 38964 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_776
timestamp 1581449086
transform 1 0 38760 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_777
timestamp 1581449086
transform 1 0 38556 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_778
timestamp 1581449086
transform 1 0 38352 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_779
timestamp 1581449086
transform 1 0 38148 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_780
timestamp 1581449086
transform 1 0 37944 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_781
timestamp 1581449086
transform 1 0 37536 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_782
timestamp 1581449086
transform 1 0 37128 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_783
timestamp 1581449086
transform 1 0 36720 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_784
timestamp 1581449086
transform 1 0 36516 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_785
timestamp 1581449086
transform 1 0 36312 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_786
timestamp 1581449086
transform 1 0 36108 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_787
timestamp 1581449086
transform 1 0 34884 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_788
timestamp 1581449086
transform 1 0 34680 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_789
timestamp 1581449086
transform 1 0 34476 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_790
timestamp 1581449086
transform 1 0 34068 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_791
timestamp 1581449086
transform 1 0 33456 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_792
timestamp 1581449086
transform 1 0 33252 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_793
timestamp 1581449086
transform 1 0 32028 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_794
timestamp 1581449086
transform 1 0 31620 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_795
timestamp 1581449086
transform 1 0 31008 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_796
timestamp 1581449086
transform 1 0 30804 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_797
timestamp 1581449086
transform 1 0 30600 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_798
timestamp 1581449086
transform 1 0 29988 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_799
timestamp 1581449086
transform 1 0 29784 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_800
timestamp 1581449086
transform 1 0 28968 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_801
timestamp 1581449086
transform 1 0 28356 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_802
timestamp 1581449086
transform 1 0 27948 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_803
timestamp 1581449086
transform 1 0 27744 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_804
timestamp 1581449086
transform 1 0 27132 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_805
timestamp 1581449086
transform 1 0 26316 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_806
timestamp 1581449086
transform 1 0 25908 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_807
timestamp 1581449086
transform 1 0 25500 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_808
timestamp 1581449086
transform 1 0 25092 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_809
timestamp 1581449086
transform 1 0 24888 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_810
timestamp 1581449086
transform 1 0 24684 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_811
timestamp 1581449086
transform 1 0 24072 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_812
timestamp 1581449086
transform 1 0 23868 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_813
timestamp 1581449086
transform 1 0 23256 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_814
timestamp 1581449086
transform 1 0 22848 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_815
timestamp 1581449086
transform 1 0 22236 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_816
timestamp 1581449086
transform 1 0 21216 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_817
timestamp 1581449086
transform 1 0 21012 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_818
timestamp 1581449086
transform 1 0 20808 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_819
timestamp 1581449086
transform 1 0 20196 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_820
timestamp 1581449086
transform 1 0 19584 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_821
timestamp 1581449086
transform 1 0 18564 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_822
timestamp 1581449086
transform 1 0 18156 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_823
timestamp 1581449086
transform 1 0 17952 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_824
timestamp 1581449086
transform 1 0 17748 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_825
timestamp 1581449086
transform 1 0 17340 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_826
timestamp 1581449086
transform 1 0 17136 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_827
timestamp 1581449086
transform 1 0 16524 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_828
timestamp 1581449086
transform 1 0 16320 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_829
timestamp 1581449086
transform 1 0 15912 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_830
timestamp 1581449086
transform 1 0 15504 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_831
timestamp 1581449086
transform 1 0 15300 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_832
timestamp 1581449086
transform 1 0 14280 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_833
timestamp 1581449086
transform 1 0 14076 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_834
timestamp 1581449086
transform 1 0 13872 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_835
timestamp 1581449086
transform 1 0 12444 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_836
timestamp 1581449086
transform 1 0 12036 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_837
timestamp 1581449086
transform 1 0 11016 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_838
timestamp 1581449086
transform 1 0 10608 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_839
timestamp 1581449086
transform 1 0 10404 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_840
timestamp 1581449086
transform 1 0 9588 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_841
timestamp 1581449086
transform 1 0 9384 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_842
timestamp 1581449086
transform 1 0 9180 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_843
timestamp 1581449086
transform 1 0 8976 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_844
timestamp 1581449086
transform 1 0 8772 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_845
timestamp 1581449086
transform 1 0 7140 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_846
timestamp 1581449086
transform 1 0 6732 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_847
timestamp 1581449086
transform 1 0 6528 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_848
timestamp 1581449086
transform 1 0 6324 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_849
timestamp 1581449086
transform 1 0 5916 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_850
timestamp 1581449086
transform 1 0 5508 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_851
timestamp 1581449086
transform 1 0 5304 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_852
timestamp 1581449086
transform 1 0 4896 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_853
timestamp 1581449086
transform 1 0 3876 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_854
timestamp 1581449086
transform 1 0 3672 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_855
timestamp 1581449086
transform 1 0 3468 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_856
timestamp 1581449086
transform 1 0 2652 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_857
timestamp 1581449086
transform 1 0 2448 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_858
timestamp 1581449086
transform 1 0 1020 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_859
timestamp 1581449086
transform 1 0 816 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_860
timestamp 1581449086
transform 1 0 612 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_861
timestamp 1581449086
transform 1 0 408 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_862
timestamp 1581449086
transform 1 0 204 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_863
timestamp 1581449086
transform 1 0 0 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_864
timestamp 1581449086
transform 1 0 51408 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_865
timestamp 1581449086
transform 1 0 50592 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_866
timestamp 1581449086
transform 1 0 50388 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_867
timestamp 1581449086
transform 1 0 49980 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_868
timestamp 1581449086
transform 1 0 49776 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_869
timestamp 1581449086
transform 1 0 49368 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_870
timestamp 1581449086
transform 1 0 49164 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_871
timestamp 1581449086
transform 1 0 48552 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_872
timestamp 1581449086
transform 1 0 48144 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_873
timestamp 1581449086
transform 1 0 47940 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_874
timestamp 1581449086
transform 1 0 47736 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_875
timestamp 1581449086
transform 1 0 47532 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_876
timestamp 1581449086
transform 1 0 47124 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_877
timestamp 1581449086
transform 1 0 46920 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_878
timestamp 1581449086
transform 1 0 46716 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_879
timestamp 1581449086
transform 1 0 46512 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_880
timestamp 1581449086
transform 1 0 46308 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_881
timestamp 1581449086
transform 1 0 45492 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_882
timestamp 1581449086
transform 1 0 45288 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_883
timestamp 1581449086
transform 1 0 43452 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_884
timestamp 1581449086
transform 1 0 43248 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_885
timestamp 1581449086
transform 1 0 42228 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_886
timestamp 1581449086
transform 1 0 42024 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_887
timestamp 1581449086
transform 1 0 41616 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_888
timestamp 1581449086
transform 1 0 41412 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_889
timestamp 1581449086
transform 1 0 41208 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_890
timestamp 1581449086
transform 1 0 40800 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_891
timestamp 1581449086
transform 1 0 40596 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_892
timestamp 1581449086
transform 1 0 40392 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_893
timestamp 1581449086
transform 1 0 40188 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_894
timestamp 1581449086
transform 1 0 39780 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_895
timestamp 1581449086
transform 1 0 39576 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_896
timestamp 1581449086
transform 1 0 39372 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_897
timestamp 1581449086
transform 1 0 39168 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_898
timestamp 1581449086
transform 1 0 38760 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_899
timestamp 1581449086
transform 1 0 38148 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_900
timestamp 1581449086
transform 1 0 37944 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_901
timestamp 1581449086
transform 1 0 37740 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_902
timestamp 1581449086
transform 1 0 37536 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_903
timestamp 1581449086
transform 1 0 36108 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_904
timestamp 1581449086
transform 1 0 35292 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_905
timestamp 1581449086
transform 1 0 35088 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_906
timestamp 1581449086
transform 1 0 34680 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_907
timestamp 1581449086
transform 1 0 34476 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_908
timestamp 1581449086
transform 1 0 34068 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_909
timestamp 1581449086
transform 1 0 33864 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_910
timestamp 1581449086
transform 1 0 33456 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_911
timestamp 1581449086
transform 1 0 33048 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_912
timestamp 1581449086
transform 1 0 32640 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_913
timestamp 1581449086
transform 1 0 31416 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_914
timestamp 1581449086
transform 1 0 30600 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_915
timestamp 1581449086
transform 1 0 30192 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_916
timestamp 1581449086
transform 1 0 29988 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_917
timestamp 1581449086
transform 1 0 29376 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_918
timestamp 1581449086
transform 1 0 27948 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_919
timestamp 1581449086
transform 1 0 27744 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_920
timestamp 1581449086
transform 1 0 27540 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_921
timestamp 1581449086
transform 1 0 27336 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_922
timestamp 1581449086
transform 1 0 27132 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_923
timestamp 1581449086
transform 1 0 26724 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_924
timestamp 1581449086
transform 1 0 26520 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_925
timestamp 1581449086
transform 1 0 25908 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_926
timestamp 1581449086
transform 1 0 25296 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_927
timestamp 1581449086
transform 1 0 24888 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_928
timestamp 1581449086
transform 1 0 24480 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_929
timestamp 1581449086
transform 1 0 23052 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_930
timestamp 1581449086
transform 1 0 22848 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_931
timestamp 1581449086
transform 1 0 22236 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_932
timestamp 1581449086
transform 1 0 21828 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_933
timestamp 1581449086
transform 1 0 21420 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_934
timestamp 1581449086
transform 1 0 21012 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_935
timestamp 1581449086
transform 1 0 20400 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_936
timestamp 1581449086
transform 1 0 20196 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_937
timestamp 1581449086
transform 1 0 19788 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_938
timestamp 1581449086
transform 1 0 19584 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_939
timestamp 1581449086
transform 1 0 19380 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_940
timestamp 1581449086
transform 1 0 19176 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_941
timestamp 1581449086
transform 1 0 18972 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_942
timestamp 1581449086
transform 1 0 18156 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_943
timestamp 1581449086
transform 1 0 17952 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_944
timestamp 1581449086
transform 1 0 17748 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_945
timestamp 1581449086
transform 1 0 17544 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_946
timestamp 1581449086
transform 1 0 17340 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_947
timestamp 1581449086
transform 1 0 17136 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_948
timestamp 1581449086
transform 1 0 16524 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_949
timestamp 1581449086
transform 1 0 16116 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_950
timestamp 1581449086
transform 1 0 15708 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_951
timestamp 1581449086
transform 1 0 15504 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_952
timestamp 1581449086
transform 1 0 15096 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_953
timestamp 1581449086
transform 1 0 14484 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_954
timestamp 1581449086
transform 1 0 14280 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_955
timestamp 1581449086
transform 1 0 13872 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_956
timestamp 1581449086
transform 1 0 13464 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_957
timestamp 1581449086
transform 1 0 13260 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_958
timestamp 1581449086
transform 1 0 13056 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_959
timestamp 1581449086
transform 1 0 12240 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_960
timestamp 1581449086
transform 1 0 11832 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_961
timestamp 1581449086
transform 1 0 11628 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_962
timestamp 1581449086
transform 1 0 11220 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_963
timestamp 1581449086
transform 1 0 10812 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_964
timestamp 1581449086
transform 1 0 10200 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_965
timestamp 1581449086
transform 1 0 9996 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_966
timestamp 1581449086
transform 1 0 9588 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_967
timestamp 1581449086
transform 1 0 9384 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_968
timestamp 1581449086
transform 1 0 8976 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_969
timestamp 1581449086
transform 1 0 8772 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_970
timestamp 1581449086
transform 1 0 8568 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_971
timestamp 1581449086
transform 1 0 8364 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_972
timestamp 1581449086
transform 1 0 8160 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_973
timestamp 1581449086
transform 1 0 7752 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_974
timestamp 1581449086
transform 1 0 7548 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_975
timestamp 1581449086
transform 1 0 7344 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_976
timestamp 1581449086
transform 1 0 6936 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_977
timestamp 1581449086
transform 1 0 6732 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_978
timestamp 1581449086
transform 1 0 6324 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_979
timestamp 1581449086
transform 1 0 6120 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_980
timestamp 1581449086
transform 1 0 4692 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_981
timestamp 1581449086
transform 1 0 4080 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_982
timestamp 1581449086
transform 1 0 3876 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_983
timestamp 1581449086
transform 1 0 3468 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_984
timestamp 1581449086
transform 1 0 3264 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_985
timestamp 1581449086
transform 1 0 3060 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_986
timestamp 1581449086
transform 1 0 2856 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_987
timestamp 1581449086
transform 1 0 2652 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_988
timestamp 1581449086
transform 1 0 1836 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_989
timestamp 1581449086
transform 1 0 1632 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_990
timestamp 1581449086
transform 1 0 204 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_991
timestamp 1581449086
transform 1 0 0 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_992
timestamp 1581449086
transform 1 0 51816 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_993
timestamp 1581449086
transform 1 0 51204 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_994
timestamp 1581449086
transform 1 0 50796 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_995
timestamp 1581449086
transform 1 0 50184 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_996
timestamp 1581449086
transform 1 0 49980 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_997
timestamp 1581449086
transform 1 0 49572 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_998
timestamp 1581449086
transform 1 0 49368 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_999
timestamp 1581449086
transform 1 0 48756 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1000
timestamp 1581449086
transform 1 0 48552 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1001
timestamp 1581449086
transform 1 0 48348 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1002
timestamp 1581449086
transform 1 0 48144 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1003
timestamp 1581449086
transform 1 0 47736 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1004
timestamp 1581449086
transform 1 0 46716 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1005
timestamp 1581449086
transform 1 0 46104 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1006
timestamp 1581449086
transform 1 0 45696 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1007
timestamp 1581449086
transform 1 0 45492 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1008
timestamp 1581449086
transform 1 0 45084 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1009
timestamp 1581449086
transform 1 0 44880 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1010
timestamp 1581449086
transform 1 0 44472 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1011
timestamp 1581449086
transform 1 0 44064 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1012
timestamp 1581449086
transform 1 0 43860 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1013
timestamp 1581449086
transform 1 0 43656 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1014
timestamp 1581449086
transform 1 0 43452 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1015
timestamp 1581449086
transform 1 0 43248 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1016
timestamp 1581449086
transform 1 0 42840 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1017
timestamp 1581449086
transform 1 0 42228 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1018
timestamp 1581449086
transform 1 0 41820 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1019
timestamp 1581449086
transform 1 0 41616 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1020
timestamp 1581449086
transform 1 0 41412 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1021
timestamp 1581449086
transform 1 0 40392 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1022
timestamp 1581449086
transform 1 0 40188 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1023
timestamp 1581449086
transform 1 0 39780 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1024
timestamp 1581449086
transform 1 0 39576 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1025
timestamp 1581449086
transform 1 0 39168 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1026
timestamp 1581449086
transform 1 0 38964 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1027
timestamp 1581449086
transform 1 0 38556 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1028
timestamp 1581449086
transform 1 0 38352 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1029
timestamp 1581449086
transform 1 0 38148 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1030
timestamp 1581449086
transform 1 0 37944 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1031
timestamp 1581449086
transform 1 0 37740 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1032
timestamp 1581449086
transform 1 0 37128 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1033
timestamp 1581449086
transform 1 0 36108 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1034
timestamp 1581449086
transform 1 0 35904 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1035
timestamp 1581449086
transform 1 0 35496 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1036
timestamp 1581449086
transform 1 0 35088 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1037
timestamp 1581449086
transform 1 0 34884 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1038
timestamp 1581449086
transform 1 0 34680 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1039
timestamp 1581449086
transform 1 0 33456 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1040
timestamp 1581449086
transform 1 0 33252 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1041
timestamp 1581449086
transform 1 0 32844 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1042
timestamp 1581449086
transform 1 0 32640 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1043
timestamp 1581449086
transform 1 0 32436 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1044
timestamp 1581449086
transform 1 0 32028 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1045
timestamp 1581449086
transform 1 0 31824 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1046
timestamp 1581449086
transform 1 0 31620 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1047
timestamp 1581449086
transform 1 0 31212 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1048
timestamp 1581449086
transform 1 0 30804 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1049
timestamp 1581449086
transform 1 0 30396 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1050
timestamp 1581449086
transform 1 0 29988 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1051
timestamp 1581449086
transform 1 0 29376 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1052
timestamp 1581449086
transform 1 0 29172 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1053
timestamp 1581449086
transform 1 0 28560 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1054
timestamp 1581449086
transform 1 0 28356 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1055
timestamp 1581449086
transform 1 0 27948 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1056
timestamp 1581449086
transform 1 0 27540 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1057
timestamp 1581449086
transform 1 0 27132 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1058
timestamp 1581449086
transform 1 0 26520 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1059
timestamp 1581449086
transform 1 0 26112 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1060
timestamp 1581449086
transform 1 0 25908 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1061
timestamp 1581449086
transform 1 0 24888 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1062
timestamp 1581449086
transform 1 0 24684 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1063
timestamp 1581449086
transform 1 0 24480 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1064
timestamp 1581449086
transform 1 0 24276 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1065
timestamp 1581449086
transform 1 0 23868 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1066
timestamp 1581449086
transform 1 0 23664 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1067
timestamp 1581449086
transform 1 0 23052 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1068
timestamp 1581449086
transform 1 0 22848 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1069
timestamp 1581449086
transform 1 0 22440 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1070
timestamp 1581449086
transform 1 0 22236 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1071
timestamp 1581449086
transform 1 0 22032 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1072
timestamp 1581449086
transform 1 0 21828 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1073
timestamp 1581449086
transform 1 0 21216 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1074
timestamp 1581449086
transform 1 0 21012 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1075
timestamp 1581449086
transform 1 0 20808 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1076
timestamp 1581449086
transform 1 0 20604 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1077
timestamp 1581449086
transform 1 0 20400 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1078
timestamp 1581449086
transform 1 0 20196 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1079
timestamp 1581449086
transform 1 0 19380 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1080
timestamp 1581449086
transform 1 0 19176 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1081
timestamp 1581449086
transform 1 0 18972 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1082
timestamp 1581449086
transform 1 0 18768 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1083
timestamp 1581449086
transform 1 0 18360 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1084
timestamp 1581449086
transform 1 0 17136 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1085
timestamp 1581449086
transform 1 0 16728 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1086
timestamp 1581449086
transform 1 0 15912 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1087
timestamp 1581449086
transform 1 0 15708 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1088
timestamp 1581449086
transform 1 0 14484 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1089
timestamp 1581449086
transform 1 0 14280 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1090
timestamp 1581449086
transform 1 0 14076 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1091
timestamp 1581449086
transform 1 0 13872 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1092
timestamp 1581449086
transform 1 0 13260 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1093
timestamp 1581449086
transform 1 0 12852 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1094
timestamp 1581449086
transform 1 0 12648 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1095
timestamp 1581449086
transform 1 0 12036 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1096
timestamp 1581449086
transform 1 0 11016 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1097
timestamp 1581449086
transform 1 0 10608 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1098
timestamp 1581449086
transform 1 0 9996 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1099
timestamp 1581449086
transform 1 0 8772 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1100
timestamp 1581449086
transform 1 0 8568 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1101
timestamp 1581449086
transform 1 0 7752 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1102
timestamp 1581449086
transform 1 0 6528 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1103
timestamp 1581449086
transform 1 0 6120 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1104
timestamp 1581449086
transform 1 0 5712 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1105
timestamp 1581449086
transform 1 0 5508 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1106
timestamp 1581449086
transform 1 0 5100 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1107
timestamp 1581449086
transform 1 0 4896 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1108
timestamp 1581449086
transform 1 0 4080 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1109
timestamp 1581449086
transform 1 0 3672 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1110
timestamp 1581449086
transform 1 0 3060 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1111
timestamp 1581449086
transform 1 0 2448 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1112
timestamp 1581449086
transform 1 0 2244 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1113
timestamp 1581449086
transform 1 0 1632 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1114
timestamp 1581449086
transform 1 0 1428 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1115
timestamp 1581449086
transform 1 0 1224 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1116
timestamp 1581449086
transform 1 0 1020 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1117
timestamp 1581449086
transform 1 0 0 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1118
timestamp 1581449086
transform 1 0 52020 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1119
timestamp 1581449086
transform 1 0 51612 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1120
timestamp 1581449086
transform 1 0 51408 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1121
timestamp 1581449086
transform 1 0 51204 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1122
timestamp 1581449086
transform 1 0 51000 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1123
timestamp 1581449086
transform 1 0 50796 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1124
timestamp 1581449086
transform 1 0 49776 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1125
timestamp 1581449086
transform 1 0 49368 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1126
timestamp 1581449086
transform 1 0 48756 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1127
timestamp 1581449086
transform 1 0 48552 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1128
timestamp 1581449086
transform 1 0 47940 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1129
timestamp 1581449086
transform 1 0 47736 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1130
timestamp 1581449086
transform 1 0 46512 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1131
timestamp 1581449086
transform 1 0 46104 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1132
timestamp 1581449086
transform 1 0 45696 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1133
timestamp 1581449086
transform 1 0 45492 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1134
timestamp 1581449086
transform 1 0 45084 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1135
timestamp 1581449086
transform 1 0 44880 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1136
timestamp 1581449086
transform 1 0 44268 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1137
timestamp 1581449086
transform 1 0 44064 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1138
timestamp 1581449086
transform 1 0 43656 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1139
timestamp 1581449086
transform 1 0 43452 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1140
timestamp 1581449086
transform 1 0 43044 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1141
timestamp 1581449086
transform 1 0 42228 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1142
timestamp 1581449086
transform 1 0 41820 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1143
timestamp 1581449086
transform 1 0 41616 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1144
timestamp 1581449086
transform 1 0 41208 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1145
timestamp 1581449086
transform 1 0 40596 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1146
timestamp 1581449086
transform 1 0 40392 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1147
timestamp 1581449086
transform 1 0 40188 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1148
timestamp 1581449086
transform 1 0 39780 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1149
timestamp 1581449086
transform 1 0 39576 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1150
timestamp 1581449086
transform 1 0 39372 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1151
timestamp 1581449086
transform 1 0 39168 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1152
timestamp 1581449086
transform 1 0 38556 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1153
timestamp 1581449086
transform 1 0 38148 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1154
timestamp 1581449086
transform 1 0 37944 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1155
timestamp 1581449086
transform 1 0 37536 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1156
timestamp 1581449086
transform 1 0 37332 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1157
timestamp 1581449086
transform 1 0 37128 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1158
timestamp 1581449086
transform 1 0 36720 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1159
timestamp 1581449086
transform 1 0 36516 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1160
timestamp 1581449086
transform 1 0 36312 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1161
timestamp 1581449086
transform 1 0 35904 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1162
timestamp 1581449086
transform 1 0 35700 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1163
timestamp 1581449086
transform 1 0 34476 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1164
timestamp 1581449086
transform 1 0 34272 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1165
timestamp 1581449086
transform 1 0 34068 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1166
timestamp 1581449086
transform 1 0 33252 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1167
timestamp 1581449086
transform 1 0 33048 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1168
timestamp 1581449086
transform 1 0 32640 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1169
timestamp 1581449086
transform 1 0 32436 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1170
timestamp 1581449086
transform 1 0 32028 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1171
timestamp 1581449086
transform 1 0 31620 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1172
timestamp 1581449086
transform 1 0 31416 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1173
timestamp 1581449086
transform 1 0 29784 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1174
timestamp 1581449086
transform 1 0 29376 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1175
timestamp 1581449086
transform 1 0 29172 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1176
timestamp 1581449086
transform 1 0 28560 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1177
timestamp 1581449086
transform 1 0 28356 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1178
timestamp 1581449086
transform 1 0 28152 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1179
timestamp 1581449086
transform 1 0 27948 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1180
timestamp 1581449086
transform 1 0 27336 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1181
timestamp 1581449086
transform 1 0 26928 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1182
timestamp 1581449086
transform 1 0 26724 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1183
timestamp 1581449086
transform 1 0 26520 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1184
timestamp 1581449086
transform 1 0 25704 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1185
timestamp 1581449086
transform 1 0 25500 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1186
timestamp 1581449086
transform 1 0 25092 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1187
timestamp 1581449086
transform 1 0 24684 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1188
timestamp 1581449086
transform 1 0 24072 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1189
timestamp 1581449086
transform 1 0 23664 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1190
timestamp 1581449086
transform 1 0 23052 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1191
timestamp 1581449086
transform 1 0 22848 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1192
timestamp 1581449086
transform 1 0 22644 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1193
timestamp 1581449086
transform 1 0 22440 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1194
timestamp 1581449086
transform 1 0 22032 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1195
timestamp 1581449086
transform 1 0 21828 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1196
timestamp 1581449086
transform 1 0 21420 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1197
timestamp 1581449086
transform 1 0 21012 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1198
timestamp 1581449086
transform 1 0 20808 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1199
timestamp 1581449086
transform 1 0 19584 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1200
timestamp 1581449086
transform 1 0 19380 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1201
timestamp 1581449086
transform 1 0 19176 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1202
timestamp 1581449086
transform 1 0 18972 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1203
timestamp 1581449086
transform 1 0 18768 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1204
timestamp 1581449086
transform 1 0 18564 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1205
timestamp 1581449086
transform 1 0 18156 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1206
timestamp 1581449086
transform 1 0 17544 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1207
timestamp 1581449086
transform 1 0 17340 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1208
timestamp 1581449086
transform 1 0 16932 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1209
timestamp 1581449086
transform 1 0 16524 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1210
timestamp 1581449086
transform 1 0 15708 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1211
timestamp 1581449086
transform 1 0 15504 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1212
timestamp 1581449086
transform 1 0 15096 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1213
timestamp 1581449086
transform 1 0 14076 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1214
timestamp 1581449086
transform 1 0 13668 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1215
timestamp 1581449086
transform 1 0 13464 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1216
timestamp 1581449086
transform 1 0 13056 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1217
timestamp 1581449086
transform 1 0 12852 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1218
timestamp 1581449086
transform 1 0 12444 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1219
timestamp 1581449086
transform 1 0 12240 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1220
timestamp 1581449086
transform 1 0 12036 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1221
timestamp 1581449086
transform 1 0 11832 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1222
timestamp 1581449086
transform 1 0 11628 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1223
timestamp 1581449086
transform 1 0 11220 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1224
timestamp 1581449086
transform 1 0 11016 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1225
timestamp 1581449086
transform 1 0 9792 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1226
timestamp 1581449086
transform 1 0 8568 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1227
timestamp 1581449086
transform 1 0 7956 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1228
timestamp 1581449086
transform 1 0 7548 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1229
timestamp 1581449086
transform 1 0 7344 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1230
timestamp 1581449086
transform 1 0 7140 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1231
timestamp 1581449086
transform 1 0 6120 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1232
timestamp 1581449086
transform 1 0 5916 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1233
timestamp 1581449086
transform 1 0 5712 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1234
timestamp 1581449086
transform 1 0 5304 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1235
timestamp 1581449086
transform 1 0 5100 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1236
timestamp 1581449086
transform 1 0 4692 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1237
timestamp 1581449086
transform 1 0 4080 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1238
timestamp 1581449086
transform 1 0 3876 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1239
timestamp 1581449086
transform 1 0 3672 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1240
timestamp 1581449086
transform 1 0 3468 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1241
timestamp 1581449086
transform 1 0 2652 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1242
timestamp 1581449086
transform 1 0 2244 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1243
timestamp 1581449086
transform 1 0 1836 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1244
timestamp 1581449086
transform 1 0 1632 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1245
timestamp 1581449086
transform 1 0 1428 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1246
timestamp 1581449086
transform 1 0 1224 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1247
timestamp 1581449086
transform 1 0 612 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1248
timestamp 1581449086
transform 1 0 408 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_0
timestamp 1581449086
transform 1 0 52020 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1
timestamp 1581449086
transform 1 0 51408 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_2
timestamp 1581449086
transform 1 0 51204 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_3
timestamp 1581449086
transform 1 0 51000 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_4
timestamp 1581449086
transform 1 0 50592 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_5
timestamp 1581449086
transform 1 0 49572 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_6
timestamp 1581449086
transform 1 0 49368 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_7
timestamp 1581449086
transform 1 0 48756 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_8
timestamp 1581449086
transform 1 0 48348 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_9
timestamp 1581449086
transform 1 0 48144 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_10
timestamp 1581449086
transform 1 0 47940 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_11
timestamp 1581449086
transform 1 0 47124 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_12
timestamp 1581449086
transform 1 0 46920 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_13
timestamp 1581449086
transform 1 0 46104 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_14
timestamp 1581449086
transform 1 0 45084 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_15
timestamp 1581449086
transform 1 0 44676 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_16
timestamp 1581449086
transform 1 0 44268 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_17
timestamp 1581449086
transform 1 0 44064 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_18
timestamp 1581449086
transform 1 0 43044 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_19
timestamp 1581449086
transform 1 0 42840 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_20
timestamp 1581449086
transform 1 0 41412 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_21
timestamp 1581449086
transform 1 0 41208 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_22
timestamp 1581449086
transform 1 0 39780 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_23
timestamp 1581449086
transform 1 0 39576 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_24
timestamp 1581449086
transform 1 0 39372 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_25
timestamp 1581449086
transform 1 0 38964 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_26
timestamp 1581449086
transform 1 0 38556 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_27
timestamp 1581449086
transform 1 0 38148 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_28
timestamp 1581449086
transform 1 0 37944 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_29
timestamp 1581449086
transform 1 0 37536 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_30
timestamp 1581449086
transform 1 0 37332 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_31
timestamp 1581449086
transform 1 0 36924 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_32
timestamp 1581449086
transform 1 0 36312 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_33
timestamp 1581449086
transform 1 0 35700 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_34
timestamp 1581449086
transform 1 0 35496 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_35
timestamp 1581449086
transform 1 0 34884 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_36
timestamp 1581449086
transform 1 0 34680 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_37
timestamp 1581449086
transform 1 0 34476 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_38
timestamp 1581449086
transform 1 0 34272 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_39
timestamp 1581449086
transform 1 0 33864 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_40
timestamp 1581449086
transform 1 0 33252 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_41
timestamp 1581449086
transform 1 0 32844 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_42
timestamp 1581449086
transform 1 0 32640 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_43
timestamp 1581449086
transform 1 0 32232 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_44
timestamp 1581449086
transform 1 0 32028 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_45
timestamp 1581449086
transform 1 0 31620 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_46
timestamp 1581449086
transform 1 0 31212 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_47
timestamp 1581449086
transform 1 0 31008 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_48
timestamp 1581449086
transform 1 0 29988 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_49
timestamp 1581449086
transform 1 0 29376 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_50
timestamp 1581449086
transform 1 0 28968 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_51
timestamp 1581449086
transform 1 0 28356 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_52
timestamp 1581449086
transform 1 0 27744 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_53
timestamp 1581449086
transform 1 0 27540 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_54
timestamp 1581449086
transform 1 0 27132 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_55
timestamp 1581449086
transform 1 0 26724 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_56
timestamp 1581449086
transform 1 0 26520 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_57
timestamp 1581449086
transform 1 0 26316 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_58
timestamp 1581449086
transform 1 0 25500 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_59
timestamp 1581449086
transform 1 0 25296 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_60
timestamp 1581449086
transform 1 0 24888 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_61
timestamp 1581449086
transform 1 0 24276 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_62
timestamp 1581449086
transform 1 0 24072 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_63
timestamp 1581449086
transform 1 0 23868 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_64
timestamp 1581449086
transform 1 0 23256 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_65
timestamp 1581449086
transform 1 0 23052 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_66
timestamp 1581449086
transform 1 0 22644 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_67
timestamp 1581449086
transform 1 0 22440 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_68
timestamp 1581449086
transform 1 0 22236 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_69
timestamp 1581449086
transform 1 0 21624 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_70
timestamp 1581449086
transform 1 0 21012 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_71
timestamp 1581449086
transform 1 0 20604 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_72
timestamp 1581449086
transform 1 0 20196 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_73
timestamp 1581449086
transform 1 0 19788 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_74
timestamp 1581449086
transform 1 0 18564 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_75
timestamp 1581449086
transform 1 0 18360 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_76
timestamp 1581449086
transform 1 0 18156 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_77
timestamp 1581449086
transform 1 0 17952 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_78
timestamp 1581449086
transform 1 0 17340 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_79
timestamp 1581449086
transform 1 0 16932 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_80
timestamp 1581449086
transform 1 0 16728 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_81
timestamp 1581449086
transform 1 0 16320 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_82
timestamp 1581449086
transform 1 0 15504 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_83
timestamp 1581449086
transform 1 0 14892 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_84
timestamp 1581449086
transform 1 0 14688 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_85
timestamp 1581449086
transform 1 0 14484 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_86
timestamp 1581449086
transform 1 0 14076 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_87
timestamp 1581449086
transform 1 0 12852 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_88
timestamp 1581449086
transform 1 0 12648 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_89
timestamp 1581449086
transform 1 0 12444 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_90
timestamp 1581449086
transform 1 0 12240 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_91
timestamp 1581449086
transform 1 0 12036 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_92
timestamp 1581449086
transform 1 0 11832 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_93
timestamp 1581449086
transform 1 0 11628 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_94
timestamp 1581449086
transform 1 0 11424 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_95
timestamp 1581449086
transform 1 0 10812 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_96
timestamp 1581449086
transform 1 0 10608 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_97
timestamp 1581449086
transform 1 0 10404 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_98
timestamp 1581449086
transform 1 0 10200 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_99
timestamp 1581449086
transform 1 0 9996 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_100
timestamp 1581449086
transform 1 0 9792 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_101
timestamp 1581449086
transform 1 0 8976 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_102
timestamp 1581449086
transform 1 0 8364 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_103
timestamp 1581449086
transform 1 0 7956 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_104
timestamp 1581449086
transform 1 0 7548 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_105
timestamp 1581449086
transform 1 0 7344 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_106
timestamp 1581449086
transform 1 0 6936 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_107
timestamp 1581449086
transform 1 0 6528 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_108
timestamp 1581449086
transform 1 0 6324 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_109
timestamp 1581449086
transform 1 0 5916 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_110
timestamp 1581449086
transform 1 0 5508 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_111
timestamp 1581449086
transform 1 0 5304 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_112
timestamp 1581449086
transform 1 0 4692 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_113
timestamp 1581449086
transform 1 0 4080 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_114
timestamp 1581449086
transform 1 0 3876 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_115
timestamp 1581449086
transform 1 0 3672 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_116
timestamp 1581449086
transform 1 0 2856 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_117
timestamp 1581449086
transform 1 0 2652 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_118
timestamp 1581449086
transform 1 0 2448 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_119
timestamp 1581449086
transform 1 0 2244 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_120
timestamp 1581449086
transform 1 0 2040 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_121
timestamp 1581449086
transform 1 0 204 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_122
timestamp 1581449086
transform 1 0 0 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_123
timestamp 1581449086
transform 1 0 51612 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_124
timestamp 1581449086
transform 1 0 51000 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_125
timestamp 1581449086
transform 1 0 50796 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_126
timestamp 1581449086
transform 1 0 50592 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_127
timestamp 1581449086
transform 1 0 49572 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_128
timestamp 1581449086
transform 1 0 49368 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_129
timestamp 1581449086
transform 1 0 49164 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_130
timestamp 1581449086
transform 1 0 48756 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_131
timestamp 1581449086
transform 1 0 48348 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_132
timestamp 1581449086
transform 1 0 48144 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_133
timestamp 1581449086
transform 1 0 47532 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_134
timestamp 1581449086
transform 1 0 47124 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_135
timestamp 1581449086
transform 1 0 46512 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_136
timestamp 1581449086
transform 1 0 46308 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_137
timestamp 1581449086
transform 1 0 45696 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_138
timestamp 1581449086
transform 1 0 45288 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_139
timestamp 1581449086
transform 1 0 45084 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_140
timestamp 1581449086
transform 1 0 44472 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_141
timestamp 1581449086
transform 1 0 44268 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_142
timestamp 1581449086
transform 1 0 43656 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_143
timestamp 1581449086
transform 1 0 43452 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_144
timestamp 1581449086
transform 1 0 42840 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_145
timestamp 1581449086
transform 1 0 42636 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_146
timestamp 1581449086
transform 1 0 42432 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_147
timestamp 1581449086
transform 1 0 41616 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_148
timestamp 1581449086
transform 1 0 41412 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_149
timestamp 1581449086
transform 1 0 41004 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_150
timestamp 1581449086
transform 1 0 40800 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_151
timestamp 1581449086
transform 1 0 40392 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_152
timestamp 1581449086
transform 1 0 40188 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_153
timestamp 1581449086
transform 1 0 39576 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_154
timestamp 1581449086
transform 1 0 39372 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_155
timestamp 1581449086
transform 1 0 39168 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_156
timestamp 1581449086
transform 1 0 38760 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_157
timestamp 1581449086
transform 1 0 38556 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_158
timestamp 1581449086
transform 1 0 38352 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_159
timestamp 1581449086
transform 1 0 38148 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_160
timestamp 1581449086
transform 1 0 37740 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_161
timestamp 1581449086
transform 1 0 36720 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_162
timestamp 1581449086
transform 1 0 36516 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_163
timestamp 1581449086
transform 1 0 36108 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_164
timestamp 1581449086
transform 1 0 35904 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_165
timestamp 1581449086
transform 1 0 35496 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_166
timestamp 1581449086
transform 1 0 35292 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_167
timestamp 1581449086
transform 1 0 34272 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_168
timestamp 1581449086
transform 1 0 33048 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_169
timestamp 1581449086
transform 1 0 32640 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_170
timestamp 1581449086
transform 1 0 32436 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_171
timestamp 1581449086
transform 1 0 32232 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_172
timestamp 1581449086
transform 1 0 32028 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_173
timestamp 1581449086
transform 1 0 31824 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_174
timestamp 1581449086
transform 1 0 31212 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_175
timestamp 1581449086
transform 1 0 31008 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_176
timestamp 1581449086
transform 1 0 30600 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_177
timestamp 1581449086
transform 1 0 30192 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_178
timestamp 1581449086
transform 1 0 29376 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_179
timestamp 1581449086
transform 1 0 28764 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_180
timestamp 1581449086
transform 1 0 28560 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_181
timestamp 1581449086
transform 1 0 28356 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_182
timestamp 1581449086
transform 1 0 27540 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_183
timestamp 1581449086
transform 1 0 26928 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_184
timestamp 1581449086
transform 1 0 26520 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_185
timestamp 1581449086
transform 1 0 26316 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_186
timestamp 1581449086
transform 1 0 25908 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_187
timestamp 1581449086
transform 1 0 25704 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_188
timestamp 1581449086
transform 1 0 25500 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_189
timestamp 1581449086
transform 1 0 25296 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_190
timestamp 1581449086
transform 1 0 25092 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_191
timestamp 1581449086
transform 1 0 24888 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_192
timestamp 1581449086
transform 1 0 24480 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_193
timestamp 1581449086
transform 1 0 24072 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_194
timestamp 1581449086
transform 1 0 23868 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_195
timestamp 1581449086
transform 1 0 23664 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_196
timestamp 1581449086
transform 1 0 23460 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_197
timestamp 1581449086
transform 1 0 23256 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_198
timestamp 1581449086
transform 1 0 22848 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_199
timestamp 1581449086
transform 1 0 22236 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_200
timestamp 1581449086
transform 1 0 21828 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_201
timestamp 1581449086
transform 1 0 21624 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_202
timestamp 1581449086
transform 1 0 20196 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_203
timestamp 1581449086
transform 1 0 19788 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_204
timestamp 1581449086
transform 1 0 19584 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_205
timestamp 1581449086
transform 1 0 19380 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_206
timestamp 1581449086
transform 1 0 18360 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_207
timestamp 1581449086
transform 1 0 17952 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_208
timestamp 1581449086
transform 1 0 17544 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_209
timestamp 1581449086
transform 1 0 17340 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_210
timestamp 1581449086
transform 1 0 17136 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_211
timestamp 1581449086
transform 1 0 16728 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_212
timestamp 1581449086
transform 1 0 16116 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_213
timestamp 1581449086
transform 1 0 15912 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_214
timestamp 1581449086
transform 1 0 15504 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_215
timestamp 1581449086
transform 1 0 15300 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_216
timestamp 1581449086
transform 1 0 14892 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_217
timestamp 1581449086
transform 1 0 14688 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_218
timestamp 1581449086
transform 1 0 14484 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_219
timestamp 1581449086
transform 1 0 13872 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_220
timestamp 1581449086
transform 1 0 13464 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_221
timestamp 1581449086
transform 1 0 13260 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_222
timestamp 1581449086
transform 1 0 12852 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_223
timestamp 1581449086
transform 1 0 12444 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_224
timestamp 1581449086
transform 1 0 12036 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_225
timestamp 1581449086
transform 1 0 11628 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_226
timestamp 1581449086
transform 1 0 11220 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_227
timestamp 1581449086
transform 1 0 10608 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_228
timestamp 1581449086
transform 1 0 10404 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_229
timestamp 1581449086
transform 1 0 9792 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_230
timestamp 1581449086
transform 1 0 9588 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_231
timestamp 1581449086
transform 1 0 9384 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_232
timestamp 1581449086
transform 1 0 8976 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_233
timestamp 1581449086
transform 1 0 8160 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_234
timestamp 1581449086
transform 1 0 7140 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_235
timestamp 1581449086
transform 1 0 6936 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_236
timestamp 1581449086
transform 1 0 6324 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_237
timestamp 1581449086
transform 1 0 5916 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_238
timestamp 1581449086
transform 1 0 5304 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_239
timestamp 1581449086
transform 1 0 4488 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_240
timestamp 1581449086
transform 1 0 4284 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_241
timestamp 1581449086
transform 1 0 3468 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_242
timestamp 1581449086
transform 1 0 3264 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_243
timestamp 1581449086
transform 1 0 2448 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_244
timestamp 1581449086
transform 1 0 2244 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_245
timestamp 1581449086
transform 1 0 2040 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_246
timestamp 1581449086
transform 1 0 1836 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_247
timestamp 1581449086
transform 1 0 1632 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_248
timestamp 1581449086
transform 1 0 1428 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_249
timestamp 1581449086
transform 1 0 1224 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_250
timestamp 1581449086
transform 1 0 1020 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_251
timestamp 1581449086
transform 1 0 816 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_252
timestamp 1581449086
transform 1 0 612 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_253
timestamp 1581449086
transform 1 0 408 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_254
timestamp 1581449086
transform 1 0 204 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_255
timestamp 1581449086
transform 1 0 0 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_256
timestamp 1581449086
transform 1 0 52020 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_257
timestamp 1581449086
transform 1 0 51612 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_258
timestamp 1581449086
transform 1 0 51000 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_259
timestamp 1581449086
transform 1 0 50388 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_260
timestamp 1581449086
transform 1 0 50184 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_261
timestamp 1581449086
transform 1 0 49980 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_262
timestamp 1581449086
transform 1 0 49776 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_263
timestamp 1581449086
transform 1 0 49368 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_264
timestamp 1581449086
transform 1 0 48960 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_265
timestamp 1581449086
transform 1 0 48756 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_266
timestamp 1581449086
transform 1 0 48144 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_267
timestamp 1581449086
transform 1 0 47940 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_268
timestamp 1581449086
transform 1 0 47736 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_269
timestamp 1581449086
transform 1 0 47532 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_270
timestamp 1581449086
transform 1 0 47328 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_271
timestamp 1581449086
transform 1 0 47124 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_272
timestamp 1581449086
transform 1 0 46920 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_273
timestamp 1581449086
transform 1 0 46716 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_274
timestamp 1581449086
transform 1 0 46308 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_275
timestamp 1581449086
transform 1 0 46104 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_276
timestamp 1581449086
transform 1 0 45696 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_277
timestamp 1581449086
transform 1 0 45288 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_278
timestamp 1581449086
transform 1 0 45084 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_279
timestamp 1581449086
transform 1 0 44676 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_280
timestamp 1581449086
transform 1 0 44268 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_281
timestamp 1581449086
transform 1 0 44064 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_282
timestamp 1581449086
transform 1 0 43656 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_283
timestamp 1581449086
transform 1 0 43248 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_284
timestamp 1581449086
transform 1 0 42636 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_285
timestamp 1581449086
transform 1 0 42024 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_286
timestamp 1581449086
transform 1 0 41820 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_287
timestamp 1581449086
transform 1 0 41616 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_288
timestamp 1581449086
transform 1 0 41412 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_289
timestamp 1581449086
transform 1 0 40800 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_290
timestamp 1581449086
transform 1 0 40596 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_291
timestamp 1581449086
transform 1 0 40188 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_292
timestamp 1581449086
transform 1 0 39984 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_293
timestamp 1581449086
transform 1 0 39576 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_294
timestamp 1581449086
transform 1 0 39372 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_295
timestamp 1581449086
transform 1 0 38964 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_296
timestamp 1581449086
transform 1 0 38556 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_297
timestamp 1581449086
transform 1 0 38352 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_298
timestamp 1581449086
transform 1 0 37740 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_299
timestamp 1581449086
transform 1 0 37536 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_300
timestamp 1581449086
transform 1 0 37332 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_301
timestamp 1581449086
transform 1 0 37128 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_302
timestamp 1581449086
transform 1 0 36720 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_303
timestamp 1581449086
transform 1 0 36516 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_304
timestamp 1581449086
transform 1 0 35904 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_305
timestamp 1581449086
transform 1 0 35700 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_306
timestamp 1581449086
transform 1 0 35088 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_307
timestamp 1581449086
transform 1 0 34884 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_308
timestamp 1581449086
transform 1 0 34680 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_309
timestamp 1581449086
transform 1 0 34272 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_310
timestamp 1581449086
transform 1 0 34068 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_311
timestamp 1581449086
transform 1 0 33864 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_312
timestamp 1581449086
transform 1 0 33660 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_313
timestamp 1581449086
transform 1 0 33252 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_314
timestamp 1581449086
transform 1 0 32844 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_315
timestamp 1581449086
transform 1 0 32436 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_316
timestamp 1581449086
transform 1 0 32028 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_317
timestamp 1581449086
transform 1 0 31824 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_318
timestamp 1581449086
transform 1 0 31416 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_319
timestamp 1581449086
transform 1 0 31212 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_320
timestamp 1581449086
transform 1 0 31008 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_321
timestamp 1581449086
transform 1 0 30396 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_322
timestamp 1581449086
transform 1 0 29988 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_323
timestamp 1581449086
transform 1 0 29784 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_324
timestamp 1581449086
transform 1 0 29172 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_325
timestamp 1581449086
transform 1 0 28968 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_326
timestamp 1581449086
transform 1 0 28764 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_327
timestamp 1581449086
transform 1 0 28152 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_328
timestamp 1581449086
transform 1 0 27336 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_329
timestamp 1581449086
transform 1 0 27132 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_330
timestamp 1581449086
transform 1 0 26724 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_331
timestamp 1581449086
transform 1 0 26316 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_332
timestamp 1581449086
transform 1 0 25908 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_333
timestamp 1581449086
transform 1 0 25704 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_334
timestamp 1581449086
transform 1 0 25296 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_335
timestamp 1581449086
transform 1 0 25092 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_336
timestamp 1581449086
transform 1 0 24684 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_337
timestamp 1581449086
transform 1 0 23868 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_338
timestamp 1581449086
transform 1 0 23460 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_339
timestamp 1581449086
transform 1 0 22644 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_340
timestamp 1581449086
transform 1 0 22236 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_341
timestamp 1581449086
transform 1 0 22032 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_342
timestamp 1581449086
transform 1 0 21624 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_343
timestamp 1581449086
transform 1 0 21420 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_344
timestamp 1581449086
transform 1 0 20400 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_345
timestamp 1581449086
transform 1 0 19380 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_346
timestamp 1581449086
transform 1 0 19176 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_347
timestamp 1581449086
transform 1 0 18564 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_348
timestamp 1581449086
transform 1 0 18360 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_349
timestamp 1581449086
transform 1 0 17544 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_350
timestamp 1581449086
transform 1 0 17340 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_351
timestamp 1581449086
transform 1 0 17136 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_352
timestamp 1581449086
transform 1 0 16728 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_353
timestamp 1581449086
transform 1 0 16524 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_354
timestamp 1581449086
transform 1 0 15912 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_355
timestamp 1581449086
transform 1 0 15708 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_356
timestamp 1581449086
transform 1 0 15504 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_357
timestamp 1581449086
transform 1 0 14892 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_358
timestamp 1581449086
transform 1 0 14688 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_359
timestamp 1581449086
transform 1 0 14484 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_360
timestamp 1581449086
transform 1 0 14280 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_361
timestamp 1581449086
transform 1 0 13668 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_362
timestamp 1581449086
transform 1 0 13464 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_363
timestamp 1581449086
transform 1 0 13260 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_364
timestamp 1581449086
transform 1 0 12852 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_365
timestamp 1581449086
transform 1 0 12648 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_366
timestamp 1581449086
transform 1 0 12444 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_367
timestamp 1581449086
transform 1 0 11832 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_368
timestamp 1581449086
transform 1 0 11628 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_369
timestamp 1581449086
transform 1 0 11424 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_370
timestamp 1581449086
transform 1 0 11220 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_371
timestamp 1581449086
transform 1 0 11016 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_372
timestamp 1581449086
transform 1 0 10608 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_373
timestamp 1581449086
transform 1 0 9996 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_374
timestamp 1581449086
transform 1 0 9588 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_375
timestamp 1581449086
transform 1 0 8976 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_376
timestamp 1581449086
transform 1 0 8568 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_377
timestamp 1581449086
transform 1 0 8364 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_378
timestamp 1581449086
transform 1 0 8160 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_379
timestamp 1581449086
transform 1 0 7956 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_380
timestamp 1581449086
transform 1 0 7752 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_381
timestamp 1581449086
transform 1 0 7548 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_382
timestamp 1581449086
transform 1 0 7344 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_383
timestamp 1581449086
transform 1 0 7140 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_384
timestamp 1581449086
transform 1 0 6936 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_385
timestamp 1581449086
transform 1 0 6528 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_386
timestamp 1581449086
transform 1 0 5508 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_387
timestamp 1581449086
transform 1 0 5304 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_388
timestamp 1581449086
transform 1 0 5100 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_389
timestamp 1581449086
transform 1 0 4896 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_390
timestamp 1581449086
transform 1 0 4692 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_391
timestamp 1581449086
transform 1 0 4284 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_392
timestamp 1581449086
transform 1 0 4080 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_393
timestamp 1581449086
transform 1 0 3876 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_394
timestamp 1581449086
transform 1 0 3672 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_395
timestamp 1581449086
transform 1 0 3060 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_396
timestamp 1581449086
transform 1 0 1836 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_397
timestamp 1581449086
transform 1 0 1632 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_398
timestamp 1581449086
transform 1 0 1428 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_399
timestamp 1581449086
transform 1 0 51816 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_400
timestamp 1581449086
transform 1 0 51408 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_401
timestamp 1581449086
transform 1 0 51000 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_402
timestamp 1581449086
transform 1 0 50796 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_403
timestamp 1581449086
transform 1 0 50388 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_404
timestamp 1581449086
transform 1 0 49776 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_405
timestamp 1581449086
transform 1 0 49368 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_406
timestamp 1581449086
transform 1 0 49164 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_407
timestamp 1581449086
transform 1 0 48960 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_408
timestamp 1581449086
transform 1 0 48348 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_409
timestamp 1581449086
transform 1 0 47940 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_410
timestamp 1581449086
transform 1 0 47532 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_411
timestamp 1581449086
transform 1 0 47124 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_412
timestamp 1581449086
transform 1 0 46512 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_413
timestamp 1581449086
transform 1 0 46308 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_414
timestamp 1581449086
transform 1 0 45696 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_415
timestamp 1581449086
transform 1 0 45492 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_416
timestamp 1581449086
transform 1 0 45288 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_417
timestamp 1581449086
transform 1 0 44064 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_418
timestamp 1581449086
transform 1 0 43860 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_419
timestamp 1581449086
transform 1 0 43248 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_420
timestamp 1581449086
transform 1 0 43044 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_421
timestamp 1581449086
transform 1 0 42432 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_422
timestamp 1581449086
transform 1 0 42228 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_423
timestamp 1581449086
transform 1 0 42024 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_424
timestamp 1581449086
transform 1 0 41820 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_425
timestamp 1581449086
transform 1 0 41412 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_426
timestamp 1581449086
transform 1 0 41004 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_427
timestamp 1581449086
transform 1 0 40800 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_428
timestamp 1581449086
transform 1 0 40392 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_429
timestamp 1581449086
transform 1 0 39984 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_430
timestamp 1581449086
transform 1 0 39780 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_431
timestamp 1581449086
transform 1 0 39372 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_432
timestamp 1581449086
transform 1 0 38964 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_433
timestamp 1581449086
transform 1 0 38556 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_434
timestamp 1581449086
transform 1 0 37536 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_435
timestamp 1581449086
transform 1 0 37332 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_436
timestamp 1581449086
transform 1 0 37128 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_437
timestamp 1581449086
transform 1 0 36516 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_438
timestamp 1581449086
transform 1 0 36312 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_439
timestamp 1581449086
transform 1 0 36108 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_440
timestamp 1581449086
transform 1 0 35496 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_441
timestamp 1581449086
transform 1 0 35292 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_442
timestamp 1581449086
transform 1 0 35088 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_443
timestamp 1581449086
transform 1 0 34476 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_444
timestamp 1581449086
transform 1 0 34272 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_445
timestamp 1581449086
transform 1 0 33456 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_446
timestamp 1581449086
transform 1 0 32844 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_447
timestamp 1581449086
transform 1 0 32436 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_448
timestamp 1581449086
transform 1 0 32232 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_449
timestamp 1581449086
transform 1 0 32028 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_450
timestamp 1581449086
transform 1 0 31620 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_451
timestamp 1581449086
transform 1 0 31416 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_452
timestamp 1581449086
transform 1 0 31212 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_453
timestamp 1581449086
transform 1 0 31008 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_454
timestamp 1581449086
transform 1 0 30600 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_455
timestamp 1581449086
transform 1 0 30396 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_456
timestamp 1581449086
transform 1 0 29988 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_457
timestamp 1581449086
transform 1 0 29376 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_458
timestamp 1581449086
transform 1 0 29172 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_459
timestamp 1581449086
transform 1 0 28764 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_460
timestamp 1581449086
transform 1 0 28356 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_461
timestamp 1581449086
transform 1 0 27948 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_462
timestamp 1581449086
transform 1 0 27744 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_463
timestamp 1581449086
transform 1 0 27540 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_464
timestamp 1581449086
transform 1 0 27132 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_465
timestamp 1581449086
transform 1 0 26928 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_466
timestamp 1581449086
transform 1 0 26724 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_467
timestamp 1581449086
transform 1 0 26520 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_468
timestamp 1581449086
transform 1 0 26316 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_469
timestamp 1581449086
transform 1 0 26112 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_470
timestamp 1581449086
transform 1 0 25908 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_471
timestamp 1581449086
transform 1 0 25704 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_472
timestamp 1581449086
transform 1 0 25500 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_473
timestamp 1581449086
transform 1 0 25296 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_474
timestamp 1581449086
transform 1 0 25092 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_475
timestamp 1581449086
transform 1 0 24888 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_476
timestamp 1581449086
transform 1 0 23460 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_477
timestamp 1581449086
transform 1 0 23256 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_478
timestamp 1581449086
transform 1 0 22644 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_479
timestamp 1581449086
transform 1 0 22440 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_480
timestamp 1581449086
transform 1 0 22236 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_481
timestamp 1581449086
transform 1 0 22032 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_482
timestamp 1581449086
transform 1 0 21828 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_483
timestamp 1581449086
transform 1 0 21420 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_484
timestamp 1581449086
transform 1 0 21012 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_485
timestamp 1581449086
transform 1 0 20808 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_486
timestamp 1581449086
transform 1 0 19584 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_487
timestamp 1581449086
transform 1 0 19176 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_488
timestamp 1581449086
transform 1 0 18972 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_489
timestamp 1581449086
transform 1 0 18768 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_490
timestamp 1581449086
transform 1 0 18360 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_491
timestamp 1581449086
transform 1 0 17544 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_492
timestamp 1581449086
transform 1 0 17136 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_493
timestamp 1581449086
transform 1 0 16524 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_494
timestamp 1581449086
transform 1 0 15504 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_495
timestamp 1581449086
transform 1 0 15300 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_496
timestamp 1581449086
transform 1 0 15096 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_497
timestamp 1581449086
transform 1 0 14892 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_498
timestamp 1581449086
transform 1 0 14688 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_499
timestamp 1581449086
transform 1 0 14484 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_500
timestamp 1581449086
transform 1 0 14076 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_501
timestamp 1581449086
transform 1 0 13872 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_502
timestamp 1581449086
transform 1 0 13668 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_503
timestamp 1581449086
transform 1 0 13464 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_504
timestamp 1581449086
transform 1 0 13260 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_505
timestamp 1581449086
transform 1 0 12852 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_506
timestamp 1581449086
transform 1 0 12444 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_507
timestamp 1581449086
transform 1 0 11628 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_508
timestamp 1581449086
transform 1 0 11016 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_509
timestamp 1581449086
transform 1 0 10608 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_510
timestamp 1581449086
transform 1 0 10200 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_511
timestamp 1581449086
transform 1 0 9588 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_512
timestamp 1581449086
transform 1 0 9384 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_513
timestamp 1581449086
transform 1 0 8772 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_514
timestamp 1581449086
transform 1 0 7956 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_515
timestamp 1581449086
transform 1 0 7752 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_516
timestamp 1581449086
transform 1 0 7548 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_517
timestamp 1581449086
transform 1 0 7344 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_518
timestamp 1581449086
transform 1 0 7140 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_519
timestamp 1581449086
transform 1 0 6528 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_520
timestamp 1581449086
transform 1 0 6120 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_521
timestamp 1581449086
transform 1 0 5712 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_522
timestamp 1581449086
transform 1 0 5304 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_523
timestamp 1581449086
transform 1 0 5100 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_524
timestamp 1581449086
transform 1 0 4896 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_525
timestamp 1581449086
transform 1 0 4692 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_526
timestamp 1581449086
transform 1 0 4488 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_527
timestamp 1581449086
transform 1 0 3876 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_528
timestamp 1581449086
transform 1 0 3672 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_529
timestamp 1581449086
transform 1 0 3060 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_530
timestamp 1581449086
transform 1 0 2856 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_531
timestamp 1581449086
transform 1 0 1836 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_532
timestamp 1581449086
transform 1 0 1632 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_533
timestamp 1581449086
transform 1 0 1020 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_534
timestamp 1581449086
transform 1 0 816 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_535
timestamp 1581449086
transform 1 0 612 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_536
timestamp 1581449086
transform 1 0 408 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_537
timestamp 1581449086
transform 1 0 204 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_538
timestamp 1581449086
transform 1 0 0 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_539
timestamp 1581449086
transform 1 0 51000 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_540
timestamp 1581449086
transform 1 0 50592 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_541
timestamp 1581449086
transform 1 0 50184 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_542
timestamp 1581449086
transform 1 0 49368 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_543
timestamp 1581449086
transform 1 0 49164 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_544
timestamp 1581449086
transform 1 0 48552 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_545
timestamp 1581449086
transform 1 0 48144 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_546
timestamp 1581449086
transform 1 0 47736 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_547
timestamp 1581449086
transform 1 0 47328 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_548
timestamp 1581449086
transform 1 0 47124 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_549
timestamp 1581449086
transform 1 0 46920 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_550
timestamp 1581449086
transform 1 0 46716 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_551
timestamp 1581449086
transform 1 0 46512 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_552
timestamp 1581449086
transform 1 0 46308 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_553
timestamp 1581449086
transform 1 0 45696 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_554
timestamp 1581449086
transform 1 0 45492 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_555
timestamp 1581449086
transform 1 0 45084 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_556
timestamp 1581449086
transform 1 0 44676 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_557
timestamp 1581449086
transform 1 0 44472 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_558
timestamp 1581449086
transform 1 0 44268 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_559
timestamp 1581449086
transform 1 0 43656 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_560
timestamp 1581449086
transform 1 0 43452 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_561
timestamp 1581449086
transform 1 0 43044 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_562
timestamp 1581449086
transform 1 0 42840 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_563
timestamp 1581449086
transform 1 0 42432 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_564
timestamp 1581449086
transform 1 0 40596 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_565
timestamp 1581449086
transform 1 0 40392 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_566
timestamp 1581449086
transform 1 0 40188 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_567
timestamp 1581449086
transform 1 0 39372 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_568
timestamp 1581449086
transform 1 0 39168 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_569
timestamp 1581449086
transform 1 0 37740 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_570
timestamp 1581449086
transform 1 0 37332 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_571
timestamp 1581449086
transform 1 0 36924 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_572
timestamp 1581449086
transform 1 0 35904 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_573
timestamp 1581449086
transform 1 0 35700 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_574
timestamp 1581449086
transform 1 0 35496 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_575
timestamp 1581449086
transform 1 0 35292 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_576
timestamp 1581449086
transform 1 0 35088 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_577
timestamp 1581449086
transform 1 0 34272 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_578
timestamp 1581449086
transform 1 0 33864 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_579
timestamp 1581449086
transform 1 0 33660 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_580
timestamp 1581449086
transform 1 0 33048 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_581
timestamp 1581449086
transform 1 0 32844 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_582
timestamp 1581449086
transform 1 0 32640 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_583
timestamp 1581449086
transform 1 0 32436 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_584
timestamp 1581449086
transform 1 0 32232 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_585
timestamp 1581449086
transform 1 0 31824 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_586
timestamp 1581449086
transform 1 0 31416 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_587
timestamp 1581449086
transform 1 0 31212 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_588
timestamp 1581449086
transform 1 0 30396 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_589
timestamp 1581449086
transform 1 0 30192 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_590
timestamp 1581449086
transform 1 0 29580 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_591
timestamp 1581449086
transform 1 0 29376 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_592
timestamp 1581449086
transform 1 0 29172 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_593
timestamp 1581449086
transform 1 0 28764 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_594
timestamp 1581449086
transform 1 0 28560 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_595
timestamp 1581449086
transform 1 0 28152 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_596
timestamp 1581449086
transform 1 0 27540 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_597
timestamp 1581449086
transform 1 0 27336 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_598
timestamp 1581449086
transform 1 0 26928 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_599
timestamp 1581449086
transform 1 0 26724 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_600
timestamp 1581449086
transform 1 0 26520 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_601
timestamp 1581449086
transform 1 0 26112 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_602
timestamp 1581449086
transform 1 0 25704 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_603
timestamp 1581449086
transform 1 0 25296 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_604
timestamp 1581449086
transform 1 0 24480 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_605
timestamp 1581449086
transform 1 0 24276 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_606
timestamp 1581449086
transform 1 0 23664 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_607
timestamp 1581449086
transform 1 0 23460 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_608
timestamp 1581449086
transform 1 0 23052 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_609
timestamp 1581449086
transform 1 0 22644 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_610
timestamp 1581449086
transform 1 0 22440 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_611
timestamp 1581449086
transform 1 0 22032 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_612
timestamp 1581449086
transform 1 0 21828 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_613
timestamp 1581449086
transform 1 0 21624 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_614
timestamp 1581449086
transform 1 0 21420 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_615
timestamp 1581449086
transform 1 0 20604 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_616
timestamp 1581449086
transform 1 0 20400 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_617
timestamp 1581449086
transform 1 0 19992 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_618
timestamp 1581449086
transform 1 0 19788 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_619
timestamp 1581449086
transform 1 0 19380 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_620
timestamp 1581449086
transform 1 0 19176 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_621
timestamp 1581449086
transform 1 0 18972 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_622
timestamp 1581449086
transform 1 0 18768 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_623
timestamp 1581449086
transform 1 0 18360 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_624
timestamp 1581449086
transform 1 0 17544 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_625
timestamp 1581449086
transform 1 0 16932 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_626
timestamp 1581449086
transform 1 0 16728 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_627
timestamp 1581449086
transform 1 0 16116 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_628
timestamp 1581449086
transform 1 0 15708 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_629
timestamp 1581449086
transform 1 0 15096 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_630
timestamp 1581449086
transform 1 0 14892 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_631
timestamp 1581449086
transform 1 0 14688 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_632
timestamp 1581449086
transform 1 0 14484 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_633
timestamp 1581449086
transform 1 0 13668 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_634
timestamp 1581449086
transform 1 0 13464 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_635
timestamp 1581449086
transform 1 0 13260 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_636
timestamp 1581449086
transform 1 0 13056 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_637
timestamp 1581449086
transform 1 0 12852 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_638
timestamp 1581449086
transform 1 0 12648 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_639
timestamp 1581449086
transform 1 0 12240 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_640
timestamp 1581449086
transform 1 0 11832 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_641
timestamp 1581449086
transform 1 0 11628 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_642
timestamp 1581449086
transform 1 0 11424 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_643
timestamp 1581449086
transform 1 0 11220 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_644
timestamp 1581449086
transform 1 0 10812 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_645
timestamp 1581449086
transform 1 0 10200 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_646
timestamp 1581449086
transform 1 0 9996 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_647
timestamp 1581449086
transform 1 0 9792 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_648
timestamp 1581449086
transform 1 0 8568 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_649
timestamp 1581449086
transform 1 0 8364 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_650
timestamp 1581449086
transform 1 0 8160 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_651
timestamp 1581449086
transform 1 0 7956 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_652
timestamp 1581449086
transform 1 0 7752 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_653
timestamp 1581449086
transform 1 0 7548 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_654
timestamp 1581449086
transform 1 0 7344 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_655
timestamp 1581449086
transform 1 0 6936 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_656
timestamp 1581449086
transform 1 0 6120 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_657
timestamp 1581449086
transform 1 0 5712 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_658
timestamp 1581449086
transform 1 0 5100 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_659
timestamp 1581449086
transform 1 0 4692 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_660
timestamp 1581449086
transform 1 0 4488 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_661
timestamp 1581449086
transform 1 0 4284 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_662
timestamp 1581449086
transform 1 0 4080 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_663
timestamp 1581449086
transform 1 0 3264 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_664
timestamp 1581449086
transform 1 0 3060 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_665
timestamp 1581449086
transform 1 0 2856 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_666
timestamp 1581449086
transform 1 0 2244 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_667
timestamp 1581449086
transform 1 0 2040 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_668
timestamp 1581449086
transform 1 0 1836 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_669
timestamp 1581449086
transform 1 0 1632 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_670
timestamp 1581449086
transform 1 0 1428 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_671
timestamp 1581449086
transform 1 0 1224 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_672
timestamp 1581449086
transform 1 0 52020 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_673
timestamp 1581449086
transform 1 0 51816 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_674
timestamp 1581449086
transform 1 0 51612 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_675
timestamp 1581449086
transform 1 0 51204 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_676
timestamp 1581449086
transform 1 0 51000 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_677
timestamp 1581449086
transform 1 0 50796 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_678
timestamp 1581449086
transform 1 0 50184 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_679
timestamp 1581449086
transform 1 0 49572 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_680
timestamp 1581449086
transform 1 0 48960 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_681
timestamp 1581449086
transform 1 0 48756 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_682
timestamp 1581449086
transform 1 0 48348 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_683
timestamp 1581449086
transform 1 0 47328 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_684
timestamp 1581449086
transform 1 0 46104 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_685
timestamp 1581449086
transform 1 0 45900 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_686
timestamp 1581449086
transform 1 0 45696 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_687
timestamp 1581449086
transform 1 0 45084 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_688
timestamp 1581449086
transform 1 0 44880 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_689
timestamp 1581449086
transform 1 0 44676 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_690
timestamp 1581449086
transform 1 0 44472 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_691
timestamp 1581449086
transform 1 0 44268 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_692
timestamp 1581449086
transform 1 0 44064 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_693
timestamp 1581449086
transform 1 0 43860 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_694
timestamp 1581449086
transform 1 0 43656 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_695
timestamp 1581449086
transform 1 0 43044 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_696
timestamp 1581449086
transform 1 0 42840 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_697
timestamp 1581449086
transform 1 0 42636 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_698
timestamp 1581449086
transform 1 0 42432 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_699
timestamp 1581449086
transform 1 0 41820 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_700
timestamp 1581449086
transform 1 0 41004 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_701
timestamp 1581449086
transform 1 0 39984 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_702
timestamp 1581449086
transform 1 0 38964 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_703
timestamp 1581449086
transform 1 0 38556 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_704
timestamp 1581449086
transform 1 0 38352 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_705
timestamp 1581449086
transform 1 0 37332 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_706
timestamp 1581449086
transform 1 0 37128 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_707
timestamp 1581449086
transform 1 0 36924 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_708
timestamp 1581449086
transform 1 0 36720 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_709
timestamp 1581449086
transform 1 0 36516 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_710
timestamp 1581449086
transform 1 0 36312 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_711
timestamp 1581449086
transform 1 0 35904 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_712
timestamp 1581449086
transform 1 0 35700 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_713
timestamp 1581449086
transform 1 0 35496 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_714
timestamp 1581449086
transform 1 0 34884 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_715
timestamp 1581449086
transform 1 0 34272 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_716
timestamp 1581449086
transform 1 0 33660 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_717
timestamp 1581449086
transform 1 0 33252 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_718
timestamp 1581449086
transform 1 0 32844 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_719
timestamp 1581449086
transform 1 0 32436 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_720
timestamp 1581449086
transform 1 0 32232 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_721
timestamp 1581449086
transform 1 0 32028 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_722
timestamp 1581449086
transform 1 0 31824 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_723
timestamp 1581449086
transform 1 0 31620 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_724
timestamp 1581449086
transform 1 0 31212 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_725
timestamp 1581449086
transform 1 0 31008 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_726
timestamp 1581449086
transform 1 0 30804 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_727
timestamp 1581449086
transform 1 0 30396 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_728
timestamp 1581449086
transform 1 0 29784 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_729
timestamp 1581449086
transform 1 0 29580 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_730
timestamp 1581449086
transform 1 0 29172 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_731
timestamp 1581449086
transform 1 0 28968 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_732
timestamp 1581449086
transform 1 0 28764 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_733
timestamp 1581449086
transform 1 0 28560 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_734
timestamp 1581449086
transform 1 0 28356 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_735
timestamp 1581449086
transform 1 0 28152 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_736
timestamp 1581449086
transform 1 0 26928 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_737
timestamp 1581449086
transform 1 0 26316 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_738
timestamp 1581449086
transform 1 0 26112 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_739
timestamp 1581449086
transform 1 0 25704 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_740
timestamp 1581449086
transform 1 0 25500 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_741
timestamp 1581449086
transform 1 0 25092 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_742
timestamp 1581449086
transform 1 0 24684 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_743
timestamp 1581449086
transform 1 0 24276 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_744
timestamp 1581449086
transform 1 0 24072 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_745
timestamp 1581449086
transform 1 0 23868 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_746
timestamp 1581449086
transform 1 0 23664 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_747
timestamp 1581449086
transform 1 0 23460 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_748
timestamp 1581449086
transform 1 0 23256 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_749
timestamp 1581449086
transform 1 0 22644 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_750
timestamp 1581449086
transform 1 0 22440 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_751
timestamp 1581449086
transform 1 0 22032 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_752
timestamp 1581449086
transform 1 0 21624 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_753
timestamp 1581449086
transform 1 0 21216 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_754
timestamp 1581449086
transform 1 0 20808 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_755
timestamp 1581449086
transform 1 0 20604 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_756
timestamp 1581449086
transform 1 0 19992 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_757
timestamp 1581449086
transform 1 0 18768 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_758
timestamp 1581449086
transform 1 0 18564 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_759
timestamp 1581449086
transform 1 0 18360 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_760
timestamp 1581449086
transform 1 0 16932 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_761
timestamp 1581449086
transform 1 0 16728 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_762
timestamp 1581449086
transform 1 0 16320 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_763
timestamp 1581449086
transform 1 0 15912 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_764
timestamp 1581449086
transform 1 0 15300 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_765
timestamp 1581449086
transform 1 0 14892 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_766
timestamp 1581449086
transform 1 0 14688 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_767
timestamp 1581449086
transform 1 0 14076 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_768
timestamp 1581449086
transform 1 0 13668 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_769
timestamp 1581449086
transform 1 0 12852 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_770
timestamp 1581449086
transform 1 0 12648 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_771
timestamp 1581449086
transform 1 0 12444 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_772
timestamp 1581449086
transform 1 0 12036 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_773
timestamp 1581449086
transform 1 0 11424 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_774
timestamp 1581449086
transform 1 0 11016 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_775
timestamp 1581449086
transform 1 0 10608 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_776
timestamp 1581449086
transform 1 0 10404 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_777
timestamp 1581449086
transform 1 0 9792 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_778
timestamp 1581449086
transform 1 0 9180 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_779
timestamp 1581449086
transform 1 0 7956 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_780
timestamp 1581449086
transform 1 0 7140 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_781
timestamp 1581449086
transform 1 0 6528 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_782
timestamp 1581449086
transform 1 0 5916 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_783
timestamp 1581449086
transform 1 0 5712 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_784
timestamp 1581449086
transform 1 0 5508 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_785
timestamp 1581449086
transform 1 0 5304 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_786
timestamp 1581449086
transform 1 0 5100 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_787
timestamp 1581449086
transform 1 0 4896 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_788
timestamp 1581449086
transform 1 0 4488 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_789
timestamp 1581449086
transform 1 0 4284 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_790
timestamp 1581449086
transform 1 0 3672 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_791
timestamp 1581449086
transform 1 0 2448 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_792
timestamp 1581449086
transform 1 0 2244 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_793
timestamp 1581449086
transform 1 0 2040 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_794
timestamp 1581449086
transform 1 0 1428 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_795
timestamp 1581449086
transform 1 0 1224 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_796
timestamp 1581449086
transform 1 0 1020 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_797
timestamp 1581449086
transform 1 0 816 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_798
timestamp 1581449086
transform 1 0 612 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_799
timestamp 1581449086
transform 1 0 408 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_800
timestamp 1581449086
transform 1 0 52020 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_801
timestamp 1581449086
transform 1 0 51612 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_802
timestamp 1581449086
transform 1 0 51408 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_803
timestamp 1581449086
transform 1 0 51000 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_804
timestamp 1581449086
transform 1 0 50592 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_805
timestamp 1581449086
transform 1 0 50388 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_806
timestamp 1581449086
transform 1 0 49776 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_807
timestamp 1581449086
transform 1 0 49164 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_808
timestamp 1581449086
transform 1 0 48960 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_809
timestamp 1581449086
transform 1 0 47940 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_810
timestamp 1581449086
transform 1 0 47532 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_811
timestamp 1581449086
transform 1 0 47328 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_812
timestamp 1581449086
transform 1 0 47124 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_813
timestamp 1581449086
transform 1 0 46920 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_814
timestamp 1581449086
transform 1 0 46512 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_815
timestamp 1581449086
transform 1 0 46308 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_816
timestamp 1581449086
transform 1 0 45900 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_817
timestamp 1581449086
transform 1 0 45288 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_818
timestamp 1581449086
transform 1 0 44676 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_819
timestamp 1581449086
transform 1 0 44268 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_820
timestamp 1581449086
transform 1 0 43044 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_821
timestamp 1581449086
transform 1 0 42636 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_822
timestamp 1581449086
transform 1 0 42432 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_823
timestamp 1581449086
transform 1 0 42024 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_824
timestamp 1581449086
transform 1 0 41208 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_825
timestamp 1581449086
transform 1 0 41004 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_826
timestamp 1581449086
transform 1 0 40800 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_827
timestamp 1581449086
transform 1 0 40596 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_828
timestamp 1581449086
transform 1 0 39984 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_829
timestamp 1581449086
transform 1 0 39372 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_830
timestamp 1581449086
transform 1 0 38760 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_831
timestamp 1581449086
transform 1 0 37536 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_832
timestamp 1581449086
transform 1 0 37332 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_833
timestamp 1581449086
transform 1 0 36924 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_834
timestamp 1581449086
transform 1 0 36720 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_835
timestamp 1581449086
transform 1 0 36516 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_836
timestamp 1581449086
transform 1 0 36312 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_837
timestamp 1581449086
transform 1 0 35700 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_838
timestamp 1581449086
transform 1 0 35292 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_839
timestamp 1581449086
transform 1 0 34476 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_840
timestamp 1581449086
transform 1 0 34272 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_841
timestamp 1581449086
transform 1 0 34068 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_842
timestamp 1581449086
transform 1 0 33864 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_843
timestamp 1581449086
transform 1 0 33660 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_844
timestamp 1581449086
transform 1 0 33048 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_845
timestamp 1581449086
transform 1 0 32232 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_846
timestamp 1581449086
transform 1 0 31416 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_847
timestamp 1581449086
transform 1 0 31008 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_848
timestamp 1581449086
transform 1 0 30600 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_849
timestamp 1581449086
transform 1 0 30192 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_850
timestamp 1581449086
transform 1 0 29784 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_851
timestamp 1581449086
transform 1 0 29580 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_852
timestamp 1581449086
transform 1 0 28968 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_853
timestamp 1581449086
transform 1 0 28764 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_854
timestamp 1581449086
transform 1 0 28152 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_855
timestamp 1581449086
transform 1 0 27744 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_856
timestamp 1581449086
transform 1 0 27336 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_857
timestamp 1581449086
transform 1 0 26928 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_858
timestamp 1581449086
transform 1 0 26724 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_859
timestamp 1581449086
transform 1 0 26316 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_860
timestamp 1581449086
transform 1 0 25704 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_861
timestamp 1581449086
transform 1 0 25500 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_862
timestamp 1581449086
transform 1 0 25296 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_863
timestamp 1581449086
transform 1 0 25092 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_864
timestamp 1581449086
transform 1 0 24072 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_865
timestamp 1581449086
transform 1 0 23460 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_866
timestamp 1581449086
transform 1 0 23256 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_867
timestamp 1581449086
transform 1 0 22644 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_868
timestamp 1581449086
transform 1 0 21624 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_869
timestamp 1581449086
transform 1 0 21420 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_870
timestamp 1581449086
transform 1 0 19992 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_871
timestamp 1581449086
transform 1 0 19788 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_872
timestamp 1581449086
transform 1 0 19584 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_873
timestamp 1581449086
transform 1 0 18564 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_874
timestamp 1581449086
transform 1 0 18156 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_875
timestamp 1581449086
transform 1 0 17952 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_876
timestamp 1581449086
transform 1 0 17748 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_877
timestamp 1581449086
transform 1 0 17544 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_878
timestamp 1581449086
transform 1 0 17340 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_879
timestamp 1581449086
transform 1 0 16932 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_880
timestamp 1581449086
transform 1 0 16524 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_881
timestamp 1581449086
transform 1 0 16320 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_882
timestamp 1581449086
transform 1 0 16116 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_883
timestamp 1581449086
transform 1 0 15504 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_884
timestamp 1581449086
transform 1 0 15300 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_885
timestamp 1581449086
transform 1 0 15096 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_886
timestamp 1581449086
transform 1 0 14892 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_887
timestamp 1581449086
transform 1 0 14688 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_888
timestamp 1581449086
transform 1 0 13668 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_889
timestamp 1581449086
transform 1 0 13464 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_890
timestamp 1581449086
transform 1 0 13056 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_891
timestamp 1581449086
transform 1 0 12444 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_892
timestamp 1581449086
transform 1 0 12240 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_893
timestamp 1581449086
transform 1 0 11832 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_894
timestamp 1581449086
transform 1 0 11628 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_895
timestamp 1581449086
transform 1 0 11424 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_896
timestamp 1581449086
transform 1 0 11220 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_897
timestamp 1581449086
transform 1 0 10812 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_898
timestamp 1581449086
transform 1 0 10404 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_899
timestamp 1581449086
transform 1 0 10200 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_900
timestamp 1581449086
transform 1 0 9792 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_901
timestamp 1581449086
transform 1 0 9588 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_902
timestamp 1581449086
transform 1 0 9384 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_903
timestamp 1581449086
transform 1 0 9180 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_904
timestamp 1581449086
transform 1 0 8976 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_905
timestamp 1581449086
transform 1 0 8364 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_906
timestamp 1581449086
transform 1 0 8160 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_907
timestamp 1581449086
transform 1 0 7956 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_908
timestamp 1581449086
transform 1 0 7548 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_909
timestamp 1581449086
transform 1 0 7344 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_910
timestamp 1581449086
transform 1 0 7140 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_911
timestamp 1581449086
transform 1 0 6936 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_912
timestamp 1581449086
transform 1 0 6732 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_913
timestamp 1581449086
transform 1 0 6324 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_914
timestamp 1581449086
transform 1 0 5916 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_915
timestamp 1581449086
transform 1 0 5304 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_916
timestamp 1581449086
transform 1 0 4692 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_917
timestamp 1581449086
transform 1 0 4488 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_918
timestamp 1581449086
transform 1 0 4284 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_919
timestamp 1581449086
transform 1 0 3876 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_920
timestamp 1581449086
transform 1 0 3468 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_921
timestamp 1581449086
transform 1 0 3264 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_922
timestamp 1581449086
transform 1 0 2856 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_923
timestamp 1581449086
transform 1 0 2652 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_924
timestamp 1581449086
transform 1 0 2040 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_925
timestamp 1581449086
transform 1 0 1836 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_926
timestamp 1581449086
transform 1 0 816 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_927
timestamp 1581449086
transform 1 0 612 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_928
timestamp 1581449086
transform 1 0 408 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_929
timestamp 1581449086
transform 1 0 204 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_930
timestamp 1581449086
transform 1 0 51816 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_931
timestamp 1581449086
transform 1 0 50592 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_932
timestamp 1581449086
transform 1 0 50388 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_933
timestamp 1581449086
transform 1 0 50184 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_934
timestamp 1581449086
transform 1 0 49980 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_935
timestamp 1581449086
transform 1 0 49572 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_936
timestamp 1581449086
transform 1 0 49164 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_937
timestamp 1581449086
transform 1 0 48960 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_938
timestamp 1581449086
transform 1 0 48348 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_939
timestamp 1581449086
transform 1 0 48144 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_940
timestamp 1581449086
transform 1 0 47532 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_941
timestamp 1581449086
transform 1 0 47328 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_942
timestamp 1581449086
transform 1 0 47124 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_943
timestamp 1581449086
transform 1 0 46920 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_944
timestamp 1581449086
transform 1 0 46716 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_945
timestamp 1581449086
transform 1 0 46308 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_946
timestamp 1581449086
transform 1 0 45900 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_947
timestamp 1581449086
transform 1 0 45288 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_948
timestamp 1581449086
transform 1 0 44676 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_949
timestamp 1581449086
transform 1 0 44472 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_950
timestamp 1581449086
transform 1 0 43860 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_951
timestamp 1581449086
transform 1 0 43248 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_952
timestamp 1581449086
transform 1 0 42840 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_953
timestamp 1581449086
transform 1 0 42636 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_954
timestamp 1581449086
transform 1 0 42432 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_955
timestamp 1581449086
transform 1 0 42024 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_956
timestamp 1581449086
transform 1 0 41412 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_957
timestamp 1581449086
transform 1 0 41004 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_958
timestamp 1581449086
transform 1 0 40800 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_959
timestamp 1581449086
transform 1 0 39984 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_960
timestamp 1581449086
transform 1 0 38964 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_961
timestamp 1581449086
transform 1 0 38760 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_962
timestamp 1581449086
transform 1 0 38352 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_963
timestamp 1581449086
transform 1 0 37740 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_964
timestamp 1581449086
transform 1 0 36924 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_965
timestamp 1581449086
transform 1 0 36108 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_966
timestamp 1581449086
transform 1 0 35496 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_967
timestamp 1581449086
transform 1 0 35292 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_968
timestamp 1581449086
transform 1 0 35088 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_969
timestamp 1581449086
transform 1 0 34884 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_970
timestamp 1581449086
transform 1 0 34680 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_971
timestamp 1581449086
transform 1 0 33864 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_972
timestamp 1581449086
transform 1 0 33660 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_973
timestamp 1581449086
transform 1 0 33456 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_974
timestamp 1581449086
transform 1 0 32844 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_975
timestamp 1581449086
transform 1 0 32232 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_976
timestamp 1581449086
transform 1 0 31824 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_977
timestamp 1581449086
transform 1 0 31212 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_978
timestamp 1581449086
transform 1 0 31008 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_979
timestamp 1581449086
transform 1 0 30804 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_980
timestamp 1581449086
transform 1 0 30600 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_981
timestamp 1581449086
transform 1 0 30396 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_982
timestamp 1581449086
transform 1 0 30192 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_983
timestamp 1581449086
transform 1 0 29988 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_984
timestamp 1581449086
transform 1 0 29580 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_985
timestamp 1581449086
transform 1 0 28968 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_986
timestamp 1581449086
transform 1 0 28764 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_987
timestamp 1581449086
transform 1 0 27744 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_988
timestamp 1581449086
transform 1 0 27540 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_989
timestamp 1581449086
transform 1 0 27132 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_990
timestamp 1581449086
transform 1 0 26316 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_991
timestamp 1581449086
transform 1 0 26112 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_992
timestamp 1581449086
transform 1 0 25908 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_993
timestamp 1581449086
transform 1 0 25296 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_994
timestamp 1581449086
transform 1 0 24888 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_995
timestamp 1581449086
transform 1 0 24480 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_996
timestamp 1581449086
transform 1 0 24276 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_997
timestamp 1581449086
transform 1 0 23868 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_998
timestamp 1581449086
transform 1 0 23460 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_999
timestamp 1581449086
transform 1 0 23256 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1000
timestamp 1581449086
transform 1 0 22236 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1001
timestamp 1581449086
transform 1 0 21624 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1002
timestamp 1581449086
transform 1 0 21216 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1003
timestamp 1581449086
transform 1 0 20604 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1004
timestamp 1581449086
transform 1 0 20400 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1005
timestamp 1581449086
transform 1 0 20196 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1006
timestamp 1581449086
transform 1 0 19992 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1007
timestamp 1581449086
transform 1 0 19788 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1008
timestamp 1581449086
transform 1 0 18360 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1009
timestamp 1581449086
transform 1 0 17952 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1010
timestamp 1581449086
transform 1 0 17748 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1011
timestamp 1581449086
transform 1 0 17136 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1012
timestamp 1581449086
transform 1 0 16728 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1013
timestamp 1581449086
transform 1 0 16320 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1014
timestamp 1581449086
transform 1 0 16116 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1015
timestamp 1581449086
transform 1 0 15912 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1016
timestamp 1581449086
transform 1 0 15300 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1017
timestamp 1581449086
transform 1 0 14892 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1018
timestamp 1581449086
transform 1 0 14688 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1019
timestamp 1581449086
transform 1 0 14484 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1020
timestamp 1581449086
transform 1 0 14280 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1021
timestamp 1581449086
transform 1 0 13872 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1022
timestamp 1581449086
transform 1 0 13260 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1023
timestamp 1581449086
transform 1 0 12648 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1024
timestamp 1581449086
transform 1 0 11424 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1025
timestamp 1581449086
transform 1 0 10812 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1026
timestamp 1581449086
transform 1 0 10608 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1027
timestamp 1581449086
transform 1 0 10404 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1028
timestamp 1581449086
transform 1 0 10200 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1029
timestamp 1581449086
transform 1 0 9996 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1030
timestamp 1581449086
transform 1 0 9588 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1031
timestamp 1581449086
transform 1 0 9384 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1032
timestamp 1581449086
transform 1 0 9180 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1033
timestamp 1581449086
transform 1 0 8976 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1034
timestamp 1581449086
transform 1 0 8772 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1035
timestamp 1581449086
transform 1 0 8364 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1036
timestamp 1581449086
transform 1 0 8160 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1037
timestamp 1581449086
transform 1 0 7752 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1038
timestamp 1581449086
transform 1 0 6936 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1039
timestamp 1581449086
transform 1 0 6732 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1040
timestamp 1581449086
transform 1 0 6528 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1041
timestamp 1581449086
transform 1 0 6324 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1042
timestamp 1581449086
transform 1 0 5508 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1043
timestamp 1581449086
transform 1 0 4896 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1044
timestamp 1581449086
transform 1 0 4488 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1045
timestamp 1581449086
transform 1 0 4284 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1046
timestamp 1581449086
transform 1 0 3264 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1047
timestamp 1581449086
transform 1 0 3060 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1048
timestamp 1581449086
transform 1 0 2856 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1049
timestamp 1581449086
transform 1 0 2448 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1050
timestamp 1581449086
transform 1 0 2040 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1051
timestamp 1581449086
transform 1 0 1020 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1052
timestamp 1581449086
transform 1 0 816 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1053
timestamp 1581449086
transform 1 0 204 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1054
timestamp 1581449086
transform 1 0 0 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_0
timestamp 1581449086
transform 1 0 52224 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_1
timestamp 1581449086
transform 1 0 50592 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_2
timestamp 1581449086
transform 1 0 48960 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_3
timestamp 1581449086
transform 1 0 47328 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_4
timestamp 1581449086
transform 1 0 45696 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_5
timestamp 1581449086
transform 1 0 44064 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_6
timestamp 1581449086
transform 1 0 42432 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_7
timestamp 1581449086
transform 1 0 40800 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_8
timestamp 1581449086
transform 1 0 39168 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_9
timestamp 1581449086
transform 1 0 37536 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_10
timestamp 1581449086
transform 1 0 35904 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_11
timestamp 1581449086
transform 1 0 34272 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_12
timestamp 1581449086
transform 1 0 32640 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_13
timestamp 1581449086
transform 1 0 31008 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_14
timestamp 1581449086
transform 1 0 29376 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_15
timestamp 1581449086
transform 1 0 27744 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_16
timestamp 1581449086
transform 1 0 26112 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_17
timestamp 1581449086
transform 1 0 24480 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_18
timestamp 1581449086
transform 1 0 22848 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_19
timestamp 1581449086
transform 1 0 21216 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_20
timestamp 1581449086
transform 1 0 19584 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_21
timestamp 1581449086
transform 1 0 17952 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_22
timestamp 1581449086
transform 1 0 16320 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_23
timestamp 1581449086
transform 1 0 14688 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_24
timestamp 1581449086
transform 1 0 13056 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_25
timestamp 1581449086
transform 1 0 11424 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_26
timestamp 1581449086
transform 1 0 9792 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_27
timestamp 1581449086
transform 1 0 8160 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_28
timestamp 1581449086
transform 1 0 6528 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_29
timestamp 1581449086
transform 1 0 4896 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_30
timestamp 1581449086
transform 1 0 3264 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_31
timestamp 1581449086
transform 1 0 1632 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_32
timestamp 1581449086
transform 1 0 0 0 1 2609
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_33
timestamp 1581449086
transform 1 0 52224 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_34
timestamp 1581449086
transform 1 0 50592 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_35
timestamp 1581449086
transform 1 0 48960 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_36
timestamp 1581449086
transform 1 0 47328 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_37
timestamp 1581449086
transform 1 0 45696 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_38
timestamp 1581449086
transform 1 0 44064 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_39
timestamp 1581449086
transform 1 0 42432 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_40
timestamp 1581449086
transform 1 0 40800 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_41
timestamp 1581449086
transform 1 0 39168 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_42
timestamp 1581449086
transform 1 0 37536 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_43
timestamp 1581449086
transform 1 0 35904 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_44
timestamp 1581449086
transform 1 0 34272 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_45
timestamp 1581449086
transform 1 0 32640 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_46
timestamp 1581449086
transform 1 0 31008 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_47
timestamp 1581449086
transform 1 0 29376 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_48
timestamp 1581449086
transform 1 0 27744 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_49
timestamp 1581449086
transform 1 0 26112 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_50
timestamp 1581449086
transform 1 0 24480 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_51
timestamp 1581449086
transform 1 0 22848 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_52
timestamp 1581449086
transform 1 0 21216 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_53
timestamp 1581449086
transform 1 0 19584 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_54
timestamp 1581449086
transform 1 0 17952 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_55
timestamp 1581449086
transform 1 0 16320 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_56
timestamp 1581449086
transform 1 0 14688 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_57
timestamp 1581449086
transform 1 0 13056 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_58
timestamp 1581449086
transform 1 0 11424 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_59
timestamp 1581449086
transform 1 0 9792 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_60
timestamp 1581449086
transform 1 0 8160 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_61
timestamp 1581449086
transform 1 0 6528 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_62
timestamp 1581449086
transform 1 0 4896 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_63
timestamp 1581449086
transform 1 0 3264 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_64
timestamp 1581449086
transform 1 0 1632 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_65
timestamp 1581449086
transform 1 0 0 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_66
timestamp 1581449086
transform 1 0 52224 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_67
timestamp 1581449086
transform 1 0 50592 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_68
timestamp 1581449086
transform 1 0 48960 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_69
timestamp 1581449086
transform 1 0 47328 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_70
timestamp 1581449086
transform 1 0 45696 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_71
timestamp 1581449086
transform 1 0 44064 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_72
timestamp 1581449086
transform 1 0 42432 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_73
timestamp 1581449086
transform 1 0 40800 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_74
timestamp 1581449086
transform 1 0 39168 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_75
timestamp 1581449086
transform 1 0 37536 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_76
timestamp 1581449086
transform 1 0 35904 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_77
timestamp 1581449086
transform 1 0 34272 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_78
timestamp 1581449086
transform 1 0 32640 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_79
timestamp 1581449086
transform 1 0 31008 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_80
timestamp 1581449086
transform 1 0 29376 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_81
timestamp 1581449086
transform 1 0 27744 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_82
timestamp 1581449086
transform 1 0 26112 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_83
timestamp 1581449086
transform 1 0 24480 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_84
timestamp 1581449086
transform 1 0 22848 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_85
timestamp 1581449086
transform 1 0 21216 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_86
timestamp 1581449086
transform 1 0 19584 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_87
timestamp 1581449086
transform 1 0 17952 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_88
timestamp 1581449086
transform 1 0 16320 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_89
timestamp 1581449086
transform 1 0 14688 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_90
timestamp 1581449086
transform 1 0 13056 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_91
timestamp 1581449086
transform 1 0 11424 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_92
timestamp 1581449086
transform 1 0 9792 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_93
timestamp 1581449086
transform 1 0 8160 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_94
timestamp 1581449086
transform 1 0 6528 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_95
timestamp 1581449086
transform 1 0 4896 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_96
timestamp 1581449086
transform 1 0 3264 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_97
timestamp 1581449086
transform 1 0 1632 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_98
timestamp 1581449086
transform 1 0 0 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_99
timestamp 1581449086
transform 1 0 52224 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_100
timestamp 1581449086
transform 1 0 50592 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_101
timestamp 1581449086
transform 1 0 48960 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_102
timestamp 1581449086
transform 1 0 47328 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_103
timestamp 1581449086
transform 1 0 45696 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_104
timestamp 1581449086
transform 1 0 44064 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_105
timestamp 1581449086
transform 1 0 42432 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_106
timestamp 1581449086
transform 1 0 40800 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_107
timestamp 1581449086
transform 1 0 39168 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_108
timestamp 1581449086
transform 1 0 37536 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_109
timestamp 1581449086
transform 1 0 35904 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_110
timestamp 1581449086
transform 1 0 34272 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_111
timestamp 1581449086
transform 1 0 32640 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_112
timestamp 1581449086
transform 1 0 31008 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_113
timestamp 1581449086
transform 1 0 29376 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_114
timestamp 1581449086
transform 1 0 27744 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_115
timestamp 1581449086
transform 1 0 26112 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_116
timestamp 1581449086
transform 1 0 24480 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_117
timestamp 1581449086
transform 1 0 22848 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_118
timestamp 1581449086
transform 1 0 21216 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_119
timestamp 1581449086
transform 1 0 19584 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_120
timestamp 1581449086
transform 1 0 17952 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_121
timestamp 1581449086
transform 1 0 16320 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_122
timestamp 1581449086
transform 1 0 14688 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_123
timestamp 1581449086
transform 1 0 13056 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_124
timestamp 1581449086
transform 1 0 11424 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_125
timestamp 1581449086
transform 1 0 9792 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_126
timestamp 1581449086
transform 1 0 8160 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_127
timestamp 1581449086
transform 1 0 6528 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_128
timestamp 1581449086
transform 1 0 4896 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_129
timestamp 1581449086
transform 1 0 3264 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_130
timestamp 1581449086
transform 1 0 1632 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_131
timestamp 1581449086
transform 1 0 0 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_132
timestamp 1581449086
transform 1 0 52224 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_133
timestamp 1581449086
transform 1 0 50592 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_134
timestamp 1581449086
transform 1 0 48960 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_135
timestamp 1581449086
transform 1 0 47328 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_136
timestamp 1581449086
transform 1 0 45696 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_137
timestamp 1581449086
transform 1 0 44064 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_138
timestamp 1581449086
transform 1 0 42432 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_139
timestamp 1581449086
transform 1 0 40800 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_140
timestamp 1581449086
transform 1 0 39168 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_141
timestamp 1581449086
transform 1 0 37536 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_142
timestamp 1581449086
transform 1 0 35904 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_143
timestamp 1581449086
transform 1 0 34272 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_144
timestamp 1581449086
transform 1 0 32640 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_145
timestamp 1581449086
transform 1 0 31008 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_146
timestamp 1581449086
transform 1 0 29376 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_147
timestamp 1581449086
transform 1 0 27744 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_148
timestamp 1581449086
transform 1 0 26112 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_149
timestamp 1581449086
transform 1 0 24480 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_150
timestamp 1581449086
transform 1 0 22848 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_151
timestamp 1581449086
transform 1 0 21216 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_152
timestamp 1581449086
transform 1 0 19584 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_153
timestamp 1581449086
transform 1 0 17952 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_154
timestamp 1581449086
transform 1 0 16320 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_155
timestamp 1581449086
transform 1 0 14688 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_156
timestamp 1581449086
transform 1 0 13056 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_157
timestamp 1581449086
transform 1 0 11424 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_158
timestamp 1581449086
transform 1 0 9792 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_159
timestamp 1581449086
transform 1 0 8160 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_160
timestamp 1581449086
transform 1 0 6528 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_161
timestamp 1581449086
transform 1 0 4896 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_162
timestamp 1581449086
transform 1 0 3264 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_163
timestamp 1581449086
transform 1 0 1632 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_164
timestamp 1581449086
transform 1 0 0 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_165
timestamp 1581449086
transform 1 0 52224 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_166
timestamp 1581449086
transform 1 0 50592 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_167
timestamp 1581449086
transform 1 0 48960 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_168
timestamp 1581449086
transform 1 0 47328 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_169
timestamp 1581449086
transform 1 0 45696 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_170
timestamp 1581449086
transform 1 0 44064 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_171
timestamp 1581449086
transform 1 0 42432 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_172
timestamp 1581449086
transform 1 0 40800 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_173
timestamp 1581449086
transform 1 0 39168 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_174
timestamp 1581449086
transform 1 0 37536 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_175
timestamp 1581449086
transform 1 0 35904 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_176
timestamp 1581449086
transform 1 0 34272 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_177
timestamp 1581449086
transform 1 0 32640 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_178
timestamp 1581449086
transform 1 0 31008 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_179
timestamp 1581449086
transform 1 0 29376 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_180
timestamp 1581449086
transform 1 0 27744 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_181
timestamp 1581449086
transform 1 0 26112 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_182
timestamp 1581449086
transform 1 0 24480 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_183
timestamp 1581449086
transform 1 0 22848 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_184
timestamp 1581449086
transform 1 0 21216 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_185
timestamp 1581449086
transform 1 0 19584 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_186
timestamp 1581449086
transform 1 0 17952 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_187
timestamp 1581449086
transform 1 0 16320 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_188
timestamp 1581449086
transform 1 0 14688 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_189
timestamp 1581449086
transform 1 0 13056 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_190
timestamp 1581449086
transform 1 0 11424 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_191
timestamp 1581449086
transform 1 0 9792 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_192
timestamp 1581449086
transform 1 0 8160 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_193
timestamp 1581449086
transform 1 0 6528 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_194
timestamp 1581449086
transform 1 0 4896 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_195
timestamp 1581449086
transform 1 0 3264 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_196
timestamp 1581449086
transform 1 0 1632 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_197
timestamp 1581449086
transform 1 0 0 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_198
timestamp 1581449086
transform 1 0 52224 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_199
timestamp 1581449086
transform 1 0 50592 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_200
timestamp 1581449086
transform 1 0 48960 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_201
timestamp 1581449086
transform 1 0 47328 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_202
timestamp 1581449086
transform 1 0 45696 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_203
timestamp 1581449086
transform 1 0 44064 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_204
timestamp 1581449086
transform 1 0 42432 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_205
timestamp 1581449086
transform 1 0 40800 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_206
timestamp 1581449086
transform 1 0 39168 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_207
timestamp 1581449086
transform 1 0 37536 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_208
timestamp 1581449086
transform 1 0 35904 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_209
timestamp 1581449086
transform 1 0 34272 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_210
timestamp 1581449086
transform 1 0 32640 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_211
timestamp 1581449086
transform 1 0 31008 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_212
timestamp 1581449086
transform 1 0 29376 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_213
timestamp 1581449086
transform 1 0 27744 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_214
timestamp 1581449086
transform 1 0 26112 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_215
timestamp 1581449086
transform 1 0 24480 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_216
timestamp 1581449086
transform 1 0 22848 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_217
timestamp 1581449086
transform 1 0 21216 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_218
timestamp 1581449086
transform 1 0 19584 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_219
timestamp 1581449086
transform 1 0 17952 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_220
timestamp 1581449086
transform 1 0 16320 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_221
timestamp 1581449086
transform 1 0 14688 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_222
timestamp 1581449086
transform 1 0 13056 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_223
timestamp 1581449086
transform 1 0 11424 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_224
timestamp 1581449086
transform 1 0 9792 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_225
timestamp 1581449086
transform 1 0 8160 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_226
timestamp 1581449086
transform 1 0 6528 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_227
timestamp 1581449086
transform 1 0 4896 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_228
timestamp 1581449086
transform 1 0 3264 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_229
timestamp 1581449086
transform 1 0 1632 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_230
timestamp 1581449086
transform 1 0 0 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_231
timestamp 1581449086
transform 1 0 52224 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_232
timestamp 1581449086
transform 1 0 50592 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_233
timestamp 1581449086
transform 1 0 48960 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_234
timestamp 1581449086
transform 1 0 47328 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_235
timestamp 1581449086
transform 1 0 45696 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_236
timestamp 1581449086
transform 1 0 44064 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_237
timestamp 1581449086
transform 1 0 42432 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_238
timestamp 1581449086
transform 1 0 40800 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_239
timestamp 1581449086
transform 1 0 39168 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_240
timestamp 1581449086
transform 1 0 37536 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_241
timestamp 1581449086
transform 1 0 35904 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_242
timestamp 1581449086
transform 1 0 34272 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_243
timestamp 1581449086
transform 1 0 32640 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_244
timestamp 1581449086
transform 1 0 31008 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_245
timestamp 1581449086
transform 1 0 29376 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_246
timestamp 1581449086
transform 1 0 27744 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_247
timestamp 1581449086
transform 1 0 26112 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_248
timestamp 1581449086
transform 1 0 24480 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_249
timestamp 1581449086
transform 1 0 22848 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_250
timestamp 1581449086
transform 1 0 21216 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_251
timestamp 1581449086
transform 1 0 19584 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_252
timestamp 1581449086
transform 1 0 17952 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_253
timestamp 1581449086
transform 1 0 16320 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_254
timestamp 1581449086
transform 1 0 14688 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_255
timestamp 1581449086
transform 1 0 13056 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_256
timestamp 1581449086
transform 1 0 11424 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_257
timestamp 1581449086
transform 1 0 9792 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_258
timestamp 1581449086
transform 1 0 8160 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_259
timestamp 1581449086
transform 1 0 6528 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_260
timestamp 1581449086
transform 1 0 4896 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_261
timestamp 1581449086
transform 1 0 3264 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_262
timestamp 1581449086
transform 1 0 1632 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_263
timestamp 1581449086
transform 1 0 0 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_264
timestamp 1581449086
transform 1 0 52224 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_265
timestamp 1581449086
transform 1 0 50592 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_266
timestamp 1581449086
transform 1 0 48960 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_267
timestamp 1581449086
transform 1 0 47328 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_268
timestamp 1581449086
transform 1 0 45696 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_269
timestamp 1581449086
transform 1 0 44064 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_270
timestamp 1581449086
transform 1 0 42432 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_271
timestamp 1581449086
transform 1 0 40800 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_272
timestamp 1581449086
transform 1 0 39168 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_273
timestamp 1581449086
transform 1 0 37536 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_274
timestamp 1581449086
transform 1 0 35904 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_275
timestamp 1581449086
transform 1 0 34272 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_276
timestamp 1581449086
transform 1 0 32640 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_277
timestamp 1581449086
transform 1 0 31008 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_278
timestamp 1581449086
transform 1 0 29376 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_279
timestamp 1581449086
transform 1 0 27744 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_280
timestamp 1581449086
transform 1 0 26112 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_281
timestamp 1581449086
transform 1 0 24480 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_282
timestamp 1581449086
transform 1 0 22848 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_283
timestamp 1581449086
transform 1 0 21216 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_284
timestamp 1581449086
transform 1 0 19584 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_285
timestamp 1581449086
transform 1 0 17952 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_286
timestamp 1581449086
transform 1 0 16320 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_287
timestamp 1581449086
transform 1 0 14688 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_288
timestamp 1581449086
transform 1 0 13056 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_289
timestamp 1581449086
transform 1 0 11424 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_290
timestamp 1581449086
transform 1 0 9792 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_291
timestamp 1581449086
transform 1 0 8160 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_292
timestamp 1581449086
transform 1 0 6528 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_293
timestamp 1581449086
transform 1 0 4896 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_294
timestamp 1581449086
transform 1 0 3264 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_295
timestamp 1581449086
transform 1 0 1632 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_296
timestamp 1581449086
transform 1 0 0 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_precharge_array  sky130_rom_krom_rom_precharge_array_0
timestamp 1581449086
transform 1 0 0 0 1 128
box 0 -212 52332 408
<< labels >>
rlabel metal2 s 61 368 89 396 4 precharge
port 3 nsew
rlabel metal2 s 19 1013 47 1041 4 wl_0_0
port 5 nsew
rlabel metal2 s 19 1217 47 1245 4 wl_0_1
port 7 nsew
rlabel metal2 s 19 1421 47 1449 4 wl_0_2
port 9 nsew
rlabel metal2 s 19 1625 47 1653 4 wl_0_3
port 11 nsew
rlabel metal2 s 19 1829 47 1857 4 wl_0_4
port 13 nsew
rlabel metal2 s 19 2033 47 2061 4 wl_0_5
port 15 nsew
rlabel metal2 s 19 2237 47 2265 4 wl_0_6
port 17 nsew
rlabel metal2 s 19 2441 47 2469 4 wl_0_7
port 19 nsew
rlabel metal1 s 128 -14 156 14 4 bl_0_0
port 21 nsew
rlabel metal1 s 332 -14 360 14 4 bl_0_1
port 23 nsew
rlabel metal1 s 536 -14 564 14 4 bl_0_2
port 25 nsew
rlabel metal1 s 740 -14 768 14 4 bl_0_3
port 27 nsew
rlabel metal1 s 944 -14 972 14 4 bl_0_4
port 29 nsew
rlabel metal1 s 1148 -14 1176 14 4 bl_0_5
port 31 nsew
rlabel metal1 s 1352 -14 1380 14 4 bl_0_6
port 33 nsew
rlabel metal1 s 1556 -14 1584 14 4 bl_0_7
port 35 nsew
rlabel metal1 s 1760 -14 1788 14 4 bl_0_8
port 37 nsew
rlabel metal1 s 1964 -14 1992 14 4 bl_0_9
port 39 nsew
rlabel metal1 s 2168 -14 2196 14 4 bl_0_10
port 41 nsew
rlabel metal1 s 2372 -14 2400 14 4 bl_0_11
port 43 nsew
rlabel metal1 s 2576 -14 2604 14 4 bl_0_12
port 45 nsew
rlabel metal1 s 2780 -14 2808 14 4 bl_0_13
port 47 nsew
rlabel metal1 s 2984 -14 3012 14 4 bl_0_14
port 49 nsew
rlabel metal1 s 3188 -14 3216 14 4 bl_0_15
port 51 nsew
rlabel metal1 s 3392 -14 3420 14 4 bl_0_16
port 53 nsew
rlabel metal1 s 3596 -14 3624 14 4 bl_0_17
port 55 nsew
rlabel metal1 s 3800 -14 3828 14 4 bl_0_18
port 57 nsew
rlabel metal1 s 4004 -14 4032 14 4 bl_0_19
port 59 nsew
rlabel metal1 s 4208 -14 4236 14 4 bl_0_20
port 61 nsew
rlabel metal1 s 4412 -14 4440 14 4 bl_0_21
port 63 nsew
rlabel metal1 s 4616 -14 4644 14 4 bl_0_22
port 65 nsew
rlabel metal1 s 4820 -14 4848 14 4 bl_0_23
port 67 nsew
rlabel metal1 s 5024 -14 5052 14 4 bl_0_24
port 69 nsew
rlabel metal1 s 5228 -14 5256 14 4 bl_0_25
port 71 nsew
rlabel metal1 s 5432 -14 5460 14 4 bl_0_26
port 73 nsew
rlabel metal1 s 5636 -14 5664 14 4 bl_0_27
port 75 nsew
rlabel metal1 s 5840 -14 5868 14 4 bl_0_28
port 77 nsew
rlabel metal1 s 6044 -14 6072 14 4 bl_0_29
port 79 nsew
rlabel metal1 s 6248 -14 6276 14 4 bl_0_30
port 81 nsew
rlabel metal1 s 6452 -14 6480 14 4 bl_0_31
port 83 nsew
rlabel metal1 s 6656 -14 6684 14 4 bl_0_32
port 85 nsew
rlabel metal1 s 6860 -14 6888 14 4 bl_0_33
port 87 nsew
rlabel metal1 s 7064 -14 7092 14 4 bl_0_34
port 89 nsew
rlabel metal1 s 7268 -14 7296 14 4 bl_0_35
port 91 nsew
rlabel metal1 s 7472 -14 7500 14 4 bl_0_36
port 93 nsew
rlabel metal1 s 7676 -14 7704 14 4 bl_0_37
port 95 nsew
rlabel metal1 s 7880 -14 7908 14 4 bl_0_38
port 97 nsew
rlabel metal1 s 8084 -14 8112 14 4 bl_0_39
port 99 nsew
rlabel metal1 s 8288 -14 8316 14 4 bl_0_40
port 101 nsew
rlabel metal1 s 8492 -14 8520 14 4 bl_0_41
port 103 nsew
rlabel metal1 s 8696 -14 8724 14 4 bl_0_42
port 105 nsew
rlabel metal1 s 8900 -14 8928 14 4 bl_0_43
port 107 nsew
rlabel metal1 s 9104 -14 9132 14 4 bl_0_44
port 109 nsew
rlabel metal1 s 9308 -14 9336 14 4 bl_0_45
port 111 nsew
rlabel metal1 s 9512 -14 9540 14 4 bl_0_46
port 113 nsew
rlabel metal1 s 9716 -14 9744 14 4 bl_0_47
port 115 nsew
rlabel metal1 s 9920 -14 9948 14 4 bl_0_48
port 117 nsew
rlabel metal1 s 10124 -14 10152 14 4 bl_0_49
port 119 nsew
rlabel metal1 s 10328 -14 10356 14 4 bl_0_50
port 121 nsew
rlabel metal1 s 10532 -14 10560 14 4 bl_0_51
port 123 nsew
rlabel metal1 s 10736 -14 10764 14 4 bl_0_52
port 125 nsew
rlabel metal1 s 10940 -14 10968 14 4 bl_0_53
port 127 nsew
rlabel metal1 s 11144 -14 11172 14 4 bl_0_54
port 129 nsew
rlabel metal1 s 11348 -14 11376 14 4 bl_0_55
port 131 nsew
rlabel metal1 s 11552 -14 11580 14 4 bl_0_56
port 133 nsew
rlabel metal1 s 11756 -14 11784 14 4 bl_0_57
port 135 nsew
rlabel metal1 s 11960 -14 11988 14 4 bl_0_58
port 137 nsew
rlabel metal1 s 12164 -14 12192 14 4 bl_0_59
port 139 nsew
rlabel metal1 s 12368 -14 12396 14 4 bl_0_60
port 141 nsew
rlabel metal1 s 12572 -14 12600 14 4 bl_0_61
port 143 nsew
rlabel metal1 s 12776 -14 12804 14 4 bl_0_62
port 145 nsew
rlabel metal1 s 12980 -14 13008 14 4 bl_0_63
port 147 nsew
rlabel metal1 s 13184 -14 13212 14 4 bl_0_64
port 149 nsew
rlabel metal1 s 13388 -14 13416 14 4 bl_0_65
port 151 nsew
rlabel metal1 s 13592 -14 13620 14 4 bl_0_66
port 153 nsew
rlabel metal1 s 13796 -14 13824 14 4 bl_0_67
port 155 nsew
rlabel metal1 s 14000 -14 14028 14 4 bl_0_68
port 157 nsew
rlabel metal1 s 14204 -14 14232 14 4 bl_0_69
port 159 nsew
rlabel metal1 s 14408 -14 14436 14 4 bl_0_70
port 161 nsew
rlabel metal1 s 14612 -14 14640 14 4 bl_0_71
port 163 nsew
rlabel metal1 s 14816 -14 14844 14 4 bl_0_72
port 165 nsew
rlabel metal1 s 15020 -14 15048 14 4 bl_0_73
port 167 nsew
rlabel metal1 s 15224 -14 15252 14 4 bl_0_74
port 169 nsew
rlabel metal1 s 15428 -14 15456 14 4 bl_0_75
port 171 nsew
rlabel metal1 s 15632 -14 15660 14 4 bl_0_76
port 173 nsew
rlabel metal1 s 15836 -14 15864 14 4 bl_0_77
port 175 nsew
rlabel metal1 s 16040 -14 16068 14 4 bl_0_78
port 177 nsew
rlabel metal1 s 16244 -14 16272 14 4 bl_0_79
port 179 nsew
rlabel metal1 s 16448 -14 16476 14 4 bl_0_80
port 181 nsew
rlabel metal1 s 16652 -14 16680 14 4 bl_0_81
port 183 nsew
rlabel metal1 s 16856 -14 16884 14 4 bl_0_82
port 185 nsew
rlabel metal1 s 17060 -14 17088 14 4 bl_0_83
port 187 nsew
rlabel metal1 s 17264 -14 17292 14 4 bl_0_84
port 189 nsew
rlabel metal1 s 17468 -14 17496 14 4 bl_0_85
port 191 nsew
rlabel metal1 s 17672 -14 17700 14 4 bl_0_86
port 193 nsew
rlabel metal1 s 17876 -14 17904 14 4 bl_0_87
port 195 nsew
rlabel metal1 s 18080 -14 18108 14 4 bl_0_88
port 197 nsew
rlabel metal1 s 18284 -14 18312 14 4 bl_0_89
port 199 nsew
rlabel metal1 s 18488 -14 18516 14 4 bl_0_90
port 201 nsew
rlabel metal1 s 18692 -14 18720 14 4 bl_0_91
port 203 nsew
rlabel metal1 s 18896 -14 18924 14 4 bl_0_92
port 205 nsew
rlabel metal1 s 19100 -14 19128 14 4 bl_0_93
port 207 nsew
rlabel metal1 s 19304 -14 19332 14 4 bl_0_94
port 209 nsew
rlabel metal1 s 19508 -14 19536 14 4 bl_0_95
port 211 nsew
rlabel metal1 s 19712 -14 19740 14 4 bl_0_96
port 213 nsew
rlabel metal1 s 19916 -14 19944 14 4 bl_0_97
port 215 nsew
rlabel metal1 s 20120 -14 20148 14 4 bl_0_98
port 217 nsew
rlabel metal1 s 20324 -14 20352 14 4 bl_0_99
port 219 nsew
rlabel metal1 s 20528 -14 20556 14 4 bl_0_100
port 221 nsew
rlabel metal1 s 20732 -14 20760 14 4 bl_0_101
port 223 nsew
rlabel metal1 s 20936 -14 20964 14 4 bl_0_102
port 225 nsew
rlabel metal1 s 21140 -14 21168 14 4 bl_0_103
port 227 nsew
rlabel metal1 s 21344 -14 21372 14 4 bl_0_104
port 229 nsew
rlabel metal1 s 21548 -14 21576 14 4 bl_0_105
port 231 nsew
rlabel metal1 s 21752 -14 21780 14 4 bl_0_106
port 233 nsew
rlabel metal1 s 21956 -14 21984 14 4 bl_0_107
port 235 nsew
rlabel metal1 s 22160 -14 22188 14 4 bl_0_108
port 237 nsew
rlabel metal1 s 22364 -14 22392 14 4 bl_0_109
port 239 nsew
rlabel metal1 s 22568 -14 22596 14 4 bl_0_110
port 241 nsew
rlabel metal1 s 22772 -14 22800 14 4 bl_0_111
port 243 nsew
rlabel metal1 s 22976 -14 23004 14 4 bl_0_112
port 245 nsew
rlabel metal1 s 23180 -14 23208 14 4 bl_0_113
port 247 nsew
rlabel metal1 s 23384 -14 23412 14 4 bl_0_114
port 249 nsew
rlabel metal1 s 23588 -14 23616 14 4 bl_0_115
port 251 nsew
rlabel metal1 s 23792 -14 23820 14 4 bl_0_116
port 253 nsew
rlabel metal1 s 23996 -14 24024 14 4 bl_0_117
port 255 nsew
rlabel metal1 s 24200 -14 24228 14 4 bl_0_118
port 257 nsew
rlabel metal1 s 24404 -14 24432 14 4 bl_0_119
port 259 nsew
rlabel metal1 s 24608 -14 24636 14 4 bl_0_120
port 261 nsew
rlabel metal1 s 24812 -14 24840 14 4 bl_0_121
port 263 nsew
rlabel metal1 s 25016 -14 25044 14 4 bl_0_122
port 265 nsew
rlabel metal1 s 25220 -14 25248 14 4 bl_0_123
port 267 nsew
rlabel metal1 s 25424 -14 25452 14 4 bl_0_124
port 269 nsew
rlabel metal1 s 25628 -14 25656 14 4 bl_0_125
port 271 nsew
rlabel metal1 s 25832 -14 25860 14 4 bl_0_126
port 273 nsew
rlabel metal1 s 26036 -14 26064 14 4 bl_0_127
port 275 nsew
rlabel metal1 s 26240 -14 26268 14 4 bl_0_128
port 277 nsew
rlabel metal1 s 26444 -14 26472 14 4 bl_0_129
port 279 nsew
rlabel metal1 s 26648 -14 26676 14 4 bl_0_130
port 281 nsew
rlabel metal1 s 26852 -14 26880 14 4 bl_0_131
port 283 nsew
rlabel metal1 s 27056 -14 27084 14 4 bl_0_132
port 285 nsew
rlabel metal1 s 27260 -14 27288 14 4 bl_0_133
port 287 nsew
rlabel metal1 s 27464 -14 27492 14 4 bl_0_134
port 289 nsew
rlabel metal1 s 27668 -14 27696 14 4 bl_0_135
port 291 nsew
rlabel metal1 s 27872 -14 27900 14 4 bl_0_136
port 293 nsew
rlabel metal1 s 28076 -14 28104 14 4 bl_0_137
port 295 nsew
rlabel metal1 s 28280 -14 28308 14 4 bl_0_138
port 297 nsew
rlabel metal1 s 28484 -14 28512 14 4 bl_0_139
port 299 nsew
rlabel metal1 s 28688 -14 28716 14 4 bl_0_140
port 301 nsew
rlabel metal1 s 28892 -14 28920 14 4 bl_0_141
port 303 nsew
rlabel metal1 s 29096 -14 29124 14 4 bl_0_142
port 305 nsew
rlabel metal1 s 29300 -14 29328 14 4 bl_0_143
port 307 nsew
rlabel metal1 s 29504 -14 29532 14 4 bl_0_144
port 309 nsew
rlabel metal1 s 29708 -14 29736 14 4 bl_0_145
port 311 nsew
rlabel metal1 s 29912 -14 29940 14 4 bl_0_146
port 313 nsew
rlabel metal1 s 30116 -14 30144 14 4 bl_0_147
port 315 nsew
rlabel metal1 s 30320 -14 30348 14 4 bl_0_148
port 317 nsew
rlabel metal1 s 30524 -14 30552 14 4 bl_0_149
port 319 nsew
rlabel metal1 s 30728 -14 30756 14 4 bl_0_150
port 321 nsew
rlabel metal1 s 30932 -14 30960 14 4 bl_0_151
port 323 nsew
rlabel metal1 s 31136 -14 31164 14 4 bl_0_152
port 325 nsew
rlabel metal1 s 31340 -14 31368 14 4 bl_0_153
port 327 nsew
rlabel metal1 s 31544 -14 31572 14 4 bl_0_154
port 329 nsew
rlabel metal1 s 31748 -14 31776 14 4 bl_0_155
port 331 nsew
rlabel metal1 s 31952 -14 31980 14 4 bl_0_156
port 333 nsew
rlabel metal1 s 32156 -14 32184 14 4 bl_0_157
port 335 nsew
rlabel metal1 s 32360 -14 32388 14 4 bl_0_158
port 337 nsew
rlabel metal1 s 32564 -14 32592 14 4 bl_0_159
port 339 nsew
rlabel metal1 s 32768 -14 32796 14 4 bl_0_160
port 341 nsew
rlabel metal1 s 32972 -14 33000 14 4 bl_0_161
port 343 nsew
rlabel metal1 s 33176 -14 33204 14 4 bl_0_162
port 345 nsew
rlabel metal1 s 33380 -14 33408 14 4 bl_0_163
port 347 nsew
rlabel metal1 s 33584 -14 33612 14 4 bl_0_164
port 349 nsew
rlabel metal1 s 33788 -14 33816 14 4 bl_0_165
port 351 nsew
rlabel metal1 s 33992 -14 34020 14 4 bl_0_166
port 353 nsew
rlabel metal1 s 34196 -14 34224 14 4 bl_0_167
port 355 nsew
rlabel metal1 s 34400 -14 34428 14 4 bl_0_168
port 357 nsew
rlabel metal1 s 34604 -14 34632 14 4 bl_0_169
port 359 nsew
rlabel metal1 s 34808 -14 34836 14 4 bl_0_170
port 361 nsew
rlabel metal1 s 35012 -14 35040 14 4 bl_0_171
port 363 nsew
rlabel metal1 s 35216 -14 35244 14 4 bl_0_172
port 365 nsew
rlabel metal1 s 35420 -14 35448 14 4 bl_0_173
port 367 nsew
rlabel metal1 s 35624 -14 35652 14 4 bl_0_174
port 369 nsew
rlabel metal1 s 35828 -14 35856 14 4 bl_0_175
port 371 nsew
rlabel metal1 s 36032 -14 36060 14 4 bl_0_176
port 373 nsew
rlabel metal1 s 36236 -14 36264 14 4 bl_0_177
port 375 nsew
rlabel metal1 s 36440 -14 36468 14 4 bl_0_178
port 377 nsew
rlabel metal1 s 36644 -14 36672 14 4 bl_0_179
port 379 nsew
rlabel metal1 s 36848 -14 36876 14 4 bl_0_180
port 381 nsew
rlabel metal1 s 37052 -14 37080 14 4 bl_0_181
port 383 nsew
rlabel metal1 s 37256 -14 37284 14 4 bl_0_182
port 385 nsew
rlabel metal1 s 37460 -14 37488 14 4 bl_0_183
port 387 nsew
rlabel metal1 s 37664 -14 37692 14 4 bl_0_184
port 389 nsew
rlabel metal1 s 37868 -14 37896 14 4 bl_0_185
port 391 nsew
rlabel metal1 s 38072 -14 38100 14 4 bl_0_186
port 393 nsew
rlabel metal1 s 38276 -14 38304 14 4 bl_0_187
port 395 nsew
rlabel metal1 s 38480 -14 38508 14 4 bl_0_188
port 397 nsew
rlabel metal1 s 38684 -14 38712 14 4 bl_0_189
port 399 nsew
rlabel metal1 s 38888 -14 38916 14 4 bl_0_190
port 401 nsew
rlabel metal1 s 39092 -14 39120 14 4 bl_0_191
port 403 nsew
rlabel metal1 s 39296 -14 39324 14 4 bl_0_192
port 405 nsew
rlabel metal1 s 39500 -14 39528 14 4 bl_0_193
port 407 nsew
rlabel metal1 s 39704 -14 39732 14 4 bl_0_194
port 409 nsew
rlabel metal1 s 39908 -14 39936 14 4 bl_0_195
port 411 nsew
rlabel metal1 s 40112 -14 40140 14 4 bl_0_196
port 413 nsew
rlabel metal1 s 40316 -14 40344 14 4 bl_0_197
port 415 nsew
rlabel metal1 s 40520 -14 40548 14 4 bl_0_198
port 417 nsew
rlabel metal1 s 40724 -14 40752 14 4 bl_0_199
port 419 nsew
rlabel metal1 s 40928 -14 40956 14 4 bl_0_200
port 421 nsew
rlabel metal1 s 41132 -14 41160 14 4 bl_0_201
port 423 nsew
rlabel metal1 s 41336 -14 41364 14 4 bl_0_202
port 425 nsew
rlabel metal1 s 41540 -14 41568 14 4 bl_0_203
port 427 nsew
rlabel metal1 s 41744 -14 41772 14 4 bl_0_204
port 429 nsew
rlabel metal1 s 41948 -14 41976 14 4 bl_0_205
port 431 nsew
rlabel metal1 s 42152 -14 42180 14 4 bl_0_206
port 433 nsew
rlabel metal1 s 42356 -14 42384 14 4 bl_0_207
port 435 nsew
rlabel metal1 s 42560 -14 42588 14 4 bl_0_208
port 437 nsew
rlabel metal1 s 42764 -14 42792 14 4 bl_0_209
port 439 nsew
rlabel metal1 s 42968 -14 42996 14 4 bl_0_210
port 441 nsew
rlabel metal1 s 43172 -14 43200 14 4 bl_0_211
port 443 nsew
rlabel metal1 s 43376 -14 43404 14 4 bl_0_212
port 445 nsew
rlabel metal1 s 43580 -14 43608 14 4 bl_0_213
port 447 nsew
rlabel metal1 s 43784 -14 43812 14 4 bl_0_214
port 449 nsew
rlabel metal1 s 43988 -14 44016 14 4 bl_0_215
port 451 nsew
rlabel metal1 s 44192 -14 44220 14 4 bl_0_216
port 453 nsew
rlabel metal1 s 44396 -14 44424 14 4 bl_0_217
port 455 nsew
rlabel metal1 s 44600 -14 44628 14 4 bl_0_218
port 457 nsew
rlabel metal1 s 44804 -14 44832 14 4 bl_0_219
port 459 nsew
rlabel metal1 s 45008 -14 45036 14 4 bl_0_220
port 461 nsew
rlabel metal1 s 45212 -14 45240 14 4 bl_0_221
port 463 nsew
rlabel metal1 s 45416 -14 45444 14 4 bl_0_222
port 465 nsew
rlabel metal1 s 45620 -14 45648 14 4 bl_0_223
port 467 nsew
rlabel metal1 s 45824 -14 45852 14 4 bl_0_224
port 469 nsew
rlabel metal1 s 46028 -14 46056 14 4 bl_0_225
port 471 nsew
rlabel metal1 s 46232 -14 46260 14 4 bl_0_226
port 473 nsew
rlabel metal1 s 46436 -14 46464 14 4 bl_0_227
port 475 nsew
rlabel metal1 s 46640 -14 46668 14 4 bl_0_228
port 477 nsew
rlabel metal1 s 46844 -14 46872 14 4 bl_0_229
port 479 nsew
rlabel metal1 s 47048 -14 47076 14 4 bl_0_230
port 481 nsew
rlabel metal1 s 47252 -14 47280 14 4 bl_0_231
port 483 nsew
rlabel metal1 s 47456 -14 47484 14 4 bl_0_232
port 485 nsew
rlabel metal1 s 47660 -14 47688 14 4 bl_0_233
port 487 nsew
rlabel metal1 s 47864 -14 47892 14 4 bl_0_234
port 489 nsew
rlabel metal1 s 48068 -14 48096 14 4 bl_0_235
port 491 nsew
rlabel metal1 s 48272 -14 48300 14 4 bl_0_236
port 493 nsew
rlabel metal1 s 48476 -14 48504 14 4 bl_0_237
port 495 nsew
rlabel metal1 s 48680 -14 48708 14 4 bl_0_238
port 497 nsew
rlabel metal1 s 48884 -14 48912 14 4 bl_0_239
port 499 nsew
rlabel metal1 s 49088 -14 49116 14 4 bl_0_240
port 501 nsew
rlabel metal1 s 49292 -14 49320 14 4 bl_0_241
port 503 nsew
rlabel metal1 s 49496 -14 49524 14 4 bl_0_242
port 505 nsew
rlabel metal1 s 49700 -14 49728 14 4 bl_0_243
port 507 nsew
rlabel metal1 s 49904 -14 49932 14 4 bl_0_244
port 509 nsew
rlabel metal1 s 50108 -14 50136 14 4 bl_0_245
port 511 nsew
rlabel metal1 s 50312 -14 50340 14 4 bl_0_246
port 513 nsew
rlabel metal1 s 50516 -14 50544 14 4 bl_0_247
port 515 nsew
rlabel metal1 s 50720 -14 50748 14 4 bl_0_248
port 517 nsew
rlabel metal1 s 50924 -14 50952 14 4 bl_0_249
port 519 nsew
rlabel metal1 s 51128 -14 51156 14 4 bl_0_250
port 521 nsew
rlabel metal1 s 51332 -14 51360 14 4 bl_0_251
port 523 nsew
rlabel metal1 s 51536 -14 51564 14 4 bl_0_252
port 525 nsew
rlabel metal1 s 51740 -14 51768 14 4 bl_0_253
port 527 nsew
rlabel metal1 s 51944 -14 51972 14 4 bl_0_254
port 529 nsew
rlabel metal1 s 52148 -14 52176 14 4 bl_0_255
port 531 nsew
rlabel metal1 s 52445 368 52473 396 4 precharge_r
port 533 nsew
rlabel metal1 s 52162 2772 52190 2800 4 gnd
port 535 nsew
rlabel metal2 s 230 859 52292 887 4 gnd
port 535 nsew
rlabel metal1 s 114 2772 142 2800 4 gnd
port 535 nsew
rlabel metal2 s 12 -32 40 32 4 vdd
port 537 nsew
<< properties >>
string FIXED_BBOX 0 0 52473 974
<< end >>
