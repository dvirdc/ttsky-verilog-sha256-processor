magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1296 -1277 4216 3436
<< nwell >>
rect -36 1017 2956 2176
<< locali >>
rect 0 2101 2920 2135
rect 64 988 98 1054
rect 196 1004 449 1038
rect 547 1016 817 1050
rect 919 1006 1293 1040
rect 1503 992 1985 1026
rect 2409 992 2443 1026
rect 0 -17 2920 17
use sky130_rom_krom_pinv  sky130_rom_krom_pinv_0
timestamp 1581321264
transform 1 0 368 0 1 0
box -36 -17 404 2176
use sky130_rom_krom_pinv_0  sky130_rom_krom_pinv_0_0
timestamp 1581321264
transform 1 0 736 0 1 0
box -36 -17 512 2176
use sky130_rom_krom_pinv  sky130_rom_krom_pinv_1
timestamp 1581321264
transform 1 0 0 0 1 0
box -36 -17 404 2176
use sky130_rom_krom_pinv_1  sky130_rom_krom_pinv_1_0
timestamp 1581321264
transform 1 0 1212 0 1 0
box -36 -17 728 2176
use sky130_rom_krom_pinv_3  sky130_rom_krom_pinv_3_0
timestamp 1581321264
transform 1 0 1904 0 1 0
box -36 -17 1052 2176
<< labels >>
rlabel locali s 2426 1009 2426 1009 4 Z
port 1 nsew
rlabel locali s 81 1021 81 1021 4 A
port 2 nsew
rlabel locali s 1460 0 1460 0 4 gnd
port 3 nsew
rlabel locali s 1460 2118 1460 2118 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2920 2118
<< end >>
