magic
tech sky130A
magscale 1 2
timestamp 1581582910
<< checkpaint >>
rect -1296 -1277 1674 3946
<< nwell >>
rect -36 1262 414 2686
<< pwell >>
rect 28 25 330 225
<< scnmos >>
rect 114 51 144 199
rect 214 51 244 199
<< scpmos >>
rect 114 2354 144 2578
rect 214 2354 244 2578
<< ndiff >>
rect 54 142 114 199
rect 54 108 62 142
rect 96 108 114 142
rect 54 51 114 108
rect 144 51 214 199
rect 244 142 304 199
rect 244 108 262 142
rect 296 108 304 142
rect 244 51 304 108
<< pdiff >>
rect 54 2483 114 2578
rect 54 2449 62 2483
rect 96 2449 114 2483
rect 54 2354 114 2449
rect 144 2483 214 2578
rect 144 2449 162 2483
rect 196 2449 214 2483
rect 144 2354 214 2449
rect 244 2483 304 2578
rect 244 2449 262 2483
rect 296 2449 304 2483
rect 244 2354 304 2449
<< ndiffc >>
rect 62 108 96 142
rect 262 108 296 142
<< pdiffc >>
rect 62 2449 96 2483
rect 162 2449 196 2483
rect 262 2449 296 2483
<< poly >>
rect 114 2578 144 2604
rect 214 2578 244 2604
rect 114 303 144 2354
rect 214 551 244 2354
rect 196 535 262 551
rect 196 501 212 535
rect 246 501 262 535
rect 196 485 262 501
rect 96 287 162 303
rect 96 253 112 287
rect 146 253 162 287
rect 96 237 162 253
rect 114 199 144 237
rect 214 199 244 485
rect 114 25 144 51
rect 214 25 244 51
<< polycont >>
rect 212 501 246 535
rect 112 253 146 287
<< locali >>
rect 0 2612 378 2646
rect 62 2483 96 2612
rect 62 2433 96 2449
rect 162 2483 196 2499
rect 162 2383 196 2449
rect 262 2483 296 2612
rect 262 2433 296 2449
rect 162 2349 364 2383
rect 212 535 246 551
rect 212 485 246 501
rect 112 287 146 303
rect 112 237 146 253
rect 330 243 364 2349
rect 262 209 364 243
rect 62 142 96 158
rect 62 17 96 108
rect 262 142 296 209
rect 262 92 296 108
rect 0 -17 378 17
<< labels >>
rlabel locali s 347 2366 347 2366 4 Z
port 1 nsew
rlabel locali s 189 0 189 0 4 gnd
port 2 nsew
rlabel locali s 189 2629 189 2629 4 vdd
port 3 nsew
rlabel locali s 129 270 129 270 4 A
port 4 nsew
rlabel locali s 229 518 229 518 4 B
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 378 2382
<< end >>
