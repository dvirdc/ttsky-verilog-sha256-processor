* NGSPICE file created from sky130_rom_krom.ext - technology: sky130A

.subckt sky130_rom_krom_rom_base_one_cell G D S gnd
X0 D G S gnd sky130_fd_pr__nfet_01v8 ad=0.108p pd=1.32u as=0.108p ps=1.32u w=0.36u l=0.15u
.ends

.subckt sky130_rom_krom_rom_base_zero_cell G S gnd
X0 S G S gnd sky130_fd_pr__nfet_01v8 ad=0.216p pd=2.64u as=0p ps=0u w=0.36u l=0.15u
.ends

.subckt sky130_rom_krom_precharge_cell D G vdd
X0 D G vdd vdd sky130_fd_pr__pfet_01v8 ad=0.126p pd=1.44u as=0.126p ps=1.44u w=0.42u l=0.15u
.ends

.subckt sky130_rom_krom_rom_precharge_array_0 pre_bl3_out pre_bl5_out pre_bl6_out
+ pre_bl10_out pre_bl13_out pre_bl17_out pre_bl19_out pre_bl21_out pre_bl22_out pre_bl26_out
+ pre_bl28_out pre_bl29_out pre_bl30_out pre_bl31_out vdd gate pre_bl15_out pre_bl24_out
+ pre_bl8_out pre_bl1_out pre_bl4_out pre_bl2_out pre_bl20_out pre_bl11_out pre_bl18_out
+ pre_bl27_out pre_bl16_out pre_bl9_out pre_bl25_out pre_bl14_out pre_bl7_out pre_bl23_out
+ pre_bl0_out pre_bl12_out
Xsky130_rom_krom_precharge_cell_2 pre_bl29_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_3 pre_bl28_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_4 pre_bl27_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_5 pre_bl26_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_6 pre_bl25_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_7 pre_bl24_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_8 pre_bl23_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_9 pre_bl22_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_30 pre_bl1_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_20 pre_bl11_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_31 pre_bl0_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_10 pre_bl21_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_11 pre_bl20_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_21 pre_bl10_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_22 pre_bl9_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_12 pre_bl19_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_23 pre_bl8_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_13 pre_bl18_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_24 pre_bl7_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_14 pre_bl17_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_25 pre_bl6_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_15 pre_bl16_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_26 pre_bl5_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_16 pre_bl15_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_27 pre_bl4_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_17 pre_bl14_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_28 pre_bl3_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_18 pre_bl13_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_29 pre_bl2_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_19 pre_bl12_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_0 pre_bl31_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_1 pre_bl30_out gate vdd sky130_rom_krom_precharge_cell
.ends

.subckt sky130_rom_krom_rom_row_decode_array bl_0_0 bl_0_1 bl_0_2 bl_0_3 bl_0_4 bl_0_5
+ bl_0_6 bl_0_7 bl_0_8 bl_0_9 bl_0_10 bl_0_11 bl_0_12 bl_0_13 bl_0_14 bl_0_15 bl_0_16
+ bl_0_17 bl_0_18 bl_0_19 bl_0_20 bl_0_21 bl_0_22 bl_0_23 bl_0_25 bl_0_26 bl_0_27
+ bl_0_28 bl_0_29 bl_0_30 bl_0_31 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_9 gnd precharge wl_0_0 vdd wl_0_8 bl_0_24
Xsky130_rom_krom_rom_base_one_cell_94 wl_0_6 sky130_rom_krom_rom_base_one_cell_94/D
+ sky130_rom_krom_rom_base_one_cell_94/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_72 wl_0_7 sky130_rom_krom_rom_base_one_cell_72/D
+ sky130_rom_krom_rom_base_one_cell_72/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_83 wl_0_6 sky130_rom_krom_rom_base_one_cell_83/D
+ sky130_rom_krom_rom_base_one_cell_83/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_61 wl_0_8 sky130_rom_krom_rom_base_one_cell_61/D
+ sky130_rom_krom_rom_base_one_cell_93/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_50 wl_0_8 sky130_rom_krom_rom_base_one_cell_5/S
+ sky130_rom_krom_rom_base_one_cell_67/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_95 wl_0_6 sky130_rom_krom_rom_base_one_cell_95/D
+ sky130_rom_krom_rom_base_one_cell_95/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_73 wl_0_7 sky130_rom_krom_rom_base_one_cell_73/D
+ sky130_rom_krom_rom_base_one_cell_73/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_84 wl_0_6 sky130_rom_krom_rom_base_one_cell_84/D
+ sky130_rom_krom_rom_base_one_cell_84/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_62 wl_0_8 sky130_rom_krom_rom_base_one_cell_62/D
+ sky130_rom_krom_rom_base_one_cell_79/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_51 wl_0_8 sky130_rom_krom_rom_base_one_cell_7/S
+ sky130_rom_krom_rom_base_one_cell_83/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_40 wl_0_9 sky130_rom_krom_rom_base_one_cell_40/D
+ sky130_rom_krom_rom_base_one_cell_72/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_96 wl_0_5 sky130_rom_krom_rom_base_one_cell_96/D
+ sky130_rom_krom_rom_base_one_cell_96/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_74 wl_0_7 sky130_rom_krom_rom_base_one_cell_74/D
+ sky130_rom_krom_rom_base_one_cell_74/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_85 wl_0_6 sky130_rom_krom_rom_base_one_cell_85/D
+ sky130_rom_krom_rom_base_one_cell_85/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_63 wl_0_8 sky130_rom_krom_rom_base_one_cell_63/D
+ sky130_rom_krom_rom_base_one_cell_95/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_52 wl_0_8 sky130_rom_krom_rom_base_one_cell_9/S
+ sky130_rom_krom_rom_base_one_cell_69/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_30 precharge gnd sky130_rom_krom_rom_base_one_cell_47/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_41 wl_0_9 sky130_rom_krom_rom_base_one_cell_41/D
+ sky130_rom_krom_rom_base_one_cell_88/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_97 wl_0_5 sky130_rom_krom_rom_base_one_cell_97/D
+ sky130_rom_krom_rom_base_one_cell_97/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_75 wl_0_7 sky130_rom_krom_rom_base_one_cell_75/D
+ sky130_rom_krom_rom_base_one_cell_75/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_86 wl_0_6 sky130_rom_krom_rom_base_one_cell_86/D
+ sky130_rom_krom_rom_base_one_cell_86/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_64 wl_0_7 sky130_rom_krom_rom_base_one_cell_64/D
+ sky130_rom_krom_rom_base_one_cell_96/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_53 wl_0_8 sky130_rom_krom_rom_base_zero_cell_5/S
+ sky130_rom_krom_rom_base_one_cell_85/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_31 precharge gnd sky130_rom_krom_rom_base_one_cell_63/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_20 precharge gnd sky130_rom_krom_rom_base_one_cell_42/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_42 wl_0_9 sky130_rom_krom_rom_base_one_cell_42/D
+ sky130_rom_krom_rom_base_one_cell_74/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_32 wl_0_9 sky130_rom_krom_rom_base_one_cell_0/S
+ sky130_rom_krom_rom_base_one_cell_64/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_98 wl_0_5 sky130_rom_krom_rom_base_one_cell_98/D
+ sky130_rom_krom_rom_base_one_cell_98/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_76 wl_0_7 sky130_rom_krom_rom_base_one_cell_76/D
+ sky130_rom_krom_rom_base_one_cell_76/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_87 wl_0_6 sky130_rom_krom_rom_base_one_cell_87/D
+ sky130_rom_krom_rom_base_one_cell_87/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_65 wl_0_7 sky130_rom_krom_rom_base_one_cell_65/D
+ sky130_rom_krom_rom_base_one_cell_97/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_54 wl_0_8 sky130_rom_krom_rom_base_zero_cell_6/S
+ sky130_rom_krom_rom_base_one_cell_71/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_21 precharge gnd sky130_rom_krom_rom_base_one_cell_58/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_43 wl_0_9 sky130_rom_krom_rom_base_one_cell_43/D
+ sky130_rom_krom_rom_base_one_cell_90/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_10 precharge gnd sky130_rom_krom_rom_base_one_cell_37/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_190 wl_0_0 sky130_rom_krom_rom_base_one_cell_190/D
+ bl_0_1 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_33 wl_0_9 sky130_rom_krom_rom_base_one_cell_2/S
+ sky130_rom_krom_rom_base_one_cell_80/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_99 wl_0_5 sky130_rom_krom_rom_base_one_cell_99/D
+ sky130_rom_krom_rom_base_one_cell_99/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_77 wl_0_7 sky130_rom_krom_rom_base_one_cell_77/D
+ sky130_rom_krom_rom_base_one_cell_77/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_88 wl_0_6 sky130_rom_krom_rom_base_one_cell_88/D
+ sky130_rom_krom_rom_base_one_cell_88/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_66 wl_0_7 sky130_rom_krom_rom_base_one_cell_66/D
+ sky130_rom_krom_rom_base_one_cell_66/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_55 wl_0_8 sky130_rom_krom_rom_base_zero_cell_7/S
+ sky130_rom_krom_rom_base_one_cell_87/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_44 wl_0_9 sky130_rom_krom_rom_base_one_cell_44/D
+ sky130_rom_krom_rom_base_one_cell_76/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_22 precharge gnd sky130_rom_krom_rom_base_one_cell_43/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_11 precharge gnd sky130_rom_krom_rom_base_zero_cell_5/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_180 wl_0_0 sky130_rom_krom_rom_base_one_cell_180/D
+ bl_0_11 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_191 wl_0_0 sky130_rom_krom_rom_base_one_cell_191/D
+ bl_0_0 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_34 wl_0_9 sky130_rom_krom_rom_base_one_cell_4/S
+ sky130_rom_krom_rom_base_one_cell_66/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_78 wl_0_7 sky130_rom_krom_rom_base_one_cell_78/D
+ sky130_rom_krom_rom_base_one_cell_78/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_89 wl_0_6 sky130_rom_krom_rom_base_one_cell_89/D
+ sky130_rom_krom_rom_base_one_cell_89/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_67 wl_0_7 sky130_rom_krom_rom_base_one_cell_67/D
+ sky130_rom_krom_rom_base_one_cell_67/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_56 wl_0_8 sky130_rom_krom_rom_base_zero_cell_8/S
+ sky130_rom_krom_rom_base_one_cell_73/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_45 wl_0_9 sky130_rom_krom_rom_base_one_cell_45/D
+ sky130_rom_krom_rom_base_one_cell_92/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_23 precharge gnd sky130_rom_krom_rom_base_one_cell_59/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_12 precharge gnd sky130_rom_krom_rom_base_one_cell_38/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_0 precharge gnd sky130_rom_krom_rom_base_one_cell_0/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_170 wl_0_1 sky130_rom_krom_rom_base_one_cell_170/D
+ bl_0_21 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_181 wl_0_0 sky130_rom_krom_rom_base_one_cell_181/D
+ bl_0_10 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_13 precharge gnd sky130_rom_krom_rom_base_zero_cell_6/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_35 wl_0_9 sky130_rom_krom_rom_base_one_cell_6/S
+ sky130_rom_krom_rom_base_one_cell_82/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_79 wl_0_7 sky130_rom_krom_rom_base_one_cell_79/D
+ sky130_rom_krom_rom_base_one_cell_79/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_68 wl_0_7 sky130_rom_krom_rom_base_one_cell_68/D
+ sky130_rom_krom_rom_base_one_cell_68/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_57 wl_0_8 sky130_rom_krom_rom_base_zero_cell_9/S
+ sky130_rom_krom_rom_base_one_cell_89/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_46 wl_0_9 sky130_rom_krom_rom_base_one_cell_46/D
+ sky130_rom_krom_rom_base_one_cell_78/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_24 precharge gnd sky130_rom_krom_rom_base_one_cell_44/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1 precharge gnd sky130_rom_krom_rom_base_one_cell_1/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_160 wl_0_1 sky130_rom_krom_rom_base_one_cell_160/D
+ bl_0_31 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_171 wl_0_1 sky130_rom_krom_rom_base_one_cell_171/D
+ bl_0_20 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_182 wl_0_0 sky130_rom_krom_rom_base_one_cell_182/D
+ bl_0_9 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_0 wl_0_9 sky130_rom_krom_rom_base_one_cell_1/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_36 wl_0_9 sky130_rom_krom_rom_base_one_cell_8/S
+ sky130_rom_krom_rom_base_one_cell_68/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_69 wl_0_7 sky130_rom_krom_rom_base_one_cell_69/D
+ sky130_rom_krom_rom_base_one_cell_69/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_58 wl_0_8 sky130_rom_krom_rom_base_one_cell_58/D
+ sky130_rom_krom_rom_base_one_cell_75/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_47 wl_0_9 sky130_rom_krom_rom_base_one_cell_47/D
+ sky130_rom_krom_rom_base_one_cell_94/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_25 precharge gnd sky130_rom_krom_rom_base_one_cell_60/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_14 precharge gnd sky130_rom_krom_rom_base_one_cell_39/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_2 precharge gnd sky130_rom_krom_rom_base_one_cell_2/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_90 wl_0_4 sky130_rom_krom_rom_base_zero_cell_90/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_150 wl_0_2 sky130_rom_krom_rom_base_one_cell_150/D
+ sky130_rom_krom_rom_base_one_cell_174/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_161 wl_0_1 sky130_rom_krom_rom_base_one_cell_161/D
+ bl_0_30 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_172 wl_0_1 sky130_rom_krom_rom_base_one_cell_172/D
+ bl_0_19 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_183 wl_0_0 sky130_rom_krom_rom_base_one_cell_183/D
+ bl_0_8 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1 wl_0_9 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_precharge_array_0_0 bl_0_3 bl_0_5 bl_0_6 bl_0_10 bl_0_13 bl_0_17
+ bl_0_19 bl_0_21 bl_0_22 bl_0_26 bl_0_28 bl_0_29 bl_0_30 bl_0_31 vdd precharge bl_0_15
+ bl_0_24 bl_0_8 bl_0_1 bl_0_4 bl_0_2 bl_0_20 bl_0_11 bl_0_18 bl_0_27 bl_0_16 bl_0_9
+ bl_0_25 bl_0_14 bl_0_7 bl_0_23 bl_0_0 bl_0_12 sky130_rom_krom_rom_precharge_array_0
Xsky130_rom_krom_rom_base_one_cell_59 wl_0_8 sky130_rom_krom_rom_base_one_cell_59/D
+ sky130_rom_krom_rom_base_one_cell_91/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_48 wl_0_8 sky130_rom_krom_rom_base_one_cell_1/S
+ sky130_rom_krom_rom_base_one_cell_65/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_26 precharge gnd sky130_rom_krom_rom_base_one_cell_45/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_15 precharge gnd sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_37 wl_0_9 sky130_rom_krom_rom_base_one_cell_37/D
+ sky130_rom_krom_rom_base_one_cell_84/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_91 wl_0_4 sky130_rom_krom_rom_base_zero_cell_91/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_80 wl_0_4 sky130_rom_krom_rom_base_one_cell_96/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_3 precharge gnd sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_151 wl_0_2 sky130_rom_krom_rom_base_one_cell_151/D
+ sky130_rom_krom_rom_base_one_cell_175/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_162 wl_0_1 sky130_rom_krom_rom_base_one_cell_162/D
+ bl_0_29 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_173 wl_0_1 sky130_rom_krom_rom_base_one_cell_173/D
+ bl_0_18 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_184 wl_0_0 sky130_rom_krom_rom_base_one_cell_184/D
+ bl_0_7 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_140 wl_0_3 sky130_rom_krom_rom_base_one_cell_140/D
+ sky130_rom_krom_rom_base_one_cell_180/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_2 wl_0_9 sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_49 wl_0_8 sky130_rom_krom_rom_base_one_cell_3/S
+ sky130_rom_krom_rom_base_one_cell_81/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_27 precharge gnd sky130_rom_krom_rom_base_one_cell_61/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_16 precharge gnd sky130_rom_krom_rom_base_one_cell_40/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_38 wl_0_9 sky130_rom_krom_rom_base_one_cell_38/D
+ sky130_rom_krom_rom_base_one_cell_70/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_92 wl_0_4 sky130_rom_krom_rom_base_zero_cell_92/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_81 wl_0_4 sky130_rom_krom_rom_base_one_cell_97/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_70 wl_0_5 sky130_rom_krom_rom_base_one_cell_86/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_4 precharge gnd sky130_rom_krom_rom_base_one_cell_4/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_152 wl_0_2 sky130_rom_krom_rom_base_zero_cell_92/S
+ sky130_rom_krom_rom_base_one_cell_184/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_163 wl_0_1 sky130_rom_krom_rom_base_one_cell_163/D
+ bl_0_28 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_174 wl_0_1 sky130_rom_krom_rom_base_one_cell_174/D
+ bl_0_17 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_185 wl_0_0 sky130_rom_krom_rom_base_one_cell_185/D
+ bl_0_6 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_141 wl_0_3 sky130_rom_krom_rom_base_one_cell_141/D
+ sky130_rom_krom_rom_base_one_cell_181/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_130 wl_0_3 sky130_rom_krom_rom_base_one_cell_98/S
+ sky130_rom_krom_rom_base_one_cell_162/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_3 wl_0_9 sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_28 precharge gnd sky130_rom_krom_rom_base_one_cell_46/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_17 precharge gnd sky130_rom_krom_rom_base_zero_cell_8/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_39 wl_0_9 sky130_rom_krom_rom_base_one_cell_39/D
+ sky130_rom_krom_rom_base_one_cell_86/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_93 wl_0_4 sky130_rom_krom_rom_base_zero_cell_93/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_82 wl_0_4 sky130_rom_krom_rom_base_one_cell_98/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_71 wl_0_5 sky130_rom_krom_rom_base_one_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_60 wl_0_6 sky130_rom_krom_rom_base_one_cell_76/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_5 precharge gnd sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_153 wl_0_2 sky130_rom_krom_rom_base_zero_cell_93/S
+ sky130_rom_krom_rom_base_one_cell_185/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_164 wl_0_1 sky130_rom_krom_rom_base_one_cell_164/D
+ bl_0_27 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_175 wl_0_1 sky130_rom_krom_rom_base_one_cell_175/D
+ bl_0_16 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_186 wl_0_0 sky130_rom_krom_rom_base_one_cell_186/D
+ bl_0_5 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_142 wl_0_3 sky130_rom_krom_rom_base_one_cell_142/D
+ sky130_rom_krom_rom_base_one_cell_182/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_120 wl_0_4 sky130_rom_krom_rom_base_one_cell_74/S
+ sky130_rom_krom_rom_base_one_cell_140/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_131 wl_0_3 sky130_rom_krom_rom_base_one_cell_99/S
+ sky130_rom_krom_rom_base_one_cell_163/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_4 wl_0_9 sky130_rom_krom_rom_base_one_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_29 precharge gnd sky130_rom_krom_rom_base_one_cell_62/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_18 precharge gnd sky130_rom_krom_rom_base_one_cell_41/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_72 wl_0_5 sky130_rom_krom_rom_base_one_cell_74/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_61 wl_0_6 sky130_rom_krom_rom_base_one_cell_77/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_50 wl_0_6 sky130_rom_krom_rom_base_one_cell_66/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_6 precharge gnd sky130_rom_krom_rom_base_one_cell_6/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_94 wl_0_4 sky130_rom_krom_rom_base_zero_cell_94/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_83 wl_0_4 sky130_rom_krom_rom_base_one_cell_99/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_154 wl_0_2 sky130_rom_krom_rom_base_zero_cell_94/S
+ sky130_rom_krom_rom_base_one_cell_186/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_165 wl_0_1 sky130_rom_krom_rom_base_one_cell_165/D
+ bl_0_26 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_176 wl_0_0 sky130_rom_krom_rom_base_one_cell_176/D
+ bl_0_15 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_187 wl_0_0 sky130_rom_krom_rom_base_one_cell_187/D
+ bl_0_4 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_143 wl_0_3 sky130_rom_krom_rom_base_one_cell_143/D
+ sky130_rom_krom_rom_base_one_cell_183/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_121 wl_0_4 sky130_rom_krom_rom_base_one_cell_75/S
+ sky130_rom_krom_rom_base_one_cell_141/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_132 wl_0_3 sky130_rom_krom_rom_base_one_cell_132/D
+ sky130_rom_krom_rom_base_one_cell_164/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_110 wl_0_5 sky130_rom_krom_rom_base_one_cell_92/S
+ sky130_rom_krom_rom_base_zero_cell_94/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_5 wl_0_9 sky130_rom_krom_rom_base_zero_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_19 precharge gnd sky130_rom_krom_rom_base_zero_cell_9/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_7 precharge gnd sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_95 wl_0_4 sky130_rom_krom_rom_base_zero_cell_95/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_84 wl_0_4 sky130_rom_krom_rom_base_zero_cell_96/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_73 wl_0_5 sky130_rom_krom_rom_base_one_cell_75/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_62 wl_0_6 sky130_rom_krom_rom_base_one_cell_78/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_40 wl_0_7 sky130_rom_krom_rom_base_one_cell_88/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_51 wl_0_6 sky130_rom_krom_rom_base_one_cell_67/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_155 wl_0_2 sky130_rom_krom_rom_base_zero_cell_95/S
+ sky130_rom_krom_rom_base_one_cell_187/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_166 wl_0_1 sky130_rom_krom_rom_base_one_cell_166/D
+ bl_0_25 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_177 wl_0_0 sky130_rom_krom_rom_base_one_cell_177/D
+ bl_0_14 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_188 wl_0_0 sky130_rom_krom_rom_base_one_cell_188/D
+ bl_0_3 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_144 wl_0_2 sky130_rom_krom_rom_base_zero_cell_96/S
+ sky130_rom_krom_rom_base_one_cell_168/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_122 wl_0_4 sky130_rom_krom_rom_base_one_cell_90/S
+ sky130_rom_krom_rom_base_one_cell_142/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_133 wl_0_3 sky130_rom_krom_rom_base_one_cell_133/D
+ sky130_rom_krom_rom_base_one_cell_165/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_111 wl_0_5 sky130_rom_krom_rom_base_one_cell_93/S
+ sky130_rom_krom_rom_base_zero_cell_95/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_100 wl_0_5 sky130_rom_krom_rom_base_one_cell_68/S
+ sky130_rom_krom_rom_base_zero_cell_96/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_6 wl_0_9 sky130_rom_krom_rom_base_zero_cell_6/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_85 wl_0_4 sky130_rom_krom_rom_base_zero_cell_97/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_96 wl_0_3 sky130_rom_krom_rom_base_zero_cell_96/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_74 wl_0_5 sky130_rom_krom_rom_base_one_cell_90/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_63 wl_0_6 sky130_rom_krom_rom_base_one_cell_79/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_41 wl_0_7 sky130_rom_krom_rom_base_one_cell_89/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_52 wl_0_6 sky130_rom_krom_rom_base_one_cell_68/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_30 wl_0_8 sky130_rom_krom_rom_base_one_cell_78/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_8 precharge gnd sky130_rom_krom_rom_base_one_cell_8/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_123 wl_0_4 sky130_rom_krom_rom_base_one_cell_91/S
+ sky130_rom_krom_rom_base_one_cell_143/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_134 wl_0_3 sky130_rom_krom_rom_base_one_cell_134/D
+ sky130_rom_krom_rom_base_one_cell_166/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_112 wl_0_4 sky130_rom_krom_rom_base_one_cell_66/S
+ sky130_rom_krom_rom_base_one_cell_132/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_101 wl_0_5 sky130_rom_krom_rom_base_one_cell_69/S
+ sky130_rom_krom_rom_base_zero_cell_97/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_156 wl_0_2 sky130_rom_krom_rom_base_one_cell_156/D
+ sky130_rom_krom_rom_base_one_cell_188/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_167 wl_0_1 sky130_rom_krom_rom_base_one_cell_167/D
+ bl_0_24 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_178 wl_0_0 sky130_rom_krom_rom_base_one_cell_178/D
+ bl_0_13 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_189 wl_0_0 sky130_rom_krom_rom_base_one_cell_189/D
+ bl_0_2 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_145 wl_0_2 sky130_rom_krom_rom_base_zero_cell_97/S
+ sky130_rom_krom_rom_base_one_cell_169/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_7 wl_0_9 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_86 wl_0_4 sky130_rom_krom_rom_base_zero_cell_98/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_97 wl_0_3 sky130_rom_krom_rom_base_zero_cell_97/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_75 wl_0_5 sky130_rom_krom_rom_base_one_cell_91/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_64 wl_0_5 sky130_rom_krom_rom_base_one_cell_66/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_42 wl_0_7 sky130_rom_krom_rom_base_one_cell_90/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_53 wl_0_6 sky130_rom_krom_rom_base_one_cell_69/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_31 wl_0_8 sky130_rom_krom_rom_base_one_cell_94/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_20 wl_0_8 sky130_rom_krom_rom_base_one_cell_68/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_9 precharge gnd sky130_rom_krom_rom_base_one_cell_9/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_157 wl_0_2 sky130_rom_krom_rom_base_one_cell_157/D
+ sky130_rom_krom_rom_base_one_cell_189/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_168 wl_0_1 sky130_rom_krom_rom_base_one_cell_168/D
+ bl_0_23 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_179 wl_0_0 sky130_rom_krom_rom_base_one_cell_179/D
+ bl_0_12 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_146 wl_0_2 sky130_rom_krom_rom_base_zero_cell_98/S
+ sky130_rom_krom_rom_base_one_cell_170/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_124 wl_0_4 sky130_rom_krom_rom_base_one_cell_78/S
+ sky130_rom_krom_rom_base_one_cell_156/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_135 wl_0_3 sky130_rom_krom_rom_base_one_cell_135/D
+ sky130_rom_krom_rom_base_one_cell_167/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_113 wl_0_4 sky130_rom_krom_rom_base_one_cell_67/S
+ sky130_rom_krom_rom_base_one_cell_133/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_102 wl_0_5 sky130_rom_krom_rom_base_one_cell_84/S
+ sky130_rom_krom_rom_base_zero_cell_98/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_8 wl_0_9 sky130_rom_krom_rom_base_zero_cell_8/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_87 wl_0_4 sky130_rom_krom_rom_base_zero_cell_99/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_98 wl_0_3 sky130_rom_krom_rom_base_zero_cell_98/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_76 wl_0_5 sky130_rom_krom_rom_base_one_cell_78/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_65 wl_0_5 sky130_rom_krom_rom_base_one_cell_67/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_43 wl_0_7 sky130_rom_krom_rom_base_one_cell_91/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_54 wl_0_6 sky130_rom_krom_rom_base_one_cell_70/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_32 wl_0_7 sky130_rom_krom_rom_base_one_cell_80/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_21 wl_0_8 sky130_rom_krom_rom_base_one_cell_84/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_10 wl_0_9 sky130_rom_krom_rom_base_one_cell_58/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_158 wl_0_2 sky130_rom_krom_rom_base_one_cell_158/D
+ sky130_rom_krom_rom_base_one_cell_190/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_169 wl_0_1 sky130_rom_krom_rom_base_one_cell_169/D
+ bl_0_22 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_147 wl_0_2 sky130_rom_krom_rom_base_zero_cell_99/S
+ sky130_rom_krom_rom_base_one_cell_171/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_125 wl_0_4 sky130_rom_krom_rom_base_one_cell_79/S
+ sky130_rom_krom_rom_base_one_cell_157/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_136 wl_0_3 sky130_rom_krom_rom_base_zero_cell_88/S
+ sky130_rom_krom_rom_base_one_cell_176/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_114 wl_0_4 sky130_rom_krom_rom_base_one_cell_82/S
+ sky130_rom_krom_rom_base_one_cell_134/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_103 wl_0_5 sky130_rom_krom_rom_base_one_cell_85/S
+ sky130_rom_krom_rom_base_zero_cell_99/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_9 wl_0_9 sky130_rom_krom_rom_base_zero_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_88 wl_0_4 sky130_rom_krom_rom_base_zero_cell_88/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_77 wl_0_5 sky130_rom_krom_rom_base_one_cell_79/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_66 wl_0_5 sky130_rom_krom_rom_base_one_cell_82/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_44 wl_0_7 sky130_rom_krom_rom_base_one_cell_92/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_55 wl_0_6 sky130_rom_krom_rom_base_one_cell_71/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_33 wl_0_7 sky130_rom_krom_rom_base_one_cell_81/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_22 wl_0_8 sky130_rom_krom_rom_base_one_cell_70/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_11 wl_0_9 sky130_rom_krom_rom_base_one_cell_59/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_99 wl_0_3 sky130_rom_krom_rom_base_zero_cell_99/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_159 wl_0_2 sky130_rom_krom_rom_base_one_cell_159/D
+ sky130_rom_krom_rom_base_one_cell_191/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_148 wl_0_2 sky130_rom_krom_rom_base_one_cell_148/D
+ sky130_rom_krom_rom_base_one_cell_172/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_126 wl_0_4 sky130_rom_krom_rom_base_one_cell_94/S
+ sky130_rom_krom_rom_base_one_cell_158/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_137 wl_0_3 sky130_rom_krom_rom_base_zero_cell_89/S
+ sky130_rom_krom_rom_base_one_cell_177/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_115 wl_0_4 sky130_rom_krom_rom_base_one_cell_83/S
+ sky130_rom_krom_rom_base_one_cell_135/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_104 wl_0_5 sky130_rom_krom_rom_base_one_cell_72/S
+ sky130_rom_krom_rom_base_zero_cell_88/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_89 wl_0_4 sky130_rom_krom_rom_base_zero_cell_89/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_78 wl_0_5 sky130_rom_krom_rom_base_one_cell_94/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_67 wl_0_5 sky130_rom_krom_rom_base_one_cell_83/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_45 wl_0_7 sky130_rom_krom_rom_base_one_cell_93/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_56 wl_0_6 sky130_rom_krom_rom_base_one_cell_72/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_34 wl_0_7 sky130_rom_krom_rom_base_one_cell_82/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_23 wl_0_8 sky130_rom_krom_rom_base_one_cell_86/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_12 wl_0_9 sky130_rom_krom_rom_base_one_cell_60/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_149 wl_0_2 sky130_rom_krom_rom_base_one_cell_149/D
+ sky130_rom_krom_rom_base_one_cell_173/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_127 wl_0_4 sky130_rom_krom_rom_base_one_cell_95/S
+ sky130_rom_krom_rom_base_one_cell_159/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_138 wl_0_3 sky130_rom_krom_rom_base_zero_cell_90/S
+ sky130_rom_krom_rom_base_one_cell_178/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_116 wl_0_4 sky130_rom_krom_rom_base_one_cell_70/S
+ sky130_rom_krom_rom_base_one_cell_148/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_105 wl_0_5 sky130_rom_krom_rom_base_one_cell_73/S
+ sky130_rom_krom_rom_base_zero_cell_89/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_79 wl_0_5 sky130_rom_krom_rom_base_one_cell_95/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_68 wl_0_5 sky130_rom_krom_rom_base_one_cell_70/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_46 wl_0_7 sky130_rom_krom_rom_base_one_cell_94/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_57 wl_0_6 sky130_rom_krom_rom_base_one_cell_73/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_35 wl_0_7 sky130_rom_krom_rom_base_one_cell_83/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_24 wl_0_8 sky130_rom_krom_rom_base_one_cell_72/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_13 wl_0_9 sky130_rom_krom_rom_base_one_cell_61/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_139 wl_0_3 sky130_rom_krom_rom_base_zero_cell_91/S
+ sky130_rom_krom_rom_base_one_cell_179/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_117 wl_0_4 sky130_rom_krom_rom_base_one_cell_71/S
+ sky130_rom_krom_rom_base_one_cell_149/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_128 wl_0_3 sky130_rom_krom_rom_base_one_cell_96/S
+ sky130_rom_krom_rom_base_one_cell_160/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_106 wl_0_5 sky130_rom_krom_rom_base_one_cell_88/S
+ sky130_rom_krom_rom_base_zero_cell_90/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_69 wl_0_5 sky130_rom_krom_rom_base_one_cell_71/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_47 wl_0_7 sky130_rom_krom_rom_base_one_cell_95/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_58 wl_0_6 sky130_rom_krom_rom_base_one_cell_74/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_36 wl_0_7 sky130_rom_krom_rom_base_one_cell_84/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_25 wl_0_8 sky130_rom_krom_rom_base_one_cell_88/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_14 wl_0_9 sky130_rom_krom_rom_base_one_cell_62/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_150 wl_0_0 bl_0_25 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_118 wl_0_4 sky130_rom_krom_rom_base_one_cell_86/S
+ sky130_rom_krom_rom_base_one_cell_150/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_129 wl_0_3 sky130_rom_krom_rom_base_one_cell_97/S
+ sky130_rom_krom_rom_base_one_cell_161/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_107 wl_0_5 sky130_rom_krom_rom_base_one_cell_89/S
+ sky130_rom_krom_rom_base_zero_cell_91/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_59 wl_0_6 sky130_rom_krom_rom_base_one_cell_75/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_37 wl_0_7 sky130_rom_krom_rom_base_one_cell_85/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_48 wl_0_6 sky130_rom_krom_rom_base_one_cell_96/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_26 wl_0_8 sky130_rom_krom_rom_base_one_cell_74/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_15 wl_0_9 sky130_rom_krom_rom_base_one_cell_63/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_151 wl_0_0 bl_0_24 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_140 wl_0_1 sky130_rom_krom_rom_base_one_cell_188/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_119 wl_0_4 sky130_rom_krom_rom_base_one_cell_87/S
+ sky130_rom_krom_rom_base_one_cell_151/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_108 wl_0_5 sky130_rom_krom_rom_base_one_cell_76/S
+ sky130_rom_krom_rom_base_zero_cell_92/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_38 wl_0_7 sky130_rom_krom_rom_base_one_cell_86/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_49 wl_0_6 sky130_rom_krom_rom_base_one_cell_97/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_27 wl_0_8 sky130_rom_krom_rom_base_one_cell_90/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_16 wl_0_8 sky130_rom_krom_rom_base_one_cell_64/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_152 wl_0_0 bl_0_23 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_130 wl_0_1 sky130_rom_krom_rom_base_one_cell_178/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_141 wl_0_1 sky130_rom_krom_rom_base_one_cell_189/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_109 wl_0_5 sky130_rom_krom_rom_base_one_cell_77/S
+ sky130_rom_krom_rom_base_zero_cell_93/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_39 wl_0_7 sky130_rom_krom_rom_base_one_cell_87/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_28 wl_0_8 sky130_rom_krom_rom_base_one_cell_76/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_17 wl_0_8 sky130_rom_krom_rom_base_one_cell_80/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_120 wl_0_2 sky130_rom_krom_rom_base_one_cell_176/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_153 wl_0_0 bl_0_22 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_131 wl_0_1 sky130_rom_krom_rom_base_one_cell_179/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_142 wl_0_1 sky130_rom_krom_rom_base_one_cell_190/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_29 wl_0_8 sky130_rom_krom_rom_base_one_cell_92/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_18 wl_0_8 sky130_rom_krom_rom_base_one_cell_66/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_121 wl_0_2 sky130_rom_krom_rom_base_one_cell_177/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_154 wl_0_0 bl_0_21 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_132 wl_0_1 sky130_rom_krom_rom_base_one_cell_180/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_143 wl_0_1 sky130_rom_krom_rom_base_one_cell_191/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_110 wl_0_3 sky130_rom_krom_rom_base_one_cell_158/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_19 wl_0_8 sky130_rom_krom_rom_base_one_cell_82/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_122 wl_0_2 sky130_rom_krom_rom_base_one_cell_178/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_144 wl_0_0 bl_0_31 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_155 wl_0_0 bl_0_20 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_133 wl_0_1 sky130_rom_krom_rom_base_one_cell_181/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_111 wl_0_3 sky130_rom_krom_rom_base_one_cell_159/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_100 wl_0_3 sky130_rom_krom_rom_base_one_cell_148/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_123 wl_0_2 sky130_rom_krom_rom_base_one_cell_179/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_145 wl_0_0 bl_0_30 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_156 wl_0_0 bl_0_19 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_134 wl_0_1 sky130_rom_krom_rom_base_one_cell_182/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_112 wl_0_2 sky130_rom_krom_rom_base_one_cell_160/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_101 wl_0_3 sky130_rom_krom_rom_base_one_cell_149/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_124 wl_0_2 sky130_rom_krom_rom_base_one_cell_180/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_146 wl_0_0 bl_0_29 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_157 wl_0_0 bl_0_18 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_135 wl_0_1 sky130_rom_krom_rom_base_one_cell_183/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_113 wl_0_2 sky130_rom_krom_rom_base_one_cell_161/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_102 wl_0_3 sky130_rom_krom_rom_base_one_cell_150/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_125 wl_0_2 sky130_rom_krom_rom_base_one_cell_181/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_147 wl_0_0 bl_0_28 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_158 wl_0_0 bl_0_17 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_136 wl_0_1 sky130_rom_krom_rom_base_one_cell_184/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_114 wl_0_2 sky130_rom_krom_rom_base_one_cell_162/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_103 wl_0_3 sky130_rom_krom_rom_base_one_cell_151/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_126 wl_0_2 sky130_rom_krom_rom_base_one_cell_182/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_148 wl_0_0 bl_0_27 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_159 wl_0_0 bl_0_16 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_137 wl_0_1 sky130_rom_krom_rom_base_one_cell_185/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_115 wl_0_2 sky130_rom_krom_rom_base_one_cell_163/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_104 wl_0_3 sky130_rom_krom_rom_base_zero_cell_92/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_127 wl_0_2 sky130_rom_krom_rom_base_one_cell_183/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_149 wl_0_0 bl_0_26 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_138 wl_0_1 sky130_rom_krom_rom_base_one_cell_186/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_116 wl_0_2 sky130_rom_krom_rom_base_one_cell_164/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_105 wl_0_3 sky130_rom_krom_rom_base_zero_cell_93/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_128 wl_0_1 sky130_rom_krom_rom_base_one_cell_176/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_139 wl_0_1 sky130_rom_krom_rom_base_one_cell_187/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_117 wl_0_2 sky130_rom_krom_rom_base_one_cell_165/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_106 wl_0_3 sky130_rom_krom_rom_base_zero_cell_94/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_90 wl_0_6 sky130_rom_krom_rom_base_one_cell_90/D
+ sky130_rom_krom_rom_base_one_cell_90/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_129 wl_0_1 sky130_rom_krom_rom_base_one_cell_177/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_118 wl_0_2 sky130_rom_krom_rom_base_one_cell_166/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_107 wl_0_3 sky130_rom_krom_rom_base_zero_cell_95/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_91 wl_0_6 sky130_rom_krom_rom_base_one_cell_91/D
+ sky130_rom_krom_rom_base_one_cell_91/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_80 wl_0_6 sky130_rom_krom_rom_base_one_cell_80/D
+ sky130_rom_krom_rom_base_one_cell_98/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_119 wl_0_2 sky130_rom_krom_rom_base_one_cell_167/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_108 wl_0_3 sky130_rom_krom_rom_base_one_cell_156/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_92 wl_0_6 sky130_rom_krom_rom_base_one_cell_92/D
+ sky130_rom_krom_rom_base_one_cell_92/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_70 wl_0_7 sky130_rom_krom_rom_base_one_cell_70/D
+ sky130_rom_krom_rom_base_one_cell_70/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_81 wl_0_6 sky130_rom_krom_rom_base_one_cell_81/D
+ sky130_rom_krom_rom_base_one_cell_99/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_109 wl_0_3 sky130_rom_krom_rom_base_one_cell_157/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_93 wl_0_6 sky130_rom_krom_rom_base_one_cell_93/D
+ sky130_rom_krom_rom_base_one_cell_93/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_71 wl_0_7 sky130_rom_krom_rom_base_one_cell_71/D
+ sky130_rom_krom_rom_base_one_cell_71/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_82 wl_0_6 sky130_rom_krom_rom_base_one_cell_82/D
+ sky130_rom_krom_rom_base_one_cell_82/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_60 wl_0_8 sky130_rom_krom_rom_base_one_cell_60/D
+ sky130_rom_krom_rom_base_one_cell_77/D gnd sky130_rom_krom_rom_base_one_cell
.ends

.subckt sky130_rom_krom_inv_array_mod A Z vdd gnd w_504_0#
X0 vdd A Z w_504_0# sky130_fd_pr__pfet_01v8 ad=0.9p pd=6.6u as=0.9p ps=6.6u w=3u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.222p pd=2.08u as=0.222p ps=2.08u w=0.74u l=0.15u
.ends

.subckt sky130_fd_bd_sram__openram_sp_nand2_dec A B Z vdd gnd
X0 vdd B Z vdd sky130_fd_pr__pfet_01v8 ad=0.336p pd=2.84u as=0.6776p ps=5.69u w=1.12u l=0.15u
X1 a_174_144# B gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1554p pd=1.9u as=0.222p ps=2.08u w=0.74u l=0.15u
X2 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12u l=0.15u
X3 Z A a_174_144# gnd sky130_fd_pr__nfet_01v8 ad=0.2701p pd=2.21u as=0p ps=0u w=0.74u l=0.15u
.ends

.subckt sky130_rom_krom_rom_address_control_buf A_in A_out Abar_out clk vdd_uq0 vdd_uq1
+ vdd gnd
Xsky130_rom_krom_inv_array_mod_0 A_in sky130_rom_krom_inv_array_mod_0/Z vdd_uq1 gnd
+ vdd_uq1 sky130_rom_krom_inv_array_mod
Xsky130_fd_bd_sram__openram_sp_nand2_dec_0 clk A_out Abar_out vdd gnd sky130_fd_bd_sram__openram_sp_nand2_dec
Xsky130_fd_bd_sram__openram_sp_nand2_dec_1 clk sky130_rom_krom_inv_array_mod_0/Z A_out
+ vdd_uq0 gnd sky130_fd_bd_sram__openram_sp_nand2_dec
.ends

.subckt sky130_rom_krom_rom_address_control_array A0_in A1_in A2_in A3_in A4_in A0_out
+ A1_out A2_out A3_out A4_out Abar0_out Abar1_out Abar3_out Abar4_out vdd vdd_uq0
+ vdd_uq1 Abar2_out gnd clk
Xsky130_rom_krom_rom_address_control_buf_0 A4_in A4_out Abar4_out clk vdd vdd_uq0
+ vdd_uq1 gnd sky130_rom_krom_rom_address_control_buf
Xsky130_rom_krom_rom_address_control_buf_2 A2_in A2_out Abar2_out clk vdd vdd_uq0
+ vdd_uq1 gnd sky130_rom_krom_rom_address_control_buf
Xsky130_rom_krom_rom_address_control_buf_1 A3_in A3_out Abar3_out clk vdd vdd_uq0
+ vdd_uq1 gnd sky130_rom_krom_rom_address_control_buf
Xsky130_rom_krom_rom_address_control_buf_3 A1_in A1_out Abar1_out clk vdd vdd_uq0
+ vdd_uq1 gnd sky130_rom_krom_rom_address_control_buf
Xsky130_rom_krom_rom_address_control_buf_4 A0_in A0_out Abar0_out clk vdd vdd_uq0
+ vdd_uq1 gnd sky130_rom_krom_rom_address_control_buf
.ends

.subckt sky130_rom_krom_pinv_dec_1 A Z vdd gnd w_956_n45#
X0 vdd A Z w_956_n45# sky130_fd_pr__pfet_01v8 ad=2.1p pd=14.6u as=2.1p ps=14.6u w=7u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.9p pd=6.6u as=0.9p ps=6.6u w=3u l=0.15u
.ends

.subckt sky130_rom_krom_pinv_dec_0 A Z vdd gnd w_504_n45#
X0 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.222p pd=2.08u as=0.222p ps=2.08u w=0.74u l=0.15u
X1 vdd A Z w_504_n45# sky130_fd_pr__pfet_01v8 ad=0.9p pd=6.6u as=0.9p ps=6.6u w=3u l=0.15u
.ends

.subckt sky130_rom_krom_pbuf_dec Z vdd vdd_uq0 gnd sky130_rom_krom_pinv_dec_1_0/w_956_n45#
+ A sky130_rom_krom_pinv_dec_0_0/w_504_n45#
Xsky130_rom_krom_pinv_dec_1_0 sky130_rom_krom_pinv_dec_1_0/A Z vdd_uq0 gnd sky130_rom_krom_pinv_dec_1_0/w_956_n45#
+ sky130_rom_krom_pinv_dec_1
Xsky130_rom_krom_pinv_dec_0_0 A sky130_rom_krom_pinv_dec_1_0/A vdd gnd sky130_rom_krom_pinv_dec_0_0/w_504_n45#
+ sky130_rom_krom_pinv_dec_0
.ends

.subckt sky130_rom_krom_rom_row_decode_wordline_buffer in_0 in_1 in_2 in_3 in_4 in_6
+ in_7 in_8 in_9 in_10 in_11 in_12 in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20
+ in_21 in_22 in_23 in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 out_0 out_1 out_2
+ out_3 out_4 out_5 out_6 out_7 out_8 out_9 out_10 out_11 out_12 out_13 out_14 out_15
+ out_16 out_17 out_18 out_19 out_20 out_21 out_22 out_23 out_25 out_26 out_27 out_28
+ out_29 out_30 out_31 vdd_uq0 in_5 vdd gnd out_24
Xsky130_rom_krom_pbuf_dec_30 out_1 vdd vdd_uq0 gnd vdd_uq0 in_1 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_20 out_11 vdd vdd_uq0 gnd vdd_uq0 in_11 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_31 out_0 vdd vdd_uq0 gnd vdd_uq0 in_0 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_10 out_21 vdd vdd_uq0 gnd vdd_uq0 in_21 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_21 out_10 vdd vdd_uq0 gnd vdd_uq0 in_10 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_11 out_20 vdd vdd_uq0 gnd vdd_uq0 in_20 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_22 out_9 vdd vdd_uq0 gnd vdd_uq0 in_9 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_12 out_19 vdd vdd_uq0 gnd vdd_uq0 in_19 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_13 out_18 vdd vdd_uq0 gnd vdd_uq0 in_18 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_23 out_8 vdd vdd_uq0 gnd vdd_uq0 in_8 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_24 out_7 vdd vdd_uq0 gnd vdd_uq0 in_7 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_0 out_31 vdd vdd_uq0 gnd vdd_uq0 in_31 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_14 out_17 vdd vdd_uq0 gnd vdd_uq0 in_17 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_25 out_6 vdd vdd_uq0 gnd vdd_uq0 in_6 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_1 out_30 vdd vdd_uq0 gnd vdd_uq0 in_30 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_15 out_16 vdd vdd_uq0 gnd vdd_uq0 in_16 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_26 out_5 vdd vdd_uq0 gnd vdd_uq0 in_5 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_2 out_29 vdd vdd_uq0 gnd vdd_uq0 in_29 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_16 out_15 vdd vdd_uq0 gnd vdd_uq0 in_15 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_27 out_4 vdd vdd_uq0 gnd vdd_uq0 in_4 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_3 out_28 vdd vdd_uq0 gnd vdd_uq0 in_28 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_17 out_14 vdd vdd_uq0 gnd vdd_uq0 in_14 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_28 out_3 vdd vdd_uq0 gnd vdd_uq0 in_3 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_4 out_27 vdd vdd_uq0 gnd vdd_uq0 in_27 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_5 out_26 vdd vdd_uq0 gnd vdd_uq0 in_26 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_18 out_13 vdd vdd_uq0 gnd vdd_uq0 in_13 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_29 out_2 vdd vdd_uq0 gnd vdd_uq0 in_2 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_6 out_25 vdd vdd_uq0 gnd vdd_uq0 in_25 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_19 out_12 vdd vdd_uq0 gnd vdd_uq0 in_12 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_7 out_24 vdd vdd_uq0 gnd vdd_uq0 in_24 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_8 out_23 vdd vdd_uq0 gnd vdd_uq0 in_23 vdd sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_9 out_22 vdd vdd_uq0 gnd vdd_uq0 in_22 vdd sky130_rom_krom_pbuf_dec
.ends

.subckt sky130_rom_krom_rom_row_decode A0 A1 A2 A3 A4 wl_0 wl_1 wl_2 wl_3 wl_4 wl_6
+ wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20
+ wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 clk vdd_uq0 vdd_uq1
+ vdd_uq2 vdd_uq5 vdd_uq6 vdd wl_5 precharge gnd
Xsky130_rom_krom_rom_row_decode_array_0 sky130_rom_krom_rom_row_decode_array_0/bl_0_0
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_1 sky130_rom_krom_rom_row_decode_array_0/bl_0_2
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_3 sky130_rom_krom_rom_row_decode_array_0/bl_0_4
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_5 sky130_rom_krom_rom_row_decode_array_0/bl_0_6
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_7 sky130_rom_krom_rom_row_decode_array_0/bl_0_8
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_9 sky130_rom_krom_rom_row_decode_array_0/bl_0_10
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_11 sky130_rom_krom_rom_row_decode_array_0/bl_0_12
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_13 sky130_rom_krom_rom_row_decode_array_0/bl_0_14
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_15 sky130_rom_krom_rom_row_decode_array_0/bl_0_16
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_17 sky130_rom_krom_rom_row_decode_array_0/bl_0_18
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_19 sky130_rom_krom_rom_row_decode_array_0/bl_0_20
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_21 sky130_rom_krom_rom_row_decode_array_0/bl_0_22
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_23 sky130_rom_krom_rom_row_decode_array_0/bl_0_25
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_26 sky130_rom_krom_rom_row_decode_array_0/bl_0_27
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_28 sky130_rom_krom_rom_row_decode_array_0/bl_0_29
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_30 sky130_rom_krom_rom_row_decode_array_0/bl_0_31
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_1 sky130_rom_krom_rom_row_decode_array_0/wl_0_2
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_3 sky130_rom_krom_rom_row_decode_array_0/wl_0_4
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_5 sky130_rom_krom_rom_row_decode_array_0/wl_0_6
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_7 sky130_rom_krom_rom_row_decode_array_0/wl_0_9
+ gnd precharge sky130_rom_krom_rom_row_decode_array_0/wl_0_0 vdd_uq0 sky130_rom_krom_rom_row_decode_array_0/wl_0_8
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_24 sky130_rom_krom_rom_row_decode_array
Xsky130_rom_krom_rom_address_control_array_0 A0 A1 A2 A3 A4 sky130_rom_krom_rom_row_decode_array_0/wl_0_9
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_7 sky130_rom_krom_rom_row_decode_array_0/wl_0_5
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_3 sky130_rom_krom_rom_row_decode_array_0/wl_0_1
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_8 sky130_rom_krom_rom_row_decode_array_0/wl_0_6
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_2 sky130_rom_krom_rom_row_decode_array_0/wl_0_0
+ vdd_uq1 vdd vdd_uq2 sky130_rom_krom_rom_row_decode_array_0/wl_0_4 gnd clk sky130_rom_krom_rom_address_control_array
Xsky130_rom_krom_rom_row_decode_wordline_buffer_0 sky130_rom_krom_rom_row_decode_array_0/bl_0_0
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_1 sky130_rom_krom_rom_row_decode_array_0/bl_0_2
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_3 sky130_rom_krom_rom_row_decode_array_0/bl_0_4
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_6 sky130_rom_krom_rom_row_decode_array_0/bl_0_7
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_8 sky130_rom_krom_rom_row_decode_array_0/bl_0_9
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_10 sky130_rom_krom_rom_row_decode_array_0/bl_0_11
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_12 sky130_rom_krom_rom_row_decode_array_0/bl_0_13
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_14 sky130_rom_krom_rom_row_decode_array_0/bl_0_15
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_16 sky130_rom_krom_rom_row_decode_array_0/bl_0_17
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_18 sky130_rom_krom_rom_row_decode_array_0/bl_0_19
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_20 sky130_rom_krom_rom_row_decode_array_0/bl_0_21
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_22 sky130_rom_krom_rom_row_decode_array_0/bl_0_23
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_24 sky130_rom_krom_rom_row_decode_array_0/bl_0_25
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_26 sky130_rom_krom_rom_row_decode_array_0/bl_0_27
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_28 sky130_rom_krom_rom_row_decode_array_0/bl_0_29
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_30 sky130_rom_krom_rom_row_decode_array_0/bl_0_31
+ wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14
+ wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_25 wl_26 wl_27 wl_28 wl_29
+ wl_30 wl_31 vdd_uq5 sky130_rom_krom_rom_row_decode_array_0/bl_0_5 vdd_uq6 gnd wl_24
+ sky130_rom_krom_rom_row_decode_wordline_buffer
.ends

.subckt sky130_rom_krom_pinv_dec_4 A Z vdd gnd w_692_n45#
X0 vdd A Z w_692_n45# sky130_fd_pr__pfet_01v8 ad=1.5p pd=10.6u as=1.5p ps=10.6u w=5u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.504p pd=3.96u as=0.504p ps=3.96u w=1.68u l=0.15u
.ends

.subckt sky130_rom_krom_rom_output_buffer in_0 in_1 in_2 in_4 in_5 in_6 in_7 out_0
+ out_1 out_2 out_3 out_4 out_5 out_6 out_7 gnd vdd in_3
Xsky130_rom_krom_pinv_dec_4_0 in_7 out_7 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_1 in_6 out_6 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_2 in_5 out_5 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_3 in_4 out_4 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_4 in_3 out_3 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_5 in_2 out_2 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_6 in_1 out_1 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_7 in_0 out_0 vdd gnd vdd sky130_rom_krom_pinv_dec_4
.ends

.subckt sky130_rom_krom_pinv_2 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34p pd=13.56u as=2.97p ps=19.98u w=3u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X2 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X3 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=4.95p pd=31.98u as=3.9p ps=21.56u w=5u l=0.15u
X4 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X5 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X6 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X7 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
.ends

.subckt sky130_rom_krom_pinv_0 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.2886p pd=2.26u as=0.444p ps=4.16u w=0.74u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0.74u l=0.15u
X2 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0.756p pd=6.24u as=0.4914p ps=3.3u w=1.26u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26u l=0.15u
.ends

.subckt sky130_rom_krom_pinv_1 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.78p pd=4.78u as=1.2p ps=9.2u w=2u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=1.8p pd=13.2u as=1.17p ps=6.78u w=3u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
.ends

.subckt sky130_rom_krom_pinv A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.108p pd=1.32u as=0.108p ps=1.32u w=0.36u l=0.15u
X1 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.336p pd=2.84u as=0.336p ps=2.84u w=1.12u l=0.15u
.ends

.subckt sky130_rom_krom_rom_clock_driver A Z vdd gnd
Xsky130_rom_krom_pinv_2_0 sky130_rom_krom_pinv_2_0/A Z vdd gnd sky130_rom_krom_pinv_2
Xsky130_rom_krom_pinv_0_0 sky130_rom_krom_pinv_0/Z sky130_rom_krom_pinv_1_0/A vdd
+ gnd sky130_rom_krom_pinv_0
Xsky130_rom_krom_pinv_1_0 sky130_rom_krom_pinv_1_0/A sky130_rom_krom_pinv_2_0/A vdd
+ gnd sky130_rom_krom_pinv_1
Xsky130_rom_krom_pinv_0 A sky130_rom_krom_pinv_0/Z vdd gnd sky130_rom_krom_pinv
.ends

.subckt sky130_rom_krom_rom_control_nand A B Z vdd gnd w_n36_1262#
X0 a_144_51# A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.259p pd=2.18u as=0.222p ps=2.08u w=0.74u l=0.15u
X1 vdd B Z w_n36_1262# sky130_fd_pr__pfet_01v8 ad=0.672p pd=5.68u as=0.392p ps=2.94u w=1.12u l=0.15u
X2 Z A vdd w_n36_1262# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12u l=0.15u
X3 Z B a_144_51# gnd sky130_fd_pr__nfet_01v8 ad=0.222p pd=2.08u as=0p ps=0u w=0.74u l=0.15u
.ends

.subckt sky130_rom_krom_pinv_4 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.78p pd=4.78u as=1.2p ps=9.2u w=2u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=3p pd=21.2u as=1.95p ps=10.78u w=5u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
.ends

.subckt sky130_rom_krom_pinv_5 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=5.85p pd=32.34u as=6.9p ps=42.76u w=5u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X2 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X3 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=6.9p pd=42.76u as=5.85p ps=32.34u w=5u l=0.15u
X4 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X5 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X6 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X7 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X8 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X9 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X10 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X11 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
.ends

.subckt sky130_rom_krom_pinv_3 A Z vdd gnd
X0 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=1.2p pd=9.2u as=0.78p ps=4.78u w=2u l=0.15u
X1 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.4914p pd=3.3u as=0.756p ps=6.24u w=1.26u l=0.15u
X3 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26u l=0.15u
.ends

.subckt sky130_rom_krom_rom_precharge_driver A Z vdd gnd
Xsky130_rom_krom_pinv_4_0 sky130_rom_krom_pinv_4_0/A sky130_rom_krom_pinv_5_0/A vdd
+ gnd sky130_rom_krom_pinv_4
Xsky130_rom_krom_pinv_5_0 sky130_rom_krom_pinv_5_0/A Z vdd gnd sky130_rom_krom_pinv_5
Xsky130_rom_krom_pinv_3_0 sky130_rom_krom_pinv_0/Z sky130_rom_krom_pinv_4_0/A vdd
+ gnd sky130_rom_krom_pinv_3
Xsky130_rom_krom_pinv_0 sky130_rom_krom_pinv_1/Z sky130_rom_krom_pinv_0/Z vdd gnd
+ sky130_rom_krom_pinv
Xsky130_rom_krom_pinv_1 A sky130_rom_krom_pinv_1/Z vdd gnd sky130_rom_krom_pinv
.ends

.subckt sky130_rom_krom_rom_control_logic clk_in CS prechrg clk_out vdd gnd
Xsky130_rom_krom_rom_clock_driver_0 clk_in clk_out vdd gnd sky130_rom_krom_rom_clock_driver
Xsky130_rom_krom_rom_control_nand_0 CS clk_out sky130_rom_krom_rom_control_nand_0/Z
+ vdd gnd vdd sky130_rom_krom_rom_control_nand
Xsky130_rom_krom_rom_precharge_driver_0 sky130_rom_krom_rom_control_nand_0/Z prechrg
+ vdd gnd sky130_rom_krom_rom_precharge_driver
.ends

.subckt sky130_rom_krom_rom_column_mux bl bl_out sel gnd
X0 bl_out sel bl gnd sky130_fd_pr__nfet_01v8 ad=0.864p pd=6.36u as=0.864p ps=6.36u w=2.88u l=0.15u
.ends

.subckt sky130_rom_krom_rom_column_mux_array bl_0 bl_1 bl_2 bl_3 bl_4 bl_5 bl_6 bl_8
+ bl_9 bl_11 bl_15 bl_16 bl_17 bl_18 bl_19 bl_22 bl_26 bl_27 bl_28 bl_29 bl_30 bl_37
+ bl_38 bl_39 bl_41 bl_48 bl_49 bl_52 bl_59 bl_62 sel_3 sel_4 sel_5 bl_out_0 bl_out_1
+ bl_out_2 bl_out_3 bl_out_4 bl_out_5 bl_out_6 bl_out_7 gnd bl_24 bl_35 bl_56 bl_33
+ bl_46 bl_14 bl_12 bl_25 bl_20 bl_23 bl_54 bl_36 bl_31 bl_44 bl_57 bl_47 bl_42 bl_60
+ bl_50 bl_63 bl_53 bl_7 bl_10 bl_13 bl_21 bl_34 bl_55 bl_32 bl_58 bl_45 bl_40 bl_43
+ bl_61 bl_51 sel_7 sel_0 sel_6 sel_2 sel_1
Xsky130_rom_krom_rom_column_mux_60 bl_3 bl_out_0 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_50 bl_13 bl_out_1 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_61 bl_2 bl_out_0 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_40 bl_23 bl_out_2 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_51 bl_12 bl_out_1 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_62 bl_1 bl_out_0 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_30 bl_33 bl_out_4 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_41 bl_22 bl_out_2 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_52 bl_11 bl_out_1 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_63 bl_0 bl_out_0 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_20 bl_43 bl_out_5 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_31 bl_32 bl_out_4 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_42 bl_21 bl_out_2 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_53 bl_10 bl_out_1 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_10 bl_53 bl_out_6 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_21 bl_42 bl_out_5 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_32 bl_31 bl_out_3 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_43 bl_20 bl_out_2 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_54 bl_9 bl_out_1 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_11 bl_52 bl_out_6 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_22 bl_41 bl_out_5 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_33 bl_30 bl_out_3 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_44 bl_19 bl_out_2 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_55 bl_8 bl_out_1 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_12 bl_51 bl_out_6 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_13 bl_50 bl_out_6 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_23 bl_40 bl_out_5 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_24 bl_39 bl_out_4 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_34 bl_29 bl_out_3 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_35 bl_28 bl_out_3 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_45 bl_18 bl_out_2 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_46 bl_17 bl_out_2 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_56 bl_7 bl_out_0 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_57 bl_6 bl_out_0 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_14 bl_49 bl_out_6 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_25 bl_38 bl_out_4 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_36 bl_27 bl_out_3 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_47 bl_16 bl_out_2 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_58 bl_5 bl_out_0 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_15 bl_48 bl_out_6 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_26 bl_37 bl_out_4 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_37 bl_26 bl_out_3 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_48 bl_15 bl_out_1 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_59 bl_4 bl_out_0 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_16 bl_47 bl_out_5 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_27 bl_36 bl_out_4 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_38 bl_25 bl_out_3 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_49 bl_14 bl_out_1 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_17 bl_46 bl_out_5 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_28 bl_35 bl_out_4 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_39 bl_24 bl_out_3 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_18 bl_45 bl_out_5 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_29 bl_34 bl_out_4 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_19 bl_44 bl_out_5 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_0 bl_63 bl_out_7 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_1 bl_62 bl_out_7 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_2 bl_61 bl_out_7 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_3 bl_60 bl_out_7 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_4 bl_59 bl_out_7 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_5 bl_58 bl_out_7 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_6 bl_57 bl_out_7 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_7 bl_56 bl_out_7 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_8 bl_55 bl_out_6 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_9 bl_54 bl_out_6 sel_6 gnd sky130_rom_krom_rom_column_mux
.ends

.subckt sky130_rom_krom_rom_precharge_array pre_bl0_out pre_bl3_out pre_bl5_out pre_bl6_out
+ pre_bl10_out pre_bl12_out pre_bl17_out pre_bl19_out pre_bl21_out pre_bl22_out pre_bl24_out
+ pre_bl26_out pre_bl28_out pre_bl29_out pre_bl30_out pre_bl31_out pre_bl35_out pre_bl37_out
+ pre_bl38_out pre_bl40_out pre_bl42_out pre_bl47_out pre_bl49_out pre_bl51_out pre_bl52_out
+ pre_bl53_out pre_bl56_out pre_bl58_out pre_bl59_out pre_bl60_out pre_bl61_out pre_bl62_out
+ gate pre_bl23_out pre_bl33_out pre_bl15_out pre_bl45_out pre_bl54_out pre_bl8_out
+ pre_bl1_out pre_bl63_out pre_bl36_out pre_bl4_out pre_bl34_out pre_bl27_out pre_bl20_out
+ pre_bl50_out pre_bl13_out pre_bl43_out pre_bl25_out pre_bl18_out pre_bl48_out pre_bl11_out
+ pre_bl57_out pre_bl41_out pre_bl16_out pre_bl46_out vdd pre_bl9_out pre_bl55_out
+ pre_bl39_out pre_bl2_out pre_bl32_out pre_bl14_out pre_bl44_out pre_bl7_out
Xsky130_rom_krom_precharge_cell_2 pre_bl61_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_3 pre_bl60_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_4 pre_bl59_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_5 pre_bl58_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_60 pre_bl3_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_6 pre_bl57_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_50 pre_bl13_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_61 pre_bl2_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_7 pre_bl56_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_8 pre_bl55_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_40 pre_bl23_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_51 pre_bl12_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_62 pre_bl1_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_9 pre_bl54_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_30 pre_bl33_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_41 pre_bl22_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_52 pre_bl11_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_63 pre_bl0_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_20 pre_bl43_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_31 pre_bl32_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_42 pre_bl21_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_53 pre_bl10_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_10 pre_bl53_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_11 pre_bl52_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_21 pre_bl42_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_22 pre_bl41_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_32 pre_bl31_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_33 pre_bl30_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_43 pre_bl20_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_44 pre_bl19_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_54 pre_bl9_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_55 pre_bl8_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_12 pre_bl51_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_23 pre_bl40_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_34 pre_bl29_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_45 pre_bl18_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_56 pre_bl7_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_13 pre_bl50_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_24 pre_bl39_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_35 pre_bl28_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_46 pre_bl17_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_57 pre_bl6_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_14 pre_bl49_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_25 pre_bl38_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_36 pre_bl27_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_47 pre_bl16_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_58 pre_bl5_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_15 pre_bl48_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_26 pre_bl37_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_37 pre_bl26_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_48 pre_bl15_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_59 pre_bl4_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_16 pre_bl47_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_27 pre_bl36_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_38 pre_bl25_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_49 pre_bl14_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_17 pre_bl46_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_28 pre_bl35_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_39 pre_bl24_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_18 pre_bl45_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_29 pre_bl34_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_19 pre_bl44_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_0 pre_bl63_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_1 pre_bl62_out gate vdd sky130_rom_krom_precharge_cell
.ends

.subckt sky130_rom_krom_rom_base_array bl_0_0 bl_0_1 bl_0_2 bl_0_3 bl_0_4 bl_0_5 bl_0_6
+ bl_0_7 bl_0_8 bl_0_9 bl_0_10 bl_0_11 bl_0_12 bl_0_13 bl_0_14 bl_0_15 bl_0_16 bl_0_17
+ bl_0_18 bl_0_19 bl_0_20 bl_0_21 bl_0_22 bl_0_23 bl_0_24 bl_0_25 bl_0_26 bl_0_27
+ bl_0_28 bl_0_29 bl_0_30 bl_0_31 bl_0_32 bl_0_33 bl_0_34 bl_0_35 bl_0_36 bl_0_37
+ bl_0_38 bl_0_39 bl_0_40 bl_0_41 bl_0_42 bl_0_43 bl_0_44 bl_0_45 bl_0_46 bl_0_47
+ bl_0_48 bl_0_49 bl_0_50 bl_0_51 bl_0_52 bl_0_53 bl_0_54 bl_0_55 bl_0_56 bl_0_57
+ bl_0_58 bl_0_59 bl_0_60 bl_0_61 bl_0_62 bl_0_63 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5
+ wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_12 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_26
+ wl_0_27 wl_0_28 wl_0_31 gnd_uq0 gnd wl_0_13 wl_0_22 wl_0_23 wl_0_14 wl_0_10 wl_0_24
+ wl_0_25 wl_0_20 wl_0_0 wl_0_21 precharge wl_0_29 wl_0_11 wl_0_30 vdd
Xsky130_rom_krom_rom_base_one_cell_910 wl_0_4 sky130_rom_krom_rom_base_one_cell_910/D
+ sky130_rom_krom_rom_base_one_cell_938/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_921 wl_0_4 sky130_rom_krom_rom_base_one_cell_921/D
+ sky130_rom_krom_rom_base_one_cell_921/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_932 wl_0_3 sky130_rom_krom_rom_base_one_cell_932/D
+ sky130_rom_krom_rom_base_one_cell_966/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_943 wl_0_3 sky130_rom_krom_rom_base_one_cell_943/D
+ sky130_rom_krom_rom_base_one_cell_971/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_954 wl_0_3 sky130_rom_krom_rom_base_one_cell_954/D
+ sky130_rom_krom_rom_base_one_cell_954/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_965 wl_0_2 sky130_rom_krom_rom_base_one_cell_965/D
+ sky130_rom_krom_rom_base_one_cell_999/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_976 wl_0_2 sky130_rom_krom_rom_base_one_cell_976/D
+ bl_0_25 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_987 wl_0_2 sky130_rom_krom_rom_base_one_cell_987/D
+ sky130_rom_krom_rom_base_one_cell_987/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_998 wl_0_1 sky130_rom_krom_rom_base_one_cell_998/D
+ bl_0_51 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_206 wl_0_27 sky130_rom_krom_rom_base_one_cell_72/S
+ sky130_rom_krom_rom_base_one_cell_267/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_217 wl_0_27 sky130_rom_krom_rom_base_one_cell_78/S
+ sky130_rom_krom_rom_base_one_cell_249/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_228 wl_0_27 sky130_rom_krom_rom_base_one_cell_228/D
+ sky130_rom_krom_rom_base_one_cell_288/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_239 wl_0_26 sky130_rom_krom_rom_base_one_cell_239/D
+ sky130_rom_krom_rom_base_one_cell_299/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_260 wl_0_23 sky130_rom_krom_rom_base_one_cell_376/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_271 wl_0_23 sky130_rom_krom_rom_base_one_cell_353/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_282 wl_0_23 sky130_rom_krom_rom_base_one_cell_420/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_293 wl_0_23 sky130_rom_krom_rom_base_one_cell_369/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1052 wl_0_0 sky130_rom_krom_rom_base_one_cell_1052/D
+ bl_0_12 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1041 wl_0_0 sky130_rom_krom_rom_base_one_cell_1041/D
+ bl_0_35 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1030 wl_0_0 sky130_rom_krom_rom_base_one_cell_990/S
+ bl_0_63 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_50 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_94/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_61 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_61/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_72 wl_0_31 sky130_rom_krom_rom_base_one_cell_72/D
+ sky130_rom_krom_rom_base_one_cell_72/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_83 wl_0_31 sky130_rom_krom_rom_base_one_cell_83/D
+ sky130_rom_krom_rom_base_one_cell_83/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_94 wl_0_31 sky130_rom_krom_rom_base_one_cell_94/D
+ sky130_rom_krom_rom_base_one_cell_94/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_740 wl_0_9 sky130_rom_krom_rom_base_one_cell_740/D
+ sky130_rom_krom_rom_base_one_cell_804/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_762 wl_0_9 sky130_rom_krom_rom_base_one_cell_762/D
+ sky130_rom_krom_rom_base_one_cell_900/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_795 wl_0_8 sky130_rom_krom_rom_base_one_cell_795/D
+ sky130_rom_krom_rom_base_one_cell_829/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_784 wl_0_8 sky130_rom_krom_rom_base_one_cell_784/D
+ sky130_rom_krom_rom_base_one_cell_819/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_751 wl_0_9 sky130_rom_krom_rom_base_one_cell_751/D
+ sky130_rom_krom_rom_base_one_cell_781/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_773 wl_0_8 sky130_rom_krom_rom_base_one_cell_773/D
+ sky130_rom_krom_rom_base_one_cell_838/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1051 wl_0_0 bl_0_5 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1040 wl_0_0 bl_0_23 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_581 wl_0_14 sky130_rom_krom_rom_base_one_cell_581/D
+ sky130_rom_krom_rom_base_one_cell_614/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_570 wl_0_15 sky130_rom_krom_rom_base_one_cell_570/D
+ sky130_rom_krom_rom_base_one_cell_597/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_592 wl_0_14 sky130_rom_krom_rom_base_one_cell_592/D
+ sky130_rom_krom_rom_base_one_cell_629/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_804 wl_0_7 sky130_rom_krom_rom_base_one_cell_905/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_859 wl_0_5 sky130_rom_krom_rom_base_one_cell_963/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_848 wl_0_6 sky130_rom_krom_rom_base_one_cell_979/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_837 wl_0_6 sky130_rom_krom_rom_base_one_cell_907/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_826 wl_0_7 sky130_rom_krom_rom_base_one_cell_864/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_815 wl_0_7 sky130_rom_krom_rom_base_one_cell_847/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_656 wl_0_12 sky130_rom_krom_rom_base_one_cell_685/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_645 wl_0_12 sky130_rom_krom_rom_base_one_cell_807/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_634 wl_0_13 sky130_rom_krom_rom_base_one_cell_702/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_601 wl_0_14 sky130_rom_krom_rom_base_one_cell_633/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_623 wl_0_13 sky130_rom_krom_rom_base_one_cell_658/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_612 wl_0_13 sky130_rom_krom_rom_base_one_cell_742/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_689 wl_0_11 sky130_rom_krom_rom_base_one_cell_718/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_678 wl_0_11 sky130_rom_krom_rom_base_one_cell_770/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_667 wl_0_12 sky130_rom_krom_rom_base_one_cell_700/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_497 wl_0_17 sky130_rom_krom_rom_base_one_cell_602/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_486 wl_0_17 sky130_rom_krom_rom_base_one_cell_541/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_475 wl_0_17 sky130_rom_krom_rom_base_one_cell_583/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_464 wl_0_18 sky130_rom_krom_rom_base_one_cell_603/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_453 wl_0_18 sky130_rom_krom_rom_base_one_cell_591/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_442 wl_0_18 sky130_rom_krom_rom_base_one_cell_583/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_431 wl_0_19 sky130_rom_krom_rom_base_one_cell_485/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_420 wl_0_19 sky130_rom_krom_rom_base_one_cell_477/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_900 wl_0_5 sky130_rom_krom_rom_base_one_cell_900/D
+ sky130_rom_krom_rom_base_one_cell_924/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_911 wl_0_4 sky130_rom_krom_rom_base_one_cell_911/D
+ sky130_rom_krom_rom_base_one_cell_939/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_922 wl_0_4 sky130_rom_krom_rom_base_one_cell_922/D
+ sky130_rom_krom_rom_base_one_cell_988/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_933 wl_0_3 sky130_rom_krom_rom_base_one_cell_933/D
+ sky130_rom_krom_rom_base_one_cell_933/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_944 wl_0_3 sky130_rom_krom_rom_base_one_cell_944/D
+ sky130_rom_krom_rom_base_one_cell_972/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_955 wl_0_3 sky130_rom_krom_rom_base_one_cell_955/D
+ sky130_rom_krom_rom_base_one_cell_955/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_966 wl_0_2 sky130_rom_krom_rom_base_one_cell_966/D
+ sky130_rom_krom_rom_base_one_cell_966/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_977 wl_0_2 sky130_rom_krom_rom_base_one_cell_977/D
+ sky130_rom_krom_rom_base_one_cell_977/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_988 wl_0_2 sky130_rom_krom_rom_base_one_cell_988/D
+ sky130_rom_krom_rom_base_one_cell_988/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_999 wl_0_1 sky130_rom_krom_rom_base_one_cell_999/D
+ sky130_rom_krom_rom_base_one_cell_999/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_207 wl_0_27 sky130_rom_krom_rom_base_zero_cell_65/S
+ sky130_rom_krom_rom_base_one_cell_269/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1053 wl_0_0 sky130_rom_krom_rom_base_one_cell_921/S
+ bl_0_8 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1042 wl_0_0 sky130_rom_krom_rom_base_one_cell_1042/D
+ bl_0_34 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1031 wl_0_0 sky130_rom_krom_rom_base_one_cell_992/S
+ bl_0_61 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1020 wl_0_1 sky130_rom_krom_rom_base_one_cell_985/S
+ bl_0_10 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_218 wl_0_27 sky130_rom_krom_rom_base_one_cell_79/S
+ sky130_rom_krom_rom_base_one_cell_277/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_229 wl_0_27 sky130_rom_krom_rom_base_one_cell_229/D
+ sky130_rom_krom_rom_base_one_cell_289/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_250 wl_0_24 sky130_rom_krom_rom_base_one_cell_398/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_261 wl_0_23 sky130_rom_krom_rom_base_one_cell_347/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_272 wl_0_23 sky130_rom_krom_rom_base_one_cell_412/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_283 wl_0_23 sky130_rom_krom_rom_base_one_cell_391/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_294 wl_0_23 sky130_rom_krom_rom_base_one_cell_370/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_40 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_85/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_51 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_95/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_62 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_62/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_73 wl_0_31 sky130_rom_krom_rom_base_one_cell_73/D
+ sky130_rom_krom_rom_base_one_cell_73/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_84 wl_0_31 sky130_rom_krom_rom_base_one_cell_84/D
+ sky130_rom_krom_rom_base_one_cell_84/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_95 wl_0_31 sky130_rom_krom_rom_base_one_cell_95/D
+ sky130_rom_krom_rom_base_one_cell_95/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_763 wl_0_9 sky130_rom_krom_rom_base_one_cell_763/D
+ sky130_rom_krom_rom_base_one_cell_798/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_752 wl_0_9 sky130_rom_krom_rom_base_one_cell_752/D
+ sky130_rom_krom_rom_base_one_cell_815/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_741 wl_0_9 sky130_rom_krom_rom_base_one_cell_741/D
+ sky130_rom_krom_rom_base_one_cell_806/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_730 wl_0_10 sky130_rom_krom_rom_base_one_cell_730/D
+ sky130_rom_krom_rom_base_one_cell_862/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_796 wl_0_8 sky130_rom_krom_rom_base_one_cell_796/D
+ sky130_rom_krom_rom_base_one_cell_830/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_785 wl_0_8 sky130_rom_krom_rom_base_one_cell_785/D
+ sky130_rom_krom_rom_base_one_cell_979/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_774 wl_0_8 sky130_rom_krom_rom_base_one_cell_774/D
+ sky130_rom_krom_rom_base_one_cell_809/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1030 wl_0_0 bl_0_40 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1052 wl_0_0 bl_0_4 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1041 wl_0_0 bl_0_22 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_593 wl_0_14 sky130_rom_krom_rom_base_one_cell_593/D
+ sky130_rom_krom_rom_base_one_cell_657/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_582 wl_0_14 sky130_rom_krom_rom_base_one_cell_582/D
+ sky130_rom_krom_rom_base_one_cell_771/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_571 wl_0_15 sky130_rom_krom_rom_base_one_cell_571/D
+ sky130_rom_krom_rom_base_one_cell_599/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_560 wl_0_15 sky130_rom_krom_rom_base_one_cell_560/D
+ sky130_rom_krom_rom_base_one_cell_589/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_838 wl_0_6 sky130_rom_krom_rom_base_one_cell_877/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_827 wl_0_7 sky130_rom_krom_rom_base_one_cell_865/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_816 wl_0_7 sky130_rom_krom_rom_base_one_cell_888/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_805 wl_0_7 sky130_rom_krom_rom_base_one_cell_907/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_390 wl_0_21 sky130_rom_krom_rom_base_one_cell_390/D
+ sky130_rom_krom_rom_base_one_cell_449/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_849 wl_0_6 sky130_rom_krom_rom_base_one_cell_948/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_679 wl_0_11 sky130_rom_krom_rom_base_one_cell_771/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_668 wl_0_12 sky130_rom_krom_rom_base_one_cell_702/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_657 wl_0_12 sky130_rom_krom_rom_base_one_cell_817/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_646 wl_0_12 sky130_rom_krom_rom_base_one_cell_742/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_635 wl_0_13 sky130_rom_krom_rom_base_one_cell_704/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_602 wl_0_14 sky130_rom_krom_rom_base_one_cell_634/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_624 wl_0_13 sky130_rom_krom_rom_base_one_cell_659/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_613 wl_0_13 sky130_rom_krom_rom_base_one_cell_713/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_498 wl_0_17 sky130_rom_krom_rom_base_one_cell_603/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_487 wl_0_17 sky130_rom_krom_rom_base_one_cell_630/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_476 wl_0_17 sky130_rom_krom_rom_base_one_cell_528/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_465 wl_0_18 sky130_rom_krom_rom_base_one_cell_604/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_454 wl_0_18 sky130_rom_krom_rom_base_one_cell_509/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_443 wl_0_18 sky130_rom_krom_rom_base_one_cell_530/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_432 wl_0_19 sky130_rom_krom_rom_base_one_cell_486/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_421 wl_0_19 sky130_rom_krom_rom_base_one_cell_478/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_410 wl_0_19 sky130_rom_krom_rom_base_one_cell_499/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_901 wl_0_4 sky130_rom_krom_rom_base_one_cell_901/D
+ sky130_rom_krom_rom_base_one_cell_926/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_912 wl_0_4 sky130_rom_krom_rom_base_one_cell_912/D
+ sky130_rom_krom_rom_base_one_cell_969/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_923 wl_0_4 sky130_rom_krom_rom_base_one_cell_923/D
+ sky130_rom_krom_rom_base_one_cell_955/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_934 wl_0_3 sky130_rom_krom_rom_base_one_cell_934/D
+ sky130_rom_krom_rom_base_one_cell_934/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_945 wl_0_3 sky130_rom_krom_rom_base_one_cell_945/D
+ sky130_rom_krom_rom_base_one_cell_973/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_956 wl_0_3 sky130_rom_krom_rom_base_one_cell_956/D
+ sky130_rom_krom_rom_base_one_cell_989/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_967 wl_0_2 sky130_rom_krom_rom_base_one_cell_967/D
+ bl_0_41 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_978 wl_0_2 sky130_rom_krom_rom_base_one_cell_978/D
+ sky130_rom_krom_rom_base_one_cell_978/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_989 wl_0_2 sky130_rom_krom_rom_base_one_cell_989/D
+ sky130_rom_krom_rom_base_one_cell_989/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_208 wl_0_27 sky130_rom_krom_rom_base_one_cell_208/D
+ sky130_rom_krom_rom_base_one_cell_301/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_219 wl_0_27 sky130_rom_krom_rom_base_zero_cell_76/S
+ sky130_rom_krom_rom_base_one_cell_252/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1010 wl_0_1 sky130_rom_krom_rom_base_one_cell_853/S
+ bl_0_26 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1054 wl_0_0 sky130_rom_krom_rom_base_one_cell_1054/D
+ bl_0_7 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1043 wl_0_0 sky130_rom_krom_rom_base_one_cell_942/S
+ bl_0_33 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1032 wl_0_0 sky130_rom_krom_rom_base_one_cell_993/S
+ bl_0_60 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1021 wl_0_1 sky130_rom_krom_rom_base_one_cell_986/S
+ bl_0_9 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_240 wl_0_24 sky130_rom_krom_rom_base_one_cell_420/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_251 wl_0_24 sky130_rom_krom_rom_base_one_cell_342/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_262 wl_0_23 sky130_rom_krom_rom_base_one_cell_377/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_273 wl_0_23 sky130_rom_krom_rom_base_one_cell_443/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_284 wl_0_23 sky130_rom_krom_rom_base_one_cell_423/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_295 wl_0_22 sky130_rom_krom_rom_base_one_cell_372/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_30 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_77/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_41 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_86/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_52 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_96/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_63 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_63/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_74 wl_0_31 sky130_rom_krom_rom_base_one_cell_74/D
+ sky130_rom_krom_rom_base_one_cell_74/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_85 wl_0_31 sky130_rom_krom_rom_base_one_cell_85/D
+ sky130_rom_krom_rom_base_one_cell_85/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_96 wl_0_31 sky130_rom_krom_rom_base_one_cell_96/D
+ sky130_rom_krom_rom_base_one_cell_96/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_797 wl_0_8 sky130_rom_krom_rom_base_one_cell_797/D
+ sky130_rom_krom_rom_base_one_cell_831/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_786 wl_0_8 sky130_rom_krom_rom_base_one_cell_786/D
+ sky130_rom_krom_rom_base_one_cell_948/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_753 wl_0_9 sky130_rom_krom_rom_base_one_cell_753/D
+ sky130_rom_krom_rom_base_one_cell_853/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_775 wl_0_8 sky130_rom_krom_rom_base_one_cell_775/D
+ sky130_rom_krom_rom_base_one_cell_878/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_742 wl_0_9 sky130_rom_krom_rom_base_one_cell_742/D
+ sky130_rom_krom_rom_base_one_cell_808/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_764 wl_0_8 sky130_rom_krom_rom_base_one_cell_764/D
+ sky130_rom_krom_rom_base_one_cell_800/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_731 wl_0_10 sky130_rom_krom_rom_base_one_cell_731/D
+ sky130_rom_krom_rom_base_one_cell_790/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_720 wl_0_10 sky130_rom_krom_rom_base_one_cell_720/D
+ sky130_rom_krom_rom_base_one_cell_751/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1053 wl_0_0 bl_0_2 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1042 wl_0_0 bl_0_19 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1031 wl_0_0 bl_0_39 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1020 wl_0_0 bl_0_57 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_594 wl_0_14 sky130_rom_krom_rom_base_one_cell_594/D
+ sky130_rom_krom_rom_base_one_cell_662/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_583 wl_0_14 sky130_rom_krom_rom_base_one_cell_583/D
+ sky130_rom_krom_rom_base_one_cell_647/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_572 wl_0_15 sky130_rom_krom_rom_base_one_cell_572/D
+ sky130_rom_krom_rom_base_one_cell_668/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_561 wl_0_15 sky130_rom_krom_rom_base_one_cell_561/D
+ sky130_rom_krom_rom_base_one_cell_623/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_550 wl_0_15 sky130_rom_krom_rom_base_one_cell_550/D
+ sky130_rom_krom_rom_base_one_cell_576/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_839 wl_0_6 sky130_rom_krom_rom_base_one_cell_908/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_828 wl_0_7 sky130_rom_krom_rom_base_one_cell_866/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_817 wl_0_7 sky130_rom_krom_rom_base_one_cell_852/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_806 wl_0_7 sky130_rom_krom_rom_base_one_cell_838/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_380 wl_0_21 sky130_rom_krom_rom_base_one_cell_380/D
+ sky130_rom_krom_rom_base_one_cell_408/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_391 wl_0_21 sky130_rom_krom_rom_base_one_cell_391/D
+ sky130_rom_krom_rom_base_one_cell_421/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_669 wl_0_12 sky130_rom_krom_rom_base_one_cell_703/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_658 wl_0_12 sky130_rom_krom_rom_base_one_cell_687/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_647 wl_0_12 sky130_rom_krom_rom_base_one_cell_713/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_636 wl_0_13 sky130_rom_krom_rom_base_one_cell_705/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_603 wl_0_14 sky130_rom_krom_rom_base_one_cell_636/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_625 wl_0_13 sky130_rom_krom_rom_base_one_cell_661/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_614 wl_0_13 sky130_rom_krom_rom_base_one_cell_677/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_411 wl_0_19 sky130_rom_krom_rom_base_one_cell_500/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_400 wl_0_19 sky130_rom_krom_rom_base_one_cell_522/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_499 wl_0_17 sky130_rom_krom_rom_base_one_cell_604/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_488 wl_0_17 sky130_rom_krom_rom_base_one_cell_542/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_477 wl_0_17 sky130_rom_krom_rom_base_one_cell_529/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_466 wl_0_18 sky130_rom_krom_rom_base_one_cell_520/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_455 wl_0_18 sky130_rom_krom_rom_base_one_cell_541/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_444 wl_0_18 sky130_rom_krom_rom_base_one_cell_558/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_433 wl_0_19 sky130_rom_krom_rom_base_one_cell_488/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_422 wl_0_19 sky130_rom_krom_rom_base_one_cell_541/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_902 wl_0_4 sky130_rom_krom_rom_base_one_cell_902/D
+ sky130_rom_krom_rom_base_one_cell_959/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_913 wl_0_4 sky130_rom_krom_rom_base_one_cell_913/D
+ sky130_rom_krom_rom_base_one_cell_913/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_924 wl_0_4 sky130_rom_krom_rom_base_one_cell_924/D
+ sky130_rom_krom_rom_base_one_cell_956/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_935 wl_0_3 sky130_rom_krom_rom_base_one_cell_935/D
+ sky130_rom_krom_rom_base_one_cell_935/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_946 wl_0_3 sky130_rom_krom_rom_base_one_cell_946/D
+ sky130_rom_krom_rom_base_one_cell_976/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_957 wl_0_3 sky130_rom_krom_rom_base_one_cell_957/D
+ sky130_rom_krom_rom_base_one_cell_957/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_968 wl_0_2 sky130_rom_krom_rom_base_one_cell_968/D
+ sky130_rom_krom_rom_base_one_cell_968/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_979 wl_0_2 sky130_rom_krom_rom_base_one_cell_979/D
+ sky130_rom_krom_rom_base_one_cell_979/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_209 wl_0_27 sky130_rom_krom_rom_base_one_cell_209/D
+ sky130_rom_krom_rom_base_one_cell_271/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_230 wl_0_24 sky130_rom_krom_rom_base_one_cell_327/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_241 wl_0_24 sky130_rom_krom_rom_base_one_cell_391/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_252 wl_0_24 sky130_rom_krom_rom_base_one_cell_367/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_263 wl_0_23 sky130_rom_krom_rom_base_one_cell_348/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1000 wl_0_1 sky130_rom_krom_rom_base_one_cell_934/S
+ bl_0_47 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1011 wl_0_1 sky130_rom_krom_rom_base_one_cell_977/S
+ bl_0_24 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1055 wl_0_0 sky130_rom_krom_rom_base_one_cell_1055/D
+ bl_0_3 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1044 wl_0_0 sky130_rom_krom_rom_base_one_cell_971/S
+ bl_0_31 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1033 wl_0_0 sky130_rom_krom_rom_base_one_cell_995/S
+ bl_0_58 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1022 wl_0_1 sky130_rom_krom_rom_base_one_cell_987/S
+ sky130_rom_krom_rom_base_one_cell_1054/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_20 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_74/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_31 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_78/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_274 wl_0_23 sky130_rom_krom_rom_base_one_cell_414/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_285 wl_0_23 sky130_rom_krom_rom_base_one_cell_392/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_296 wl_0_22 sky130_rom_krom_rom_base_one_cell_373/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_42 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_87/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_53 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_53/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_64 wl_0_31 sky130_rom_krom_rom_base_one_cell_2/S
+ sky130_rom_krom_rom_base_one_cell_64/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_75 wl_0_31 sky130_rom_krom_rom_base_one_cell_75/D
+ sky130_rom_krom_rom_base_one_cell_75/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_86 wl_0_31 sky130_rom_krom_rom_base_one_cell_86/D
+ sky130_rom_krom_rom_base_one_cell_86/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_97 wl_0_31 sky130_rom_krom_rom_base_one_cell_97/D
+ sky130_rom_krom_rom_base_one_cell_97/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_798 wl_0_8 sky130_rom_krom_rom_base_one_cell_798/D
+ sky130_rom_krom_rom_base_one_cell_832/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_787 wl_0_8 sky130_rom_krom_rom_base_one_cell_787/D
+ sky130_rom_krom_rom_base_one_cell_919/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_754 wl_0_9 sky130_rom_krom_rom_base_one_cell_754/D
+ sky130_rom_krom_rom_base_one_cell_822/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_776 wl_0_8 sky130_rom_krom_rom_base_one_cell_776/D
+ sky130_rom_krom_rom_base_one_cell_841/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_743 wl_0_9 sky130_rom_krom_rom_base_one_cell_743/D
+ sky130_rom_krom_rom_base_one_cell_774/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_765 wl_0_8 sky130_rom_krom_rom_base_one_cell_765/D
+ sky130_rom_krom_rom_base_one_cell_802/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_732 wl_0_10 sky130_rom_krom_rom_base_one_cell_732/D
+ sky130_rom_krom_rom_base_one_cell_757/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_721 wl_0_10 sky130_rom_krom_rom_base_one_cell_721/D
+ sky130_rom_krom_rom_base_one_cell_782/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_710 wl_0_10 sky130_rom_krom_rom_base_one_cell_710/D
+ sky130_rom_krom_rom_base_one_cell_772/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1010 wl_0_1 sky130_rom_krom_rom_base_one_cell_975/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1054 wl_0_0 bl_0_0 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1043 wl_0_0 bl_0_17 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1032 wl_0_0 bl_0_38 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1021 wl_0_0 bl_0_56 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_595 wl_0_14 sky130_rom_krom_rom_base_one_cell_595/D
+ sky130_rom_krom_rom_base_one_cell_726/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_584 wl_0_14 sky130_rom_krom_rom_base_one_cell_584/D
+ sky130_rom_krom_rom_base_one_cell_617/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_573 wl_0_15 sky130_rom_krom_rom_base_one_cell_573/D
+ sky130_rom_krom_rom_base_one_cell_600/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_562 wl_0_15 sky130_rom_krom_rom_base_one_cell_562/D
+ sky130_rom_krom_rom_base_one_cell_624/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_551 wl_0_15 sky130_rom_krom_rom_base_one_cell_551/D
+ sky130_rom_krom_rom_base_one_cell_577/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_540 wl_0_16 sky130_rom_krom_rom_base_one_cell_540/D
+ sky130_rom_krom_rom_base_one_cell_628/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_370 wl_0_22 sky130_rom_krom_rom_base_one_cell_370/D
+ sky130_rom_krom_rom_base_one_cell_431/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_381 wl_0_21 sky130_rom_krom_rom_base_one_cell_381/D
+ sky130_rom_krom_rom_base_one_cell_409/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_829 wl_0_7 sky130_rom_krom_rom_base_one_cell_900/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_818 wl_0_7 sky130_rom_krom_rom_base_one_cell_853/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_807 wl_0_7 sky130_rom_krom_rom_base_one_cell_878/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_392 wl_0_21 sky130_rom_krom_rom_base_one_cell_392/D
+ sky130_rom_krom_rom_base_one_cell_426/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_604 wl_0_14 sky130_rom_krom_rom_base_one_cell_637/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_659 wl_0_12 sky130_rom_krom_rom_base_one_cell_754/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_648 wl_0_12 sky130_rom_krom_rom_base_one_cell_676/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_637 wl_0_12 sky130_rom_krom_rom_base_one_cell_737/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_626 wl_0_13 sky130_rom_krom_rom_base_one_cell_662/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_615 wl_0_13 sky130_rom_krom_rom_base_one_cell_651/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_445 wl_0_18 sky130_rom_krom_rom_base_one_cell_497/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_434 wl_0_19 sky130_rom_krom_rom_base_one_cell_602/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_423 wl_0_19 sky130_rom_krom_rom_base_one_cell_630/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_412 wl_0_19 sky130_rom_krom_rom_base_one_cell_470/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_401 wl_0_19 sky130_rom_krom_rom_base_one_cell_492/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_489 wl_0_17 sky130_rom_krom_rom_base_one_cell_543/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_478 wl_0_17 sky130_rom_krom_rom_base_one_cell_530/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_467 wl_0_18 sky130_rom_krom_rom_base_one_cell_704/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_456 wl_0_18 sky130_rom_krom_rom_base_one_cell_630/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_903 wl_0_4 sky130_rom_krom_rom_base_one_cell_903/D
+ sky130_rom_krom_rom_base_one_cell_960/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_914 wl_0_4 sky130_rom_krom_rom_base_one_cell_914/D
+ sky130_rom_krom_rom_base_one_cell_970/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_925 wl_0_4 sky130_rom_krom_rom_base_one_cell_925/D
+ sky130_rom_krom_rom_base_one_cell_957/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_936 wl_0_3 sky130_rom_krom_rom_base_one_cell_936/D
+ sky130_rom_krom_rom_base_one_cell_936/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_947 wl_0_3 sky130_rom_krom_rom_base_one_cell_947/D
+ sky130_rom_krom_rom_base_one_cell_977/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_958 wl_0_2 sky130_rom_krom_rom_base_one_cell_958/D
+ sky130_rom_krom_rom_base_one_cell_990/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_969 wl_0_2 sky130_rom_krom_rom_base_one_cell_969/D
+ sky130_rom_krom_rom_base_one_cell_969/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_990 wl_0_2 sky130_rom_krom_rom_base_one_cell_954/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1001 wl_0_1 sky130_rom_krom_rom_base_one_cell_936/S
+ sky130_rom_krom_rom_base_one_cell_1039/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_220 wl_0_24 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_231 wl_0_24 sky130_rom_krom_rom_base_one_cell_328/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_242 wl_0_24 sky130_rom_krom_rom_base_one_cell_337/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_253 wl_0_24 sky130_rom_krom_rom_base_one_cell_368/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_264 wl_0_23 sky130_rom_krom_rom_base_one_cell_349/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_275 wl_0_23 sky130_rom_krom_rom_base_one_cell_355/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_286 wl_0_23 sky130_rom_krom_rom_base_one_cell_364/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_297 wl_0_22 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1012 wl_0_1 sky130_rom_krom_rom_base_one_cell_978/S
+ bl_0_23 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1056 wl_0_0 sky130_rom_krom_rom_base_one_cell_1056/D
+ bl_0_1 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1045 wl_0_0 sky130_rom_krom_rom_base_one_cell_1045/D
+ bl_0_29 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1034 wl_0_0 sky130_rom_krom_rom_base_one_cell_906/S
+ bl_0_53 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1023 wl_0_1 sky130_rom_krom_rom_base_one_cell_867/S
+ bl_0_6 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_10 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_5/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_21 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_21/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_32 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_79/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_43 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_43/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_54 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_97/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_65 wl_0_31 sky130_rom_krom_rom_base_one_cell_4/S
+ sky130_rom_krom_rom_base_one_cell_65/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_76 wl_0_31 sky130_rom_krom_rom_base_one_cell_76/D
+ sky130_rom_krom_rom_base_one_cell_76/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_87 wl_0_31 sky130_rom_krom_rom_base_one_cell_87/D
+ sky130_rom_krom_rom_base_one_cell_87/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_98 wl_0_31 sky130_rom_krom_rom_base_one_cell_98/D
+ sky130_rom_krom_rom_base_one_cell_98/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_700 wl_0_11 sky130_rom_krom_rom_base_one_cell_700/D
+ sky130_rom_krom_rom_base_one_cell_734/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_711 wl_0_10 sky130_rom_krom_rom_base_one_cell_711/D
+ sky130_rom_krom_rom_base_one_cell_741/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_799 wl_0_8 sky130_rom_krom_rom_base_one_cell_799/D
+ sky130_rom_krom_rom_base_one_cell_833/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_788 wl_0_8 sky130_rom_krom_rom_base_one_cell_788/D
+ sky130_rom_krom_rom_base_one_cell_860/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_755 wl_0_9 sky130_rom_krom_rom_base_one_cell_755/D
+ sky130_rom_krom_rom_base_one_cell_786/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_777 wl_0_8 sky130_rom_krom_rom_base_one_cell_777/D
+ sky130_rom_krom_rom_base_one_cell_880/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_744 wl_0_9 sky130_rom_krom_rom_base_one_cell_744/D
+ sky130_rom_krom_rom_base_one_cell_776/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_766 wl_0_8 sky130_rom_krom_rom_base_one_cell_766/D
+ sky130_rom_krom_rom_base_one_cell_803/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_733 wl_0_10 sky130_rom_krom_rom_base_one_cell_733/D
+ sky130_rom_krom_rom_base_one_cell_758/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_722 wl_0_10 sky130_rom_krom_rom_base_one_cell_722/D
+ sky130_rom_krom_rom_base_one_cell_752/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1000 wl_0_1 sky130_rom_krom_rom_base_one_cell_935/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1011 wl_0_1 bl_0_25 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1044 wl_0_0 bl_0_16 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1033 wl_0_0 bl_0_37 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1022 wl_0_0 bl_0_55 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_563 wl_0_15 sky130_rom_krom_rom_base_one_cell_563/D
+ sky130_rom_krom_rom_base_one_cell_654/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_552 wl_0_15 sky130_rom_krom_rom_base_one_cell_552/D
+ sky130_rom_krom_rom_base_one_cell_579/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_541 wl_0_16 sky130_rom_krom_rom_base_one_cell_541/D
+ sky130_rom_krom_rom_base_one_cell_659/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_530 wl_0_16 sky130_rom_krom_rom_base_one_cell_530/D
+ sky130_rom_krom_rom_base_one_cell_557/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_596 wl_0_14 sky130_rom_krom_rom_base_one_cell_596/D
+ sky130_rom_krom_rom_base_one_cell_664/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_585 wl_0_14 sky130_rom_krom_rom_base_one_cell_585/D
+ sky130_rom_krom_rom_base_one_cell_742/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_574 wl_0_15 sky130_rom_krom_rom_base_one_cell_574/D
+ sky130_rom_krom_rom_base_one_cell_606/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_360 wl_0_22 sky130_rom_krom_rom_base_one_cell_360/D
+ sky130_rom_krom_rom_base_one_cell_418/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_371 wl_0_22 sky130_rom_krom_rom_base_one_cell_371/D
+ sky130_rom_krom_rom_base_one_cell_401/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_382 wl_0_21 sky130_rom_krom_rom_base_one_cell_382/D
+ sky130_rom_krom_rom_base_one_cell_587/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_393 wl_0_21 sky130_rom_krom_rom_base_one_cell_393/D
+ sky130_rom_krom_rom_base_one_cell_451/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_819 wl_0_7 sky130_rom_krom_rom_base_one_cell_979/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_808 wl_0_7 sky130_rom_krom_rom_base_one_cell_841/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_605 wl_0_14 sky130_rom_krom_rom_base_one_cell_668/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_627 wl_0_13 sky130_rom_krom_rom_base_one_cell_726/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_616 wl_0_13 sky130_rom_krom_rom_base_one_cell_678/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_190 wl_0_28 sky130_rom_krom_rom_base_one_cell_95/S
+ sky130_rom_krom_rom_base_one_cell_227/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_649 wl_0_12 sky130_rom_krom_rom_base_one_cell_677/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_638 wl_0_12 sky130_rom_krom_rom_base_one_cell_765/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_479 wl_0_17 sky130_rom_krom_rom_base_one_cell_558/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_468 wl_0_18 sky130_rom_krom_rom_base_one_cell_548/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_457 wl_0_18 sky130_rom_krom_rom_base_one_cell_543/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_446 wl_0_18 sky130_rom_krom_rom_base_one_cell_587/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_435 wl_0_19 sky130_rom_krom_rom_base_one_cell_603/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_424 wl_0_19 sky130_rom_krom_rom_base_one_cell_479/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_413 wl_0_19 sky130_rom_krom_rom_base_one_cell_471/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_402 wl_0_19 sky130_rom_krom_rom_base_one_cell_523/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_904 wl_0_4 sky130_rom_krom_rom_base_one_cell_904/D
+ sky130_rom_krom_rom_base_one_cell_928/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_915 wl_0_4 sky130_rom_krom_rom_base_one_cell_915/D
+ sky130_rom_krom_rom_base_one_cell_944/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_926 wl_0_3 sky130_rom_krom_rom_base_one_cell_926/D
+ sky130_rom_krom_rom_base_one_cell_958/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_937 wl_0_3 sky130_rom_krom_rom_base_one_cell_937/D
+ sky130_rom_krom_rom_base_one_cell_937/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_948 wl_0_3 sky130_rom_krom_rom_base_one_cell_948/D
+ sky130_rom_krom_rom_base_one_cell_948/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_959 wl_0_2 sky130_rom_krom_rom_base_one_cell_959/D
+ sky130_rom_krom_rom_base_one_cell_991/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_980 wl_0_2 sky130_rom_krom_rom_base_one_cell_942/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_991 wl_0_2 sky130_rom_krom_rom_base_one_cell_955/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1002 wl_0_1 sky130_rom_krom_rom_base_one_cell_937/S
+ bl_0_43 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1035 wl_0_0 sky130_rom_krom_rom_base_one_cell_999/S
+ bl_0_50 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1024 wl_0_1 sky130_rom_krom_rom_base_one_cell_988/S
+ bl_0_5 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1013 wl_0_1 sky130_rom_krom_rom_base_one_cell_979/S
+ sky130_rom_krom_rom_base_one_cell_1048/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_221 wl_0_24 sky130_rom_krom_rom_base_one_cell_320/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_232 wl_0_24 sky130_rom_krom_rom_base_one_cell_355/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_243 wl_0_24 sky130_rom_krom_rom_base_one_cell_338/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_210 wl_0_25 sky130_rom_krom_rom_base_one_cell_340/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_254 wl_0_24 sky130_rom_krom_rom_base_one_cell_343/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_265 wl_0_23 sky130_rom_krom_rom_base_one_cell_438/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_276 wl_0_23 sky130_rom_krom_rom_base_one_cell_356/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_287 wl_0_23 sky130_rom_krom_rom_base_one_cell_395/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_298 wl_0_22 sky130_rom_krom_rom_base_one_cell_375/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1046 wl_0_0 sky130_rom_krom_rom_base_one_cell_974/S
+ bl_0_28 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_11 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_69/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_22 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_22/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_33 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_80/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_44 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_88/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_55 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_55/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_66 wl_0_31 sky130_rom_krom_rom_base_one_cell_5/S
+ sky130_rom_krom_rom_base_one_cell_66/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_77 wl_0_31 sky130_rom_krom_rom_base_one_cell_77/D
+ sky130_rom_krom_rom_base_one_cell_77/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_88 wl_0_31 sky130_rom_krom_rom_base_one_cell_88/D
+ sky130_rom_krom_rom_base_one_cell_88/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_99 wl_0_31 sky130_rom_krom_rom_base_one_cell_99/D
+ sky130_rom_krom_rom_base_one_cell_99/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_745 wl_0_9 sky130_rom_krom_rom_base_one_cell_745/D
+ sky130_rom_krom_rom_base_one_cell_777/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_701 wl_0_11 sky130_rom_krom_rom_base_one_cell_701/D
+ sky130_rom_krom_rom_base_one_cell_735/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_734 wl_0_10 sky130_rom_krom_rom_base_one_cell_734/D
+ sky130_rom_krom_rom_base_one_cell_759/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_723 wl_0_10 sky130_rom_krom_rom_base_one_cell_723/D
+ sky130_rom_krom_rom_base_one_cell_783/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_712 wl_0_10 sky130_rom_krom_rom_base_one_cell_712/D
+ sky130_rom_krom_rom_base_one_cell_775/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_756 wl_0_9 sky130_rom_krom_rom_base_one_cell_756/D
+ sky130_rom_krom_rom_base_one_cell_824/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_789 wl_0_8 sky130_rom_krom_rom_base_one_cell_789/D
+ sky130_rom_krom_rom_base_one_cell_825/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_778 wl_0_8 sky130_rom_krom_rom_base_one_cell_778/D
+ sky130_rom_krom_rom_base_one_cell_883/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_767 wl_0_8 sky130_rom_krom_rom_base_one_cell_767/D
+ sky130_rom_krom_rom_base_one_cell_835/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1001 wl_0_1 bl_0_44 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1012 wl_0_1 bl_0_22 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1045 wl_0_0 bl_0_15 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1034 wl_0_0 bl_0_36 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1023 wl_0_0 bl_0_54 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_597 wl_0_14 sky130_rom_krom_rom_base_one_cell_597/D
+ sky130_rom_krom_rom_base_one_cell_635/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_586 wl_0_14 sky130_rom_krom_rom_base_one_cell_586/D
+ sky130_rom_krom_rom_base_one_cell_619/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_575 wl_0_14 sky130_rom_krom_rom_base_one_cell_575/D
+ sky130_rom_krom_rom_base_one_cell_608/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_564 wl_0_15 sky130_rom_krom_rom_base_one_cell_564/D
+ sky130_rom_krom_rom_base_one_cell_592/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_553 wl_0_15 sky130_rom_krom_rom_base_one_cell_553/D
+ sky130_rom_krom_rom_base_one_cell_580/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_542 wl_0_16 sky130_rom_krom_rom_base_one_cell_542/D
+ sky130_rom_krom_rom_base_one_cell_566/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_531 wl_0_16 sky130_rom_krom_rom_base_one_cell_531/D
+ sky130_rom_krom_rom_base_one_cell_559/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_520 wl_0_17 sky130_rom_krom_rom_base_one_cell_520/D
+ sky130_rom_krom_rom_base_one_cell_547/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_809 wl_0_7 sky130_rom_krom_rom_base_one_cell_880/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_350 wl_0_22 sky130_rom_krom_rom_base_one_cell_350/D
+ sky130_rom_krom_rom_base_one_cell_380/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_361 wl_0_22 sky130_rom_krom_rom_base_one_cell_361/D
+ sky130_rom_krom_rom_base_one_cell_630/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_372 wl_0_21 sky130_rom_krom_rom_base_one_cell_372/D
+ sky130_rom_krom_rom_base_one_cell_402/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_383 wl_0_21 sky130_rom_krom_rom_base_one_cell_383/D
+ sky130_rom_krom_rom_base_one_cell_468/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_394 wl_0_21 sky130_rom_krom_rom_base_one_cell_394/D
+ sky130_rom_krom_rom_base_one_cell_485/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_639 wl_0_12 sky130_rom_krom_rom_base_one_cell_706/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_606 wl_0_14 sky130_rom_krom_rom_base_one_cell_639/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_628 wl_0_13 sky130_rom_krom_rom_base_one_cell_664/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_617 wl_0_13 sky130_rom_krom_rom_base_one_cell_652/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_180 wl_0_28 sky130_rom_krom_rom_base_one_cell_35/S
+ sky130_rom_krom_rom_base_one_cell_280/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_191 wl_0_28 sky130_rom_krom_rom_base_zero_cell_88/S
+ sky130_rom_krom_rom_base_one_cell_228/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_469 wl_0_18 sky130_rom_krom_rom_base_one_cell_607/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_458 wl_0_18 sky130_rom_krom_rom_base_one_cell_513/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_447 wl_0_18 sky130_rom_krom_rom_base_one_cell_499/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_436 wl_0_19 sky130_rom_krom_rom_base_one_cell_520/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_425 wl_0_19 sky130_rom_krom_rom_base_one_cell_481/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_414 wl_0_19 sky130_rom_krom_rom_base_one_cell_473/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_403 wl_0_19 sky130_rom_krom_rom_base_one_cell_524/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_905 wl_0_4 sky130_rom_krom_rom_base_one_cell_905/D
+ sky130_rom_krom_rom_base_one_cell_929/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_916 wl_0_4 sky130_rom_krom_rom_base_one_cell_916/D
+ sky130_rom_krom_rom_base_one_cell_974/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_927 wl_0_3 sky130_rom_krom_rom_base_one_cell_927/D
+ sky130_rom_krom_rom_base_one_cell_961/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_938 wl_0_3 sky130_rom_krom_rom_base_one_cell_938/D
+ sky130_rom_krom_rom_base_one_cell_967/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_949 wl_0_3 sky130_rom_krom_rom_base_one_cell_949/D
+ bl_0_19 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_970 wl_0_2 sky130_rom_krom_rom_base_one_cell_935/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_981 wl_0_2 sky130_rom_krom_rom_base_one_cell_853/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_992 wl_0_2 sky130_rom_krom_rom_base_one_cell_870/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_200 wl_0_25 sky130_rom_krom_rom_base_one_cell_307/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_211 wl_0_25 sky130_rom_krom_rom_base_one_cell_364/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1003 wl_0_1 sky130_rom_krom_rom_base_one_cell_883/S
+ bl_0_40 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1047 wl_0_0 sky130_rom_krom_rom_base_one_cell_975/S
+ bl_0_27 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1036 wl_0_0 sky130_rom_krom_rom_base_one_cell_966/S
+ bl_0_49 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1025 wl_0_1 sky130_rom_krom_rom_base_one_cell_954/S
+ bl_0_4 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1014 wl_0_1 sky130_rom_krom_rom_base_one_cell_948/S
+ sky130_rom_krom_rom_base_one_cell_1049/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_222 wl_0_24 sky130_rom_krom_rom_base_one_cell_376/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_233 wl_0_24 sky130_rom_krom_rom_base_one_cell_356/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_244 wl_0_24 sky130_rom_krom_rom_base_one_cell_339/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_255 wl_0_24 sky130_rom_krom_rom_base_one_cell_344/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_266 wl_0_23 sky130_rom_krom_rom_base_one_cell_379/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_277 wl_0_23 sky130_rom_krom_rom_base_one_cell_507/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_288 wl_0_23 sky130_rom_krom_rom_base_one_cell_365/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_299 wl_0_22 sky130_rom_krom_rom_base_one_cell_376/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_12 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_70/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_23 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_75/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_34 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_81/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_45 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_89/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_56 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_98/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_67 wl_0_31 sky130_rom_krom_rom_base_one_cell_6/S
+ sky130_rom_krom_rom_base_one_cell_67/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_78 wl_0_31 sky130_rom_krom_rom_base_one_cell_78/D
+ sky130_rom_krom_rom_base_one_cell_78/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_89 wl_0_31 sky130_rom_krom_rom_base_one_cell_89/D
+ sky130_rom_krom_rom_base_one_cell_89/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_757 wl_0_9 sky130_rom_krom_rom_base_one_cell_757/D
+ sky130_rom_krom_rom_base_one_cell_791/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_779 wl_0_8 sky130_rom_krom_rom_base_one_cell_779/D
+ sky130_rom_krom_rom_base_one_cell_813/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_746 wl_0_9 sky130_rom_krom_rom_base_one_cell_746/D
+ sky130_rom_krom_rom_base_one_cell_810/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_768 wl_0_8 sky130_rom_krom_rom_base_one_cell_768/D
+ sky130_rom_krom_rom_base_one_cell_875/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_702 wl_0_11 sky130_rom_krom_rom_base_one_cell_702/D
+ sky130_rom_krom_rom_base_one_cell_795/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_735 wl_0_10 sky130_rom_krom_rom_base_one_cell_735/D
+ sky130_rom_krom_rom_base_one_cell_760/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_724 wl_0_10 sky130_rom_krom_rom_base_one_cell_724/D
+ sky130_rom_krom_rom_base_one_cell_821/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_713 wl_0_10 sky130_rom_krom_rom_base_one_cell_713/D
+ sky130_rom_krom_rom_base_one_cell_744/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1002 wl_0_1 sky130_rom_krom_rom_base_one_cell_882/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1046 wl_0_0 bl_0_13 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1035 wl_0_0 bl_0_32 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1024 wl_0_0 bl_0_52 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1013 wl_0_1 bl_0_19 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_598 wl_0_14 sky130_rom_krom_rom_base_one_cell_598/D
+ sky130_rom_krom_rom_base_one_cell_697/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_587 wl_0_14 sky130_rom_krom_rom_base_one_cell_587/D
+ sky130_rom_krom_rom_base_one_cell_713/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_576 wl_0_14 sky130_rom_krom_rom_base_one_cell_576/D
+ sky130_rom_krom_rom_base_one_cell_609/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_565 wl_0_15 sky130_rom_krom_rom_base_one_cell_565/D
+ sky130_rom_krom_rom_base_one_cell_593/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_554 wl_0_15 sky130_rom_krom_rom_base_one_cell_554/D
+ sky130_rom_krom_rom_base_one_cell_581/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_543 wl_0_16 sky130_rom_krom_rom_base_one_cell_543/D
+ sky130_rom_krom_rom_base_one_cell_567/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_532 wl_0_16 sky130_rom_krom_rom_base_one_cell_532/D
+ sky130_rom_krom_rom_base_one_cell_677/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_521 wl_0_16 sky130_rom_krom_rom_base_one_cell_521/D
+ sky130_rom_krom_rom_base_one_cell_550/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_510 wl_0_17 sky130_rom_krom_rom_base_one_cell_510/D
+ sky130_rom_krom_rom_base_one_cell_564/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_0 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_0/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_340 wl_0_23 sky130_rom_krom_rom_base_one_cell_340/D
+ sky130_rom_krom_rom_base_one_cell_393/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_351 wl_0_22 sky130_rom_krom_rom_base_one_cell_351/D
+ sky130_rom_krom_rom_base_one_cell_440/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_362 wl_0_22 sky130_rom_krom_rom_base_one_cell_362/D
+ sky130_rom_krom_rom_base_one_cell_389/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_373 wl_0_21 sky130_rom_krom_rom_base_one_cell_373/D
+ sky130_rom_krom_rom_base_one_cell_491/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_384 wl_0_21 sky130_rom_krom_rom_base_one_cell_384/D
+ sky130_rom_krom_rom_base_one_cell_413/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_395 wl_0_21 sky130_rom_krom_rom_base_one_cell_395/D
+ sky130_rom_krom_rom_base_one_cell_486/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_170 wl_0_28 sky130_rom_krom_rom_base_zero_cell_62/S
+ sky130_rom_krom_rom_base_one_cell_323/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_607 wl_0_14 sky130_rom_krom_rom_base_one_cell_704/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_629 wl_0_13 sky130_rom_krom_rom_base_one_cell_697/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_618 wl_0_13 sky130_rom_krom_rom_base_one_cell_683/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_181 wl_0_28 sky130_rom_krom_rom_base_zero_cell_77/S
+ sky130_rom_krom_rom_base_one_cell_220/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_192 wl_0_28 sky130_rom_krom_rom_base_one_cell_55/S
+ sky130_rom_krom_rom_base_one_cell_230/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_459 wl_0_18 sky130_rom_krom_rom_base_one_cell_515/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_448 wl_0_18 sky130_rom_krom_rom_base_one_cell_500/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_437 wl_0_18 sky130_rom_krom_rom_base_one_cell_491/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_426 wl_0_19 sky130_rom_krom_rom_base_one_cell_482/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_415 wl_0_19 sky130_rom_krom_rom_base_one_cell_537/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_404 wl_0_19 sky130_rom_krom_rom_base_one_cell_462/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_906 wl_0_4 sky130_rom_krom_rom_base_one_cell_906/D
+ sky130_rom_krom_rom_base_one_cell_906/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_917 wl_0_4 sky130_rom_krom_rom_base_one_cell_917/D
+ sky130_rom_krom_rom_base_one_cell_975/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_928 wl_0_3 sky130_rom_krom_rom_base_one_cell_928/D
+ bl_0_57 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_939 wl_0_3 sky130_rom_krom_rom_base_one_cell_939/D
+ sky130_rom_krom_rom_base_one_cell_939/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_960 wl_0_3 sky130_rom_krom_rom_base_one_cell_988/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_971 wl_0_2 sky130_rom_krom_rom_base_one_cell_936/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_982 wl_0_2 bl_0_22 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_993 wl_0_2 sky130_rom_krom_rom_base_one_cell_957/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_223 wl_0_24 sky130_rom_krom_rom_base_one_cell_377/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_201 wl_0_25 sky130_rom_krom_rom_base_one_cell_356/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_234 wl_0_24 sky130_rom_krom_rom_base_one_cell_329/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_245 wl_0_24 sky130_rom_krom_rom_base_one_cell_340/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_212 wl_0_25 sky130_rom_krom_rom_base_one_cell_341/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1004 wl_0_1 sky130_rom_krom_rom_base_one_cell_939/S
+ bl_0_38 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1048 wl_0_0 sky130_rom_krom_rom_base_one_cell_1048/D
+ bl_0_21 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1037 wl_0_0 sky130_rom_krom_rom_base_one_cell_933/S
+ bl_0_48 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1026 wl_0_1 sky130_rom_krom_rom_base_one_cell_955/S
+ sky130_rom_krom_rom_base_one_cell_1055/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1015 wl_0_1 sky130_rom_krom_rom_base_one_cell_919/S
+ sky130_rom_krom_rom_base_one_cell_1050/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_13 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_71/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_256 wl_0_23 sky130_rom_krom_rom_base_one_cell_372/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_267 wl_0_23 sky130_rom_krom_rom_base_one_cell_381/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_278 wl_0_23 sky130_rom_krom_rom_base_one_cell_387/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_289 wl_0_23 sky130_rom_krom_rom_base_one_cell_396/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_precharge_array_0 bl_0_0 bl_0_3 bl_0_5 bl_0_6 bl_0_10 bl_0_12
+ bl_0_17 bl_0_19 bl_0_21 bl_0_22 bl_0_24 bl_0_26 bl_0_28 bl_0_29 bl_0_30 bl_0_31
+ bl_0_35 bl_0_37 bl_0_38 bl_0_40 bl_0_42 bl_0_47 bl_0_49 bl_0_51 bl_0_52 bl_0_53
+ bl_0_56 bl_0_58 bl_0_59 bl_0_60 bl_0_61 bl_0_62 precharge bl_0_23 bl_0_33 bl_0_15
+ bl_0_45 bl_0_54 bl_0_8 bl_0_1 bl_0_63 bl_0_36 bl_0_4 bl_0_34 bl_0_27 bl_0_20 bl_0_50
+ bl_0_13 bl_0_43 bl_0_25 bl_0_18 bl_0_48 bl_0_11 bl_0_57 bl_0_41 bl_0_16 bl_0_46
+ vdd bl_0_9 bl_0_55 bl_0_39 bl_0_2 bl_0_32 bl_0_14 bl_0_44 bl_0_7 sky130_rom_krom_rom_precharge_array
Xsky130_rom_krom_rom_base_one_cell_24 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_24/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_35 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_35/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_46 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_90/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_57 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_57/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_68 wl_0_31 sky130_rom_krom_rom_base_one_cell_8/S
+ sky130_rom_krom_rom_base_one_cell_68/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_79 wl_0_31 sky130_rom_krom_rom_base_one_cell_79/D
+ sky130_rom_krom_rom_base_one_cell_79/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_758 wl_0_9 sky130_rom_krom_rom_base_one_cell_758/D
+ sky130_rom_krom_rom_base_one_cell_827/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_790 wl_0_8 sky130_rom_krom_rom_base_one_cell_820/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_747 wl_0_9 sky130_rom_krom_rom_base_one_cell_747/D
+ sky130_rom_krom_rom_base_one_cell_811/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_769 wl_0_8 sky130_rom_krom_rom_base_one_cell_769/D
+ sky130_rom_krom_rom_base_one_cell_836/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_736 wl_0_10 sky130_rom_krom_rom_base_one_cell_736/D
+ sky130_rom_krom_rom_base_one_cell_763/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_703 wl_0_11 sky130_rom_krom_rom_base_one_cell_703/D
+ sky130_rom_krom_rom_base_one_cell_761/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_725 wl_0_10 sky130_rom_krom_rom_base_one_cell_725/D
+ sky130_rom_krom_rom_base_one_cell_785/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_714 wl_0_10 sky130_rom_krom_rom_base_one_cell_714/D
+ sky130_rom_krom_rom_base_one_cell_746/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1003 wl_0_1 bl_0_41 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1047 wl_0_0 bl_0_11 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1036 wl_0_0 bl_0_30 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1025 wl_0_0 bl_0_51 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1014 wl_0_1 bl_0_17 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_511 wl_0_17 sky130_rom_krom_rom_base_one_cell_511/D
+ sky130_rom_krom_rom_base_one_cell_565/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_500 wl_0_17 sky130_rom_krom_rom_base_one_cell_500/D
+ sky130_rom_krom_rom_base_one_cell_533/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_599 wl_0_14 sky130_rom_krom_rom_base_one_cell_599/D
+ sky130_rom_krom_rom_base_one_cell_638/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_588 wl_0_14 sky130_rom_krom_rom_base_one_cell_588/D
+ sky130_rom_krom_rom_base_one_cell_621/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_577 wl_0_14 sky130_rom_krom_rom_base_one_cell_577/D
+ sky130_rom_krom_rom_base_one_cell_610/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_566 wl_0_15 sky130_rom_krom_rom_base_one_cell_566/D
+ sky130_rom_krom_rom_base_one_cell_661/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_555 wl_0_15 sky130_rom_krom_rom_base_one_cell_555/D
+ sky130_rom_krom_rom_base_one_cell_584/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_544 wl_0_16 sky130_rom_krom_rom_base_one_cell_544/D
+ sky130_rom_krom_rom_base_one_cell_632/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_533 wl_0_16 sky130_rom_krom_rom_base_one_cell_533/D
+ sky130_rom_krom_rom_base_one_cell_651/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_522 wl_0_16 sky130_rom_krom_rom_base_one_cell_522/D
+ sky130_rom_krom_rom_base_one_cell_551/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_1/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_330 wl_0_23 sky130_rom_krom_rom_base_one_cell_330/D
+ sky130_rom_krom_rom_base_one_cell_475/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_341 wl_0_23 sky130_rom_krom_rom_base_one_cell_341/D
+ sky130_rom_krom_rom_base_one_cell_366/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_352 wl_0_22 sky130_rom_krom_rom_base_one_cell_352/D
+ sky130_rom_krom_rom_base_one_cell_410/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_363 wl_0_22 sky130_rom_krom_rom_base_one_cell_363/D
+ sky130_rom_krom_rom_base_one_cell_422/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_374 wl_0_21 sky130_rom_krom_rom_base_one_cell_3/S
+ sky130_rom_krom_rom_base_one_cell_492/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_385 wl_0_21 sky130_rom_krom_rom_base_one_cell_385/D
+ sky130_rom_krom_rom_base_one_cell_415/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_396 wl_0_21 sky130_rom_krom_rom_base_one_cell_396/D
+ sky130_rom_krom_rom_base_one_cell_453/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_160 wl_0_29 sky130_rom_krom_rom_base_one_cell_160/D
+ sky130_rom_krom_rom_base_one_cell_196/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_171 wl_0_28 sky130_rom_krom_rom_base_zero_cell_7/S
+ sky130_rom_krom_rom_base_one_cell_268/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_182 wl_0_28 sky130_rom_krom_rom_base_zero_cell_78/S
+ sky130_rom_krom_rom_base_one_cell_221/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_193 wl_0_28 sky130_rom_krom_rom_base_one_cell_193/D
+ sky130_rom_krom_rom_base_one_cell_261/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_619 wl_0_13 sky130_rom_krom_rom_base_one_cell_654/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_608 wl_0_13 sky130_rom_krom_rom_base_one_cell_706/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_427 wl_0_19 sky130_rom_krom_rom_base_one_cell_515/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_416 wl_0_19 sky130_rom_krom_rom_base_one_cell_474/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_405 wl_0_19 sky130_rom_krom_rom_base_one_cell_463/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_449 wl_0_18 sky130_rom_krom_rom_base_one_cell_537/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_438 wl_0_18 sky130_rom_krom_rom_base_one_cell_522/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_907 wl_0_4 sky130_rom_krom_rom_base_one_cell_907/D
+ sky130_rom_krom_rom_base_one_cell_930/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_918 wl_0_4 sky130_rom_krom_rom_base_one_cell_918/D
+ sky130_rom_krom_rom_base_one_cell_947/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_929 wl_0_3 sky130_rom_krom_rom_base_one_cell_929/D
+ sky130_rom_krom_rom_base_one_cell_997/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_950 wl_0_3 sky130_rom_krom_rom_base_one_cell_979/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_961 wl_0_3 sky130_rom_krom_rom_base_one_cell_870/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_972 wl_0_2 bl_0_44 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_983 wl_0_2 sky130_rom_krom_rom_base_one_cell_948/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_0 wl_0_31 sky130_rom_krom_rom_base_one_cell_0/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_994 wl_0_1 bl_0_57 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_224 wl_0_24 sky130_rom_krom_rom_base_one_cell_348/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_202 wl_0_25 sky130_rom_krom_rom_base_one_cell_308/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_235 wl_0_24 sky130_rom_krom_rom_base_one_cell_330/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_246 wl_0_24 sky130_rom_krom_rom_base_one_cell_364/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_213 wl_0_25 sky130_rom_krom_rom_base_one_cell_368/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_257 wl_0_23 sky130_rom_krom_rom_base_one_cell_373/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_268 wl_0_23 sky130_rom_krom_rom_base_one_cell_351/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_279 wl_0_23 sky130_rom_krom_rom_base_one_cell_357/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1005 wl_0_1 sky130_rom_krom_rom_base_one_cell_968/S
+ bl_0_36 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1049 wl_0_0 sky130_rom_krom_rom_base_one_cell_1049/D
+ bl_0_20 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1038 wl_0_0 sky130_rom_krom_rom_base_one_cell_935/S
+ bl_0_46 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1027 wl_0_1 sky130_rom_krom_rom_base_one_cell_989/S
+ bl_0_2 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1016 wl_0_1 sky130_rom_krom_rom_base_one_cell_980/S
+ bl_0_16 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_14 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_6/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_25 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_76/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_36 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_82/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_47 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_91/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_58 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_58/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_69 wl_0_31 sky130_rom_krom_rom_base_one_cell_69/D
+ sky130_rom_krom_rom_base_one_cell_69/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_759 wl_0_9 sky130_rom_krom_rom_base_one_cell_759/D
+ sky130_rom_krom_rom_base_one_cell_794/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_791 wl_0_8 sky130_rom_krom_rom_base_one_cell_821/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_748 wl_0_9 sky130_rom_krom_rom_base_one_cell_748/D
+ sky130_rom_krom_rom_base_one_cell_778/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_780 wl_0_8 sky130_rom_krom_rom_base_one_cell_812/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_737 wl_0_9 sky130_rom_krom_rom_base_one_cell_737/D
+ sky130_rom_krom_rom_base_one_cell_764/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_704 wl_0_11 sky130_rom_krom_rom_base_one_cell_704/D
+ sky130_rom_krom_rom_base_one_cell_762/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_726 wl_0_10 sky130_rom_krom_rom_base_one_cell_726/D
+ sky130_rom_krom_rom_base_one_cell_823/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_715 wl_0_10 sky130_rom_krom_rom_base_one_cell_715/D
+ sky130_rom_krom_rom_base_one_cell_747/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1004 wl_0_1 bl_0_39 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1048 wl_0_0 bl_0_10 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1037 wl_0_0 bl_0_26 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1026 wl_0_0 bl_0_47 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1015 wl_0_1 bl_0_15 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_545 wl_0_16 sky130_rom_krom_rom_base_one_cell_545/D
+ sky130_rom_krom_rom_base_one_cell_596/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_534 wl_0_16 sky130_rom_krom_rom_base_one_cell_534/D
+ sky130_rom_krom_rom_base_one_cell_560/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_523 wl_0_16 sky130_rom_krom_rom_base_one_cell_523/D
+ sky130_rom_krom_rom_base_one_cell_552/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_512 wl_0_17 sky130_rom_krom_rom_base_one_cell_512/D
+ sky130_rom_krom_rom_base_one_cell_568/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_501 wl_0_17 sky130_rom_krom_rom_base_one_cell_501/D
+ sky130_rom_krom_rom_base_one_cell_534/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_589 wl_0_14 sky130_rom_krom_rom_base_one_cell_589/D
+ sky130_rom_krom_rom_base_one_cell_678/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_578 wl_0_14 sky130_rom_krom_rom_base_one_cell_578/D
+ sky130_rom_krom_rom_base_one_cell_611/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_567 wl_0_15 sky130_rom_krom_rom_base_one_cell_567/D
+ sky130_rom_krom_rom_base_one_cell_631/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_556 wl_0_15 sky130_rom_krom_rom_base_one_cell_556/D
+ sky130_rom_krom_rom_base_one_cell_618/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_90 wl_0_29 sky130_rom_krom_rom_base_zero_cell_90/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_2 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_2/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_320 wl_0_23 sky130_rom_krom_rom_base_one_cell_320/D
+ sky130_rom_krom_rom_base_one_cell_346/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_331 wl_0_23 sky130_rom_krom_rom_base_one_cell_331/D
+ sky130_rom_krom_rom_base_one_cell_358/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_342 wl_0_23 sky130_rom_krom_rom_base_one_cell_342/D
+ sky130_rom_krom_rom_base_one_cell_602/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_353 wl_0_22 sky130_rom_krom_rom_base_one_cell_353/D
+ sky130_rom_krom_rom_base_one_cell_383/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_364 wl_0_22 sky130_rom_krom_rom_base_one_cell_364/D
+ sky130_rom_krom_rom_base_one_cell_394/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_375 wl_0_21 sky130_rom_krom_rom_base_one_cell_375/D
+ sky130_rom_krom_rom_base_one_cell_434/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_386 wl_0_21 sky130_rom_krom_rom_base_one_cell_386/D
+ sky130_rom_krom_rom_base_one_cell_416/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_397 wl_0_21 sky130_rom_krom_rom_base_one_cell_397/D
+ sky130_rom_krom_rom_base_one_cell_488/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_609 wl_0_13 sky130_rom_krom_rom_base_one_cell_708/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_150 wl_0_29 sky130_rom_krom_rom_base_one_cell_150/D
+ sky130_rom_krom_rom_base_one_cell_215/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_161 wl_0_29 sky130_rom_krom_rom_base_one_cell_161/D
+ sky130_rom_krom_rom_base_one_cell_344/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_172 wl_0_28 sky130_rom_krom_rom_base_one_cell_172/D
+ sky130_rom_krom_rom_base_one_cell_208/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_183 wl_0_28 sky130_rom_krom_rom_base_zero_cell_79/S
+ sky130_rom_krom_rom_base_one_cell_222/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_194 wl_0_28 sky130_rom_krom_rom_base_zero_cell_92/S
+ sky130_rom_krom_rom_base_one_cell_262/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_439 wl_0_18 sky130_rom_krom_rom_base_one_cell_492/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_428 wl_0_19 sky130_rom_krom_rom_base_one_cell_483/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_417 wl_0_19 sky130_rom_krom_rom_base_one_cell_507/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_406 wl_0_19 sky130_rom_krom_rom_base_one_cell_466/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_908 wl_0_4 sky130_rom_krom_rom_base_one_cell_908/D
+ sky130_rom_krom_rom_base_one_cell_931/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_919 wl_0_4 sky130_rom_krom_rom_base_one_cell_919/D
+ sky130_rom_krom_rom_base_one_cell_919/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_940 wl_0_3 sky130_rom_krom_rom_base_one_cell_883/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_951 wl_0_3 sky130_rom_krom_rom_base_one_cell_919/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_962 wl_0_2 sky130_rom_krom_rom_base_one_cell_995/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_973 wl_0_2 sky130_rom_krom_rom_base_one_cell_937/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_984 wl_0_2 bl_0_19 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_995 wl_0_1 bl_0_55 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1 wl_0_31 sky130_rom_krom_rom_base_one_cell_1/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1006 wl_0_1 sky130_rom_krom_rom_base_one_cell_969/S
+ sky130_rom_krom_rom_base_one_cell_1041/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1017 wl_0_1 sky130_rom_krom_rom_base_one_cell_952/S
+ sky130_rom_krom_rom_base_one_cell_1051/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_225 wl_0_24 sky130_rom_krom_rom_base_one_cell_379/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_236 wl_0_24 sky130_rom_krom_rom_base_one_cell_387/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_203 wl_0_25 sky130_rom_krom_rom_base_one_cell_311/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_247 wl_0_24 sky130_rom_krom_rom_base_one_cell_395/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_214 wl_0_25 sky130_rom_krom_rom_base_one_cell_343/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_258 wl_0_23 sky130_rom_krom_rom_base_one_cell_345/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_269 wl_0_23 sky130_rom_krom_rom_base_one_cell_352/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1039 wl_0_0 sky130_rom_krom_rom_base_one_cell_1039/D
+ bl_0_45 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1028 wl_0_1 sky130_rom_krom_rom_base_one_cell_870/S
+ sky130_rom_krom_rom_base_one_cell_1056/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_15 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_72/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_26 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_26/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_37 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_37/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_48 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_92/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_59 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_99/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_705 wl_0_11 sky130_rom_krom_rom_base_one_cell_705/D
+ sky130_rom_krom_rom_base_one_cell_736/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_727 wl_0_10 sky130_rom_krom_rom_base_one_cell_727/D
+ sky130_rom_krom_rom_base_one_cell_787/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_716 wl_0_10 sky130_rom_krom_rom_base_one_cell_716/D
+ sky130_rom_krom_rom_base_one_cell_748/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_770 wl_0_9 sky130_rom_krom_rom_base_one_cell_796/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_792 wl_0_8 sky130_rom_krom_rom_base_one_cell_822/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_749 wl_0_9 sky130_rom_krom_rom_base_one_cell_749/D
+ sky130_rom_krom_rom_base_one_cell_845/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_781 wl_0_8 sky130_rom_krom_rom_base_one_cell_845/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_738 wl_0_9 sky130_rom_krom_rom_base_one_cell_738/D
+ sky130_rom_krom_rom_base_one_cell_767/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1005 wl_0_1 bl_0_37 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1049 wl_0_0 bl_0_9 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1038 wl_0_0 bl_0_25 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1027 wl_0_0 bl_0_44 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1016 wl_0_1 bl_0_13 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_579 wl_0_14 sky130_rom_krom_rom_base_one_cell_579/D
+ sky130_rom_krom_rom_base_one_cell_706/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_568 wl_0_15 sky130_rom_krom_rom_base_one_cell_568/D
+ sky130_rom_krom_rom_base_one_cell_594/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_557 wl_0_15 sky130_rom_krom_rom_base_one_cell_557/D
+ sky130_rom_krom_rom_base_one_cell_585/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_546 wl_0_16 sky130_rom_krom_rom_base_one_cell_546/D
+ sky130_rom_krom_rom_base_one_cell_634/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_535 wl_0_16 sky130_rom_krom_rom_base_one_cell_535/D
+ sky130_rom_krom_rom_base_one_cell_652/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_524 wl_0_16 sky130_rom_krom_rom_base_one_cell_524/D
+ sky130_rom_krom_rom_base_one_cell_613/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_513 wl_0_17 sky130_rom_krom_rom_base_one_cell_513/D
+ sky130_rom_krom_rom_base_one_cell_595/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_502 wl_0_17 sky130_rom_krom_rom_base_one_cell_502/D
+ sky130_rom_krom_rom_base_one_cell_561/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_80 wl_0_29 sky130_rom_krom_rom_base_one_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_91 wl_0_29 sky130_rom_krom_rom_base_one_cell_57/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_3 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_310 wl_0_24 sky130_rom_krom_rom_base_one_cell_310/D
+ sky130_rom_krom_rom_base_one_cell_331/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_321 wl_0_23 sky130_rom_krom_rom_base_one_cell_321/D
+ sky130_rom_krom_rom_base_one_cell_375/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_332 wl_0_23 sky130_rom_krom_rom_base_one_cell_332/D
+ sky130_rom_krom_rom_base_one_cell_478/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_343 wl_0_23 sky130_rom_krom_rom_base_one_cell_343/D
+ sky130_rom_krom_rom_base_one_cell_429/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_354 wl_0_22 sky130_rom_krom_rom_base_one_cell_354/D
+ sky130_rom_krom_rom_base_one_cell_384/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_365 wl_0_22 sky130_rom_krom_rom_base_one_cell_365/D
+ sky130_rom_krom_rom_base_one_cell_427/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_376 wl_0_21 sky130_rom_krom_rom_base_one_cell_376/D
+ sky130_rom_krom_rom_base_one_cell_404/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_387 wl_0_21 sky130_rom_krom_rom_base_one_cell_387/D
+ sky130_rom_krom_rom_base_one_cell_591/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_398 wl_0_21 sky130_rom_krom_rom_base_one_cell_398/D
+ sky130_rom_krom_rom_base_one_cell_454/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_140 wl_0_30 sky130_rom_krom_rom_base_one_cell_140/D
+ sky130_rom_krom_rom_base_one_cell_161/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_151 wl_0_29 sky130_rom_krom_rom_base_one_cell_151/D
+ sky130_rom_krom_rom_base_one_cell_179/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_162 wl_0_28 sky130_rom_krom_rom_base_zero_cell_51/S
+ sky130_rom_krom_rom_base_one_cell_197/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_173 wl_0_28 sky130_rom_krom_rom_base_one_cell_173/D
+ sky130_rom_krom_rom_base_one_cell_209/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_184 wl_0_28 sky130_rom_krom_rom_base_one_cell_87/S
+ sky130_rom_krom_rom_base_one_cell_223/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_195 wl_0_28 sky130_rom_krom_rom_base_zero_cell_93/S
+ sky130_rom_krom_rom_base_one_cell_232/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_429 wl_0_19 sky130_rom_krom_rom_base_one_cell_570/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_418 wl_0_19 sky130_rom_krom_rom_base_one_cell_475/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_407 wl_0_19 sky130_rom_krom_rom_base_one_cell_530/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_909 wl_0_4 sky130_rom_krom_rom_base_one_cell_909/D
+ sky130_rom_krom_rom_base_one_cell_932/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_2 wl_0_31 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_930 wl_0_3 sky130_rom_krom_rom_base_one_cell_959/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_941 wl_0_3 bl_0_39 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_952 wl_0_3 sky130_rom_krom_rom_base_one_cell_980/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_963 wl_0_2 bl_0_57 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_974 wl_0_2 sky130_rom_krom_rom_base_one_cell_882/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_985 wl_0_2 sky130_rom_krom_rom_base_one_cell_919/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_996 wl_0_1 sky130_rom_krom_rom_base_one_cell_906/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1007 wl_0_1 sky130_rom_krom_rom_base_one_cell_913/S
+ sky130_rom_krom_rom_base_one_cell_1042/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1029 wl_0_1 sky130_rom_krom_rom_base_one_cell_957/S
+ bl_0_0 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1018 wl_0_1 sky130_rom_krom_rom_base_one_cell_983/S
+ sky130_rom_krom_rom_base_one_cell_1052/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_226 wl_0_24 sky130_rom_krom_rom_base_one_cell_323/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_237 wl_0_24 sky130_rom_krom_rom_base_one_cell_332/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_204 wl_0_25 sky130_rom_krom_rom_base_one_cell_360/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_248 wl_0_24 sky130_rom_krom_rom_base_one_cell_396/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_215 wl_0_25 sky130_rom_krom_rom_base_one_cell_318/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_259 wl_0_23 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_16 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_27 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_27/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_38 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_83/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_49 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_93/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_739 wl_0_9 sky130_rom_krom_rom_base_one_cell_739/D
+ sky130_rom_krom_rom_base_one_cell_768/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_728 wl_0_10 sky130_rom_krom_rom_base_one_cell_728/D
+ sky130_rom_krom_rom_base_one_cell_859/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_717 wl_0_10 sky130_rom_krom_rom_base_one_cell_717/D
+ sky130_rom_krom_rom_base_one_cell_749/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_706 wl_0_10 sky130_rom_krom_rom_base_one_cell_706/D
+ sky130_rom_krom_rom_base_one_cell_766/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_771 wl_0_9 sky130_rom_krom_rom_base_one_cell_799/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_760 wl_0_9 sky130_rom_krom_rom_base_one_cell_823/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_793 wl_0_8 sky130_rom_krom_rom_base_one_cell_823/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_782 wl_0_8 sky130_rom_krom_rom_base_one_cell_884/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1006 wl_0_1 sky130_rom_krom_rom_base_one_cell_942/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1028 wl_0_0 bl_0_43 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1017 wl_0_1 sky130_rom_krom_rom_base_one_cell_921/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1039 wl_0_0 bl_0_24 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_590 wl_0_14 sky130_rom_krom_rom_base_one_cell_626/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_569 wl_0_15 sky130_rom_krom_rom_base_one_cell_569/D
+ sky130_rom_krom_rom_base_one_cell_633/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_558 wl_0_15 sky130_rom_krom_rom_base_one_cell_558/D
+ sky130_rom_krom_rom_base_one_cell_586/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_547 wl_0_16 sky130_rom_krom_rom_base_one_cell_547/D
+ sky130_rom_krom_rom_base_one_cell_605/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_536 wl_0_16 sky130_rom_krom_rom_base_one_cell_536/D
+ sky130_rom_krom_rom_base_one_cell_562/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_525 wl_0_16 sky130_rom_krom_rom_base_one_cell_525/D
+ sky130_rom_krom_rom_base_one_cell_708/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_514 wl_0_17 sky130_rom_krom_rom_base_one_cell_514/D
+ sky130_rom_krom_rom_base_one_cell_569/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_503 wl_0_17 sky130_rom_krom_rom_base_one_cell_503/D
+ sky130_rom_krom_rom_base_one_cell_536/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_70 wl_0_29 sky130_rom_krom_rom_base_zero_cell_70/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_81 wl_0_29 sky130_rom_krom_rom_base_zero_cell_81/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_92 wl_0_29 sky130_rom_krom_rom_base_zero_cell_92/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_4 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_4/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_300 wl_0_24 sky130_rom_krom_rom_base_one_cell_300/D
+ sky130_rom_krom_rom_base_one_cell_352/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_311 wl_0_24 sky130_rom_krom_rom_base_one_cell_311/D
+ sky130_rom_krom_rom_base_one_cell_359/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_322 wl_0_23 sky130_rom_krom_rom_base_one_cell_322/D
+ sky130_rom_krom_rom_base_one_cell_407/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_333 wl_0_23 sky130_rom_krom_rom_base_one_cell_333/D
+ sky130_rom_krom_rom_base_one_cell_361/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_344 wl_0_23 sky130_rom_krom_rom_base_one_cell_344/D
+ sky130_rom_krom_rom_base_one_cell_371/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_355 wl_0_22 sky130_rom_krom_rom_base_one_cell_355/D
+ sky130_rom_krom_rom_base_one_cell_444/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_366 wl_0_22 sky130_rom_krom_rom_base_one_cell_366/D
+ sky130_rom_krom_rom_base_one_cell_397/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_377 wl_0_21 sky130_rom_krom_rom_base_one_cell_377/D
+ sky130_rom_krom_rom_base_one_cell_405/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_388 wl_0_21 sky130_rom_krom_rom_base_one_cell_388/D
+ sky130_rom_krom_rom_base_one_cell_477/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_399 wl_0_21 sky130_rom_krom_rom_base_one_cell_399/D
+ sky130_rom_krom_rom_base_one_cell_428/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_130 wl_0_30 sky130_rom_krom_rom_base_one_cell_92/S
+ sky130_rom_krom_rom_base_zero_cell_85/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_141 wl_0_29 sky130_rom_krom_rom_base_one_cell_64/S
+ sky130_rom_krom_rom_base_one_cell_164/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_152 wl_0_29 sky130_rom_krom_rom_base_one_cell_152/D
+ sky130_rom_krom_rom_base_one_cell_251/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_163 wl_0_28 sky130_rom_krom_rom_base_one_cell_1/S
+ sky130_rom_krom_rom_base_one_cell_198/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_174 wl_0_28 sky130_rom_krom_rom_base_zero_cell_67/S
+ sky130_rom_krom_rom_base_one_cell_210/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_185 wl_0_28 sky130_rom_krom_rom_base_zero_cell_81/S
+ sky130_rom_krom_rom_base_one_cell_224/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_196 wl_0_28 sky130_rom_krom_rom_base_one_cell_196/D
+ sky130_rom_krom_rom_base_one_cell_233/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_419 wl_0_19 sky130_rom_krom_rom_base_one_cell_591/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_408 wl_0_19 sky130_rom_krom_rom_base_one_cell_587/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_920 wl_0_4 sky130_rom_krom_rom_base_one_cell_951/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_931 wl_0_3 sky130_rom_krom_rom_base_one_cell_960/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_3 wl_0_31 sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_942 wl_0_3 sky130_rom_krom_rom_base_one_cell_969/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_953 wl_0_3 sky130_rom_krom_rom_base_one_cell_982/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_964 wl_0_2 bl_0_55 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_975 wl_0_2 sky130_rom_krom_rom_base_one_cell_883/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_986 wl_0_2 bl_0_17 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_997 wl_0_1 bl_0_52 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_227 wl_0_24 sky130_rom_krom_rom_base_one_cell_381/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_205 wl_0_25 sky130_rom_krom_rom_base_one_cell_312/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_216 wl_0_25 sky130_rom_krom_rom_base_one_cell_319/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1008 wl_0_1 sky130_rom_krom_rom_base_one_cell_972/S
+ bl_0_30 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1019 wl_0_1 sky130_rom_krom_rom_base_one_cell_984/S
+ bl_0_11 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_238 wl_0_24 sky130_rom_krom_rom_base_one_cell_360/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_249 wl_0_24 sky130_rom_krom_rom_base_one_cell_341/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_17 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_8/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_28 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_28/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_39 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_84/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_761 wl_0_9 sky130_rom_krom_rom_base_one_cell_787/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_750 wl_0_9 sky130_rom_krom_rom_base_one_cell_782/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_783 wl_0_8 sky130_rom_krom_rom_base_one_cell_886/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_772 wl_0_8 sky130_rom_krom_rom_base_one_cell_871/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_729 wl_0_10 sky130_rom_krom_rom_base_one_cell_729/D
+ sky130_rom_krom_rom_base_one_cell_788/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_718 wl_0_10 sky130_rom_krom_rom_base_one_cell_718/D
+ sky130_rom_krom_rom_base_one_cell_780/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_707 wl_0_10 sky130_rom_krom_rom_base_one_cell_707/D
+ sky130_rom_krom_rom_base_one_cell_739/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_794 wl_0_8 sky130_rom_krom_rom_base_one_cell_859/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1007 wl_0_1 bl_0_32 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1029 wl_0_0 bl_0_41 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1018 wl_0_0 bl_0_62 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_591 wl_0_14 sky130_rom_krom_rom_base_one_cell_654/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_580 wl_0_14 sky130_rom_krom_rom_base_one_cell_616/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_559 wl_0_15 sky130_rom_krom_rom_base_one_cell_559/D
+ sky130_rom_krom_rom_base_one_cell_588/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_548 wl_0_16 sky130_rom_krom_rom_base_one_cell_548/D
+ sky130_rom_krom_rom_base_one_cell_574/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_537 wl_0_16 sky130_rom_krom_rom_base_one_cell_537/D
+ sky130_rom_krom_rom_base_one_cell_625/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_526 wl_0_16 sky130_rom_krom_rom_base_one_cell_526/D
+ sky130_rom_krom_rom_base_one_cell_582/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_515 wl_0_17 sky130_rom_krom_rom_base_one_cell_515/D
+ sky130_rom_krom_rom_base_one_cell_545/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_504 wl_0_17 sky130_rom_krom_rom_base_one_cell_504/D
+ sky130_rom_krom_rom_base_one_cell_626/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_60 wl_0_29 sky130_rom_krom_rom_base_zero_cell_60/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_71 wl_0_29 sky130_rom_krom_rom_base_one_cell_78/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_82 wl_0_29 sky130_rom_krom_rom_base_zero_cell_82/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_93 wl_0_29 sky130_rom_krom_rom_base_zero_cell_93/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_5 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_301 wl_0_24 sky130_rom_krom_rom_base_one_cell_301/D
+ sky130_rom_krom_rom_base_one_cell_382/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_312 wl_0_24 sky130_rom_krom_rom_base_one_cell_312/D
+ sky130_rom_krom_rom_base_one_cell_333/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_323 wl_0_23 sky130_rom_krom_rom_base_one_cell_323/D
+ sky130_rom_krom_rom_base_one_cell_350/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_334 wl_0_23 sky130_rom_krom_rom_base_one_cell_334/D
+ sky130_rom_krom_rom_base_one_cell_362/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_345 wl_0_22 sky130_rom_krom_rom_base_one_cell_345/D
+ sky130_rom_krom_rom_base_one_cell_522/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_356 wl_0_22 sky130_rom_krom_rom_base_one_cell_356/D
+ sky130_rom_krom_rom_base_one_cell_385/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_367 wl_0_22 sky130_rom_krom_rom_base_one_cell_367/D
+ sky130_rom_krom_rom_base_one_cell_603/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_378 wl_0_21 sky130_rom_krom_rom_base_one_cell_378/D
+ sky130_rom_krom_rom_base_one_cell_437/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_389 wl_0_21 sky130_rom_krom_rom_base_one_cell_389/D
+ sky130_rom_krom_rom_base_one_cell_479/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_890 wl_0_5 sky130_rom_krom_rom_base_one_cell_890/D
+ sky130_rom_krom_rom_base_one_cell_946/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_120 wl_0_30 sky130_rom_krom_rom_base_one_cell_82/S
+ sky130_rom_krom_rom_base_one_cell_152/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_131 wl_0_30 sky130_rom_krom_rom_base_one_cell_93/S
+ sky130_rom_krom_rom_base_zero_cell_86/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_142 wl_0_29 sky130_rom_krom_rom_base_one_cell_9/S
+ sky130_rom_krom_rom_base_one_cell_167/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_153 wl_0_29 sky130_rom_krom_rom_base_one_cell_153/D
+ sky130_rom_krom_rom_base_one_cell_281/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_164 wl_0_28 sky130_rom_krom_rom_base_one_cell_164/D
+ sky130_rom_krom_rom_base_one_cell_294/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_175 wl_0_28 sky130_rom_krom_rom_base_one_cell_175/D
+ sky130_rom_krom_rom_base_one_cell_273/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_186 wl_0_28 sky130_rom_krom_rom_base_zero_cell_82/S
+ sky130_rom_krom_rom_base_one_cell_255/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_197 wl_0_27 sky130_rom_krom_rom_base_one_cell_197/D
+ sky130_rom_krom_rom_base_one_cell_263/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_409 wl_0_19 sky130_rom_krom_rom_base_one_cell_468/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_910 wl_0_4 sky130_rom_krom_rom_base_one_cell_945/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_921 wl_0_4 sky130_rom_krom_rom_base_one_cell_982/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_932 wl_0_3 sky130_rom_krom_rom_base_one_cell_962/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_943 wl_0_3 sky130_rom_krom_rom_base_one_cell_913/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_954 wl_0_3 sky130_rom_krom_rom_base_one_cell_983/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_965 wl_0_2 sky130_rom_krom_rom_base_one_cell_997/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_4 wl_0_31 sky130_rom_krom_rom_base_one_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_976 wl_0_2 bl_0_39 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_987 wl_0_2 sky130_rom_krom_rom_base_one_cell_952/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_998 wl_0_1 sky130_rom_krom_rom_base_one_cell_966/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_228 wl_0_24 sky130_rom_krom_rom_base_one_cell_351/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_239 wl_0_24 sky130_rom_krom_rom_base_one_cell_334/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_206 wl_0_25 sky130_rom_krom_rom_base_one_cell_391/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_217 wl_0_25 sky130_rom_krom_rom_base_one_cell_344/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1009 wl_0_1 sky130_rom_krom_rom_base_one_cell_973/S
+ sky130_rom_krom_rom_base_one_cell_1045/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_18 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_9/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_29 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_29/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_795 wl_0_8 sky130_rom_krom_rom_base_one_cell_824/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_762 wl_0_9 sky130_rom_krom_rom_base_one_cell_859/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_751 wl_0_9 sky130_rom_krom_rom_base_one_cell_816/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_784 wl_0_8 sky130_rom_krom_rom_base_one_cell_815/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_740 wl_0_9 sky130_rom_krom_rom_base_one_cell_770/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_773 wl_0_8 sky130_rom_krom_rom_base_one_cell_801/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_719 wl_0_10 sky130_rom_krom_rom_base_one_cell_719/D
+ sky130_rom_krom_rom_base_one_cell_886/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_708 wl_0_10 sky130_rom_krom_rom_base_one_cell_708/D
+ sky130_rom_krom_rom_base_one_cell_740/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1008 wl_0_1 sky130_rom_krom_rom_base_one_cell_971/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1019 wl_0_0 bl_0_59 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_527 wl_0_16 sky130_rom_krom_rom_base_one_cell_527/D
+ sky130_rom_krom_rom_base_one_cell_616/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_516 wl_0_17 sky130_rom_krom_rom_base_one_cell_516/D
+ sky130_rom_krom_rom_base_one_cell_598/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_505 wl_0_17 sky130_rom_krom_rom_base_one_cell_505/D
+ sky130_rom_krom_rom_base_one_cell_538/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_592 wl_0_14 sky130_rom_krom_rom_base_one_cell_655/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_581 wl_0_14 sky130_rom_krom_rom_base_one_cell_618/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_570 wl_0_15 sky130_rom_krom_rom_base_one_cell_639/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_549 wl_0_15 sky130_rom_krom_rom_base_one_cell_549/D
+ sky130_rom_krom_rom_base_one_cell_575/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_538 wl_0_16 sky130_rom_krom_rom_base_one_cell_538/D
+ sky130_rom_krom_rom_base_one_cell_590/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_50 wl_0_30 sky130_rom_krom_rom_base_one_cell_58/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_61 wl_0_29 sky130_rom_krom_rom_base_zero_cell_61/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_72 wl_0_29 sky130_rom_krom_rom_base_one_cell_79/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_83 wl_0_29 sky130_rom_krom_rom_base_zero_cell_83/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_94 wl_0_28 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_6 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_6/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_302 wl_0_24 sky130_rom_krom_rom_base_one_cell_302/D
+ sky130_rom_krom_rom_base_one_cell_353/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_313 wl_0_24 sky130_rom_krom_rom_base_one_cell_313/D
+ sky130_rom_krom_rom_base_one_cell_335/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_324 wl_0_23 sky130_rom_krom_rom_base_one_cell_324/D
+ sky130_rom_krom_rom_base_one_cell_442/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_335 wl_0_23 sky130_rom_krom_rom_base_one_cell_335/D
+ sky130_rom_krom_rom_base_one_cell_419/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_346 wl_0_22 sky130_rom_krom_rom_base_one_cell_346/D
+ sky130_rom_krom_rom_base_one_cell_403/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_357 wl_0_22 sky130_rom_krom_rom_base_one_cell_357/D
+ sky130_rom_krom_rom_base_one_cell_417/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_368 wl_0_22 sky130_rom_krom_rom_base_one_cell_368/D
+ sky130_rom_krom_rom_base_one_cell_399/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_379 wl_0_21 sky130_rom_krom_rom_base_one_cell_379/D
+ sky130_rom_krom_rom_base_one_cell_466/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_891 wl_0_5 sky130_rom_krom_rom_base_one_cell_891/D
+ bl_0_22 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_880 wl_0_5 sky130_rom_krom_rom_base_one_cell_880/D
+ bl_0_44 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_110 wl_0_30 sky130_rom_krom_rom_base_zero_cell_8/S
+ sky130_rom_krom_rom_base_zero_cell_65/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_121 wl_0_30 sky130_rom_krom_rom_base_one_cell_37/S
+ sky130_rom_krom_rom_base_one_cell_153/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_132 wl_0_30 sky130_rom_krom_rom_base_one_cell_94/S
+ sky130_rom_krom_rom_base_one_cell_155/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_143 wl_0_29 sky130_rom_krom_rom_base_zero_cell_5/S
+ sky130_rom_krom_rom_base_zero_cell_98/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_154 wl_0_29 sky130_rom_krom_rom_base_one_cell_154/D
+ sky130_rom_krom_rom_base_one_cell_286/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_165 wl_0_28 sky130_rom_krom_rom_base_one_cell_67/S
+ sky130_rom_krom_rom_base_one_cell_376/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_176 wl_0_28 sky130_rom_krom_rom_base_one_cell_176/D
+ sky130_rom_krom_rom_base_one_cell_243/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_187 wl_0_28 sky130_rom_krom_rom_base_one_cell_91/S
+ sky130_rom_krom_rom_base_one_cell_256/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_198 wl_0_27 sky130_rom_krom_rom_base_one_cell_198/D
+ sky130_rom_krom_rom_base_one_cell_373/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_900 wl_0_4 sky130_rom_krom_rom_base_one_cell_936/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_911 wl_0_4 sky130_rom_krom_rom_base_one_cell_853/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_922 wl_0_4 sky130_rom_krom_rom_base_one_cell_983/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_933 wl_0_3 sky130_rom_krom_rom_base_one_cell_995/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_944 wl_0_3 sky130_rom_krom_rom_base_one_cell_970/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_955 wl_0_3 sky130_rom_krom_rom_base_one_cell_984/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_966 wl_0_2 sky130_rom_krom_rom_base_one_cell_906/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_977 wl_0_2 sky130_rom_krom_rom_base_one_cell_939/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_988 wl_0_2 sky130_rom_krom_rom_base_one_cell_921/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_999 wl_0_1 sky130_rom_krom_rom_base_one_cell_933/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_5 wl_0_31 sky130_rom_krom_rom_base_zero_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_218 wl_0_24 sky130_rom_krom_rom_base_one_cell_372/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_229 wl_0_24 sky130_rom_krom_rom_base_one_cell_325/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_207 wl_0_25 sky130_rom_krom_rom_base_zero_cell_83/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_19 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_73/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_709 wl_0_10 sky130_rom_krom_rom_base_one_cell_709/D
+ sky130_rom_krom_rom_base_one_cell_769/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_796 wl_0_8 sky130_rom_krom_rom_base_one_cell_862/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_763 wl_0_9 sky130_rom_krom_rom_base_one_cell_788/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_752 wl_0_9 sky130_rom_krom_rom_base_one_cell_817/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_785 wl_0_8 sky130_rom_krom_rom_base_one_cell_816/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_741 wl_0_9 sky130_rom_krom_rom_base_one_cell_771/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_774 wl_0_8 sky130_rom_krom_rom_base_one_cell_804/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_730 wl_0_10 sky130_rom_krom_rom_base_one_cell_795/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1009 wl_0_1 sky130_rom_krom_rom_base_one_cell_974/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_539 wl_0_16 sky130_rom_krom_rom_base_one_cell_539/D
+ sky130_rom_krom_rom_base_one_cell_685/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_528 wl_0_16 sky130_rom_krom_rom_base_one_cell_528/D
+ sky130_rom_krom_rom_base_one_cell_555/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_517 wl_0_17 sky130_rom_krom_rom_base_one_cell_517/D
+ sky130_rom_krom_rom_base_one_cell_571/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_506 wl_0_17 sky130_rom_krom_rom_base_one_cell_506/D
+ sky130_rom_krom_rom_base_one_cell_563/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_593 wl_0_14 sky130_rom_krom_rom_base_one_cell_685/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_582 wl_0_14 sky130_rom_krom_rom_base_one_cell_620/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_571 wl_0_15 sky130_rom_krom_rom_base_one_cell_602/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_560 wl_0_15 sky130_rom_krom_rom_base_one_cell_659/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_40 wl_0_30 sky130_rom_krom_rom_base_one_cell_78/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_51 wl_0_29 sky130_rom_krom_rom_base_zero_cell_51/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_62 wl_0_29 sky130_rom_krom_rom_base_zero_cell_62/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_73 wl_0_29 sky130_rom_krom_rom_base_one_cell_80/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_84 wl_0_29 sky130_rom_krom_rom_base_one_cell_91/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_95 wl_0_28 sky130_rom_krom_rom_base_one_cell_65/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_7 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_303 wl_0_24 sky130_rom_krom_rom_base_one_cell_303/D
+ sky130_rom_krom_rom_base_one_cell_324/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_314 wl_0_24 sky130_rom_krom_rom_base_one_cell_314/D
+ sky130_rom_krom_rom_base_one_cell_336/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_325 wl_0_23 sky130_rom_krom_rom_base_one_cell_325/D
+ sky130_rom_krom_rom_base_one_cell_499/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_336 wl_0_23 sky130_rom_krom_rom_base_one_cell_336/D
+ sky130_rom_krom_rom_base_one_cell_390/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_347 wl_0_22 sky130_rom_krom_rom_base_one_cell_347/D
+ sky130_rom_krom_rom_base_one_cell_435/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_358 wl_0_22 sky130_rom_krom_rom_base_one_cell_358/D
+ sky130_rom_krom_rom_base_one_cell_447/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_369 wl_0_22 sky130_rom_krom_rom_base_one_cell_369/D
+ sky130_rom_krom_rom_base_one_cell_400/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_390 wl_0_20 sky130_rom_krom_rom_base_one_cell_449/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_892 wl_0_5 sky130_rom_krom_rom_base_one_cell_892/D
+ sky130_rom_krom_rom_base_one_cell_949/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_881 wl_0_5 sky130_rom_krom_rom_base_one_cell_881/D
+ sky130_rom_krom_rom_base_one_cell_937/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_870 wl_0_6 sky130_rom_krom_rom_base_one_cell_870/D
+ sky130_rom_krom_rom_base_one_cell_870/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_100 wl_0_31 sky130_rom_krom_rom_base_one_cell_60/S
+ sky130_rom_krom_rom_base_one_cell_137/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_111 wl_0_30 sky130_rom_krom_rom_base_one_cell_73/S
+ sky130_rom_krom_rom_base_one_cell_145/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_122 wl_0_30 sky130_rom_krom_rom_base_one_cell_83/S
+ sky130_rom_krom_rom_base_zero_cell_76/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_133 wl_0_30 sky130_rom_krom_rom_base_one_cell_96/S
+ sky130_rom_krom_rom_base_zero_cell_88/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_144 wl_0_29 sky130_rom_krom_rom_base_zero_cell_9/S
+ sky130_rom_krom_rom_base_one_cell_172/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_155 wl_0_29 sky130_rom_krom_rom_base_one_cell_155/D
+ sky130_rom_krom_rom_base_one_cell_258/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_166 wl_0_28 sky130_rom_krom_rom_base_zero_cell_58/S
+ sky130_rom_krom_rom_base_one_cell_201/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_177 wl_0_28 sky130_rom_krom_rom_base_one_cell_177/D
+ sky130_rom_krom_rom_base_one_cell_213/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_188 wl_0_28 sky130_rom_krom_rom_base_zero_cell_85/S
+ sky130_rom_krom_rom_base_one_cell_225/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_199 wl_0_27 sky130_rom_krom_rom_base_one_cell_65/S
+ sky130_rom_krom_rom_base_one_cell_234/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_6 wl_0_31 sky130_rom_krom_rom_base_zero_cell_6/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_901 wl_0_4 bl_0_44 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_912 wl_0_4 sky130_rom_krom_rom_base_one_cell_946/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_923 wl_0_4 sky130_rom_krom_rom_base_one_cell_984/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_934 wl_0_3 sky130_rom_krom_rom_base_one_cell_963/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_945 wl_0_3 sky130_rom_krom_rom_base_one_cell_974/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_956 wl_0_3 sky130_rom_krom_rom_base_one_cell_985/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_967 wl_0_2 bl_0_52 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_978 wl_0_2 bl_0_37 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_989 wl_0_2 sky130_rom_krom_rom_base_one_cell_867/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_219 wl_0_24 sky130_rom_krom_rom_base_one_cell_373/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_208 wl_0_25 sky130_rom_krom_rom_base_one_cell_339/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_731 wl_0_10 sky130_rom_krom_rom_base_one_cell_796/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_720 wl_0_10 sky130_rom_krom_rom_base_one_cell_852/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_797 wl_0_8 sky130_rom_krom_rom_base_one_cell_827/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_764 wl_0_9 sky130_rom_krom_rom_base_one_cell_789/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_753 wl_0_9 sky130_rom_krom_rom_base_one_cell_783/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_786 wl_0_8 sky130_rom_krom_rom_base_one_cell_817/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_775 wl_0_8 sky130_rom_krom_rom_base_one_cell_806/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_742 wl_0_9 sky130_rom_krom_rom_base_one_cell_772/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_572 wl_0_15 sky130_rom_krom_rom_base_one_cell_603/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_561 wl_0_15 sky130_rom_krom_rom_base_one_cell_630/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_550 wl_0_15 sky130_rom_krom_rom_base_one_cell_651/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_529 wl_0_16 sky130_rom_krom_rom_base_one_cell_529/D
+ sky130_rom_krom_rom_base_one_cell_556/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_518 wl_0_17 sky130_rom_krom_rom_base_one_cell_518/D
+ sky130_rom_krom_rom_base_one_cell_572/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_507 wl_0_17 sky130_rom_krom_rom_base_one_cell_507/D
+ sky130_rom_krom_rom_base_one_cell_655/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_594 wl_0_14 sky130_rom_krom_rom_base_one_cell_628/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_583 wl_0_14 sky130_rom_krom_rom_base_one_cell_677/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_30 wl_0_30 sky130_rom_krom_rom_base_one_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_41 wl_0_30 sky130_rom_krom_rom_base_one_cell_79/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_52 wl_0_29 sky130_rom_krom_rom_base_one_cell_1/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_63 wl_0_29 sky130_rom_krom_rom_base_one_cell_72/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_74 wl_0_29 sky130_rom_krom_rom_base_zero_cell_74/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_85 wl_0_29 sky130_rom_krom_rom_base_zero_cell_85/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_96 wl_0_28 sky130_rom_krom_rom_base_zero_cell_96/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_8 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_8/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_304 wl_0_24 sky130_rom_krom_rom_base_one_cell_304/D
+ sky130_rom_krom_rom_base_one_cell_326/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_315 wl_0_24 sky130_rom_krom_rom_base_zero_cell_83/S
+ sky130_rom_krom_rom_base_one_cell_423/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_326 wl_0_23 sky130_rom_krom_rom_base_one_cell_326/D
+ sky130_rom_krom_rom_base_one_cell_411/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_337 wl_0_23 sky130_rom_krom_rom_base_one_cell_337/D
+ sky130_rom_krom_rom_base_one_cell_363/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_348 wl_0_22 sky130_rom_krom_rom_base_one_cell_348/D
+ sky130_rom_krom_rom_base_one_cell_406/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_359 wl_0_22 sky130_rom_krom_rom_base_one_cell_359/D
+ sky130_rom_krom_rom_base_one_cell_388/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_391 wl_0_20 sky130_rom_krom_rom_base_one_cell_451/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_380 wl_0_20 sky130_rom_krom_rom_base_one_cell_443/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_893 wl_0_5 sky130_rom_krom_rom_base_one_cell_893/D
+ sky130_rom_krom_rom_base_one_cell_950/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_882 wl_0_5 sky130_rom_krom_rom_base_one_cell_882/D
+ sky130_rom_krom_rom_base_one_cell_882/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_871 wl_0_5 sky130_rom_krom_rom_base_one_cell_871/D
+ sky130_rom_krom_rom_base_one_cell_901/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_860 wl_0_6 sky130_rom_krom_rom_base_one_cell_860/D
+ sky130_rom_krom_rom_base_one_cell_894/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_101 wl_0_31 sky130_rom_krom_rom_base_one_cell_61/S
+ sky130_rom_krom_rom_base_one_cell_138/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_112 wl_0_30 sky130_rom_krom_rom_base_one_cell_21/S
+ sky130_rom_krom_rom_base_zero_cell_66/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_123 wl_0_30 sky130_rom_krom_rom_base_one_cell_84/S
+ sky130_rom_krom_rom_base_zero_cell_77/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_134 wl_0_30 sky130_rom_krom_rom_base_one_cell_53/S
+ sky130_rom_krom_rom_base_one_cell_156/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_145 wl_0_29 sky130_rom_krom_rom_base_one_cell_145/D
+ sky130_rom_krom_rom_base_one_cell_240/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_156 wl_0_29 sky130_rom_krom_rom_base_one_cell_156/D
+ sky130_rom_krom_rom_base_one_cell_229/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_167 wl_0_28 sky130_rom_krom_rom_base_one_cell_167/D
+ sky130_rom_krom_rom_base_one_cell_202/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_178 wl_0_28 sky130_rom_krom_rom_base_zero_cell_70/S
+ sky130_rom_krom_rom_base_one_cell_214/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_189 wl_0_28 sky130_rom_krom_rom_base_zero_cell_86/S
+ sky130_rom_krom_rom_base_one_cell_226/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_690 wl_0_11 sky130_rom_krom_rom_base_one_cell_690/D
+ sky130_rom_krom_rom_base_one_cell_820/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_902 wl_0_4 sky130_rom_krom_rom_base_one_cell_937/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_913 wl_0_4 sky130_rom_krom_rom_base_one_cell_978/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_7 wl_0_31 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_924 wl_0_4 sky130_rom_krom_rom_base_one_cell_985/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_935 wl_0_3 bl_0_55 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_946 wl_0_3 sky130_rom_krom_rom_base_one_cell_975/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_957 wl_0_3 sky130_rom_krom_rom_base_one_cell_986/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_968 wl_0_2 sky130_rom_krom_rom_base_one_cell_933/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_979 wl_0_2 sky130_rom_krom_rom_base_one_cell_913/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_209 wl_0_25 sky130_rom_krom_rom_base_one_cell_316/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_765 wl_0_9 sky130_rom_krom_rom_base_one_cell_862/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_754 wl_0_9 sky130_rom_krom_rom_base_one_cell_888/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_743 wl_0_9 sky130_rom_krom_rom_base_one_cell_807/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_732 wl_0_10 sky130_rom_krom_rom_base_one_cell_761/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_721 wl_0_10 sky130_rom_krom_rom_base_one_cell_753/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_710 wl_0_10 sky130_rom_krom_rom_base_one_cell_773/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_798 wl_0_8 sky130_rom_krom_rom_base_one_cell_828/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_787 wl_0_8 sky130_rom_krom_rom_base_one_cell_888/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_776 wl_0_8 sky130_rom_krom_rom_base_one_cell_807/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_595 wl_0_14 sky130_rom_krom_rom_base_one_cell_658/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_584 wl_0_14 sky130_rom_krom_rom_base_one_cell_622/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_573 wl_0_15 sky130_rom_krom_rom_base_one_cell_604/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_562 wl_0_15 sky130_rom_krom_rom_base_one_cell_632/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_551 wl_0_15 sky130_rom_krom_rom_base_one_cell_652/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_540 wl_0_15 sky130_rom_krom_rom_base_one_cell_613/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_519 wl_0_17 sky130_rom_krom_rom_base_one_cell_519/D
+ sky130_rom_krom_rom_base_one_cell_601/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_508 wl_0_17 sky130_rom_krom_rom_base_one_cell_508/D
+ sky130_rom_krom_rom_base_one_cell_539/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_20 wl_0_31 sky130_rom_krom_rom_base_one_cell_53/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_31 wl_0_30 sky130_rom_krom_rom_base_zero_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_42 wl_0_30 sky130_rom_krom_rom_base_one_cell_80/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_53 wl_0_29 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_64 wl_0_29 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_75 wl_0_29 sky130_rom_krom_rom_base_one_cell_35/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_86 wl_0_29 sky130_rom_krom_rom_base_zero_cell_86/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_97 wl_0_28 sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_9 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_9/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_305 wl_0_24 sky130_rom_krom_rom_base_one_cell_305/D
+ sky130_rom_krom_rom_base_one_cell_412/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_316 wl_0_24 sky130_rom_krom_rom_base_one_cell_316/D
+ sky130_rom_krom_rom_base_one_cell_392/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_327 wl_0_23 sky130_rom_krom_rom_base_one_cell_327/D
+ sky130_rom_krom_rom_base_one_cell_470/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_338 wl_0_23 sky130_rom_krom_rom_base_one_cell_338/D
+ sky130_rom_krom_rom_base_one_cell_424/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_349 wl_0_22 sky130_rom_krom_rom_base_one_cell_349/D
+ sky130_rom_krom_rom_base_one_cell_378/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_392 wl_0_20 sky130_rom_krom_rom_base_one_cell_485/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_381 wl_0_20 sky130_rom_krom_rom_base_one_cell_444/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_370 wl_0_20 sky130_rom_krom_rom_base_one_cell_435/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_872 wl_0_5 sky130_rom_krom_rom_base_one_cell_872/D
+ sky130_rom_krom_rom_base_one_cell_902/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_861 wl_0_6 sky130_rom_krom_rom_base_one_cell_861/D
+ sky130_rom_krom_rom_base_one_cell_895/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_850 wl_0_6 sky130_rom_krom_rom_base_one_cell_850/D
+ sky130_rom_krom_rom_base_one_cell_887/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_894 wl_0_5 sky130_rom_krom_rom_base_one_cell_894/D
+ sky130_rom_krom_rom_base_one_cell_980/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_883 wl_0_5 sky130_rom_krom_rom_base_one_cell_883/D
+ sky130_rom_krom_rom_base_one_cell_883/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_102 wl_0_31 sky130_rom_krom_rom_base_one_cell_62/S
+ sky130_rom_krom_rom_base_one_cell_139/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_113 wl_0_30 sky130_rom_krom_rom_base_one_cell_22/S
+ sky130_rom_krom_rom_base_zero_cell_67/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_124 wl_0_30 sky130_rom_krom_rom_base_one_cell_85/S
+ sky130_rom_krom_rom_base_zero_cell_78/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_135 wl_0_30 sky130_rom_krom_rom_base_one_cell_98/S
+ sky130_rom_krom_rom_base_zero_cell_90/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_146 wl_0_29 sky130_rom_krom_rom_base_one_cell_74/S
+ sky130_rom_krom_rom_base_one_cell_173/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_157 wl_0_29 sky130_rom_krom_rom_base_one_cell_97/S
+ sky130_rom_krom_rom_base_one_cell_290/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_168 wl_0_28 sky130_rom_krom_rom_base_zero_cell_60/S
+ sky130_rom_krom_rom_base_one_cell_204/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_179 wl_0_28 sky130_rom_krom_rom_base_one_cell_179/D
+ sky130_rom_krom_rom_base_one_cell_216/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_691 wl_0_11 sky130_rom_krom_rom_base_one_cell_691/D
+ sky130_rom_krom_rom_base_one_cell_725/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_680 wl_0_11 sky130_rom_krom_rom_base_one_cell_680/D
+ sky130_rom_krom_rom_base_one_cell_884/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_903 wl_0_4 sky130_rom_krom_rom_base_one_cell_882/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_914 wl_0_4 bl_0_22 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_925 wl_0_4 sky130_rom_krom_rom_base_one_cell_986/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_936 wl_0_3 sky130_rom_krom_rom_base_one_cell_906/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_947 wl_0_3 sky130_rom_krom_rom_base_one_cell_853/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_8 wl_0_31 sky130_rom_krom_rom_base_zero_cell_8/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_958 wl_0_3 sky130_rom_krom_rom_base_one_cell_921/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_969 wl_0_2 sky130_rom_krom_rom_base_one_cell_934/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_766 wl_0_9 sky130_rom_krom_rom_base_one_cell_790/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_755 wl_0_9 sky130_rom_krom_rom_base_one_cell_852/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_788 wl_0_8 sky130_rom_krom_rom_base_one_cell_852/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_777 wl_0_8 sky130_rom_krom_rom_base_one_cell_808/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_744 wl_0_9 sky130_rom_krom_rom_base_one_cell_773/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_733 wl_0_10 sky130_rom_krom_rom_base_one_cell_762/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_700 wl_0_11 sky130_rom_krom_rom_base_one_cell_796/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_722 wl_0_10 sky130_rom_krom_rom_base_one_cell_784/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_711 wl_0_10 sky130_rom_krom_rom_base_one_cell_742/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_799 wl_0_8 sky130_rom_krom_rom_base_one_cell_900/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_509 wl_0_17 sky130_rom_krom_rom_base_one_cell_509/D
+ sky130_rom_krom_rom_base_one_cell_540/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_596 wl_0_14 sky130_rom_krom_rom_base_one_cell_659/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_585 wl_0_14 sky130_rom_krom_rom_base_one_cell_651/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_574 wl_0_15 sky130_rom_krom_rom_base_one_cell_605/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_563 wl_0_15 sky130_rom_krom_rom_base_one_cell_595/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_552 wl_0_15 sky130_rom_krom_rom_base_one_cell_625/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_541 wl_0_15 sky130_rom_krom_rom_base_one_cell_708/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_530 wl_0_16 sky130_rom_krom_rom_base_one_cell_572/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_10 wl_0_31 sky130_rom_krom_rom_base_one_cell_21/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_21 wl_0_31 sky130_rom_krom_rom_base_one_cell_55/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_32 wl_0_30 sky130_rom_krom_rom_base_one_cell_69/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_43 wl_0_30 sky130_rom_krom_rom_base_one_cell_35/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_54 wl_0_29 sky130_rom_krom_rom_base_one_cell_65/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_65 wl_0_29 sky130_rom_krom_rom_base_zero_cell_65/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_76 wl_0_29 sky130_rom_krom_rom_base_zero_cell_76/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_87 wl_0_29 sky130_rom_krom_rom_base_one_cell_95/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_98 wl_0_28 sky130_rom_krom_rom_base_zero_cell_98/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_306 wl_0_24 sky130_rom_krom_rom_base_one_cell_306/D
+ sky130_rom_krom_rom_base_one_cell_443/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_317 wl_0_24 sky130_rom_krom_rom_base_one_cell_317/D
+ sky130_rom_krom_rom_base_one_cell_365/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_328 wl_0_23 sky130_rom_krom_rom_base_one_cell_328/D
+ sky130_rom_krom_rom_base_one_cell_354/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_339 wl_0_23 sky130_rom_krom_rom_base_one_cell_339/D
+ sky130_rom_krom_rom_base_one_cell_425/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_360 wl_0_21 sky130_rom_krom_rom_base_one_cell_425/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_393 wl_0_20 sky130_rom_krom_rom_base_one_cell_486/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_382 wl_0_20 sky130_rom_krom_rom_base_one_cell_507/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_371 wl_0_20 sky130_rom_krom_rom_base_one_cell_437/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_895 wl_0_5 sky130_rom_krom_rom_base_one_cell_895/D
+ sky130_rom_krom_rom_base_one_cell_951/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_884 wl_0_5 sky130_rom_krom_rom_base_one_cell_884/D
+ sky130_rom_krom_rom_base_one_cell_911/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_873 wl_0_5 sky130_rom_krom_rom_base_one_cell_873/D
+ sky130_rom_krom_rom_base_one_cell_927/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_862 wl_0_6 sky130_rom_krom_rom_base_one_cell_862/D
+ sky130_rom_krom_rom_base_one_cell_982/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_851 wl_0_6 sky130_rom_krom_rom_base_one_cell_851/D
+ sky130_rom_krom_rom_base_one_cell_945/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_840 wl_0_6 sky130_rom_krom_rom_base_one_cell_840/D
+ sky130_rom_krom_rom_base_one_cell_934/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_103 wl_0_31 sky130_rom_krom_rom_base_one_cell_63/S
+ sky130_rom_krom_rom_base_one_cell_140/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_114 wl_0_30 sky130_rom_krom_rom_base_one_cell_24/S
+ sky130_rom_krom_rom_base_one_cell_148/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_125 wl_0_30 sky130_rom_krom_rom_base_one_cell_86/S
+ sky130_rom_krom_rom_base_zero_cell_79/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_136 wl_0_30 sky130_rom_krom_rom_base_one_cell_99/S
+ sky130_rom_krom_rom_base_one_cell_159/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_147 wl_0_29 sky130_rom_krom_rom_base_one_cell_75/S
+ sky130_rom_krom_rom_base_one_cell_175/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_158 wl_0_29 sky130_rom_krom_rom_base_one_cell_58/S
+ sky130_rom_krom_rom_base_one_cell_193/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_169 wl_0_28 sky130_rom_krom_rom_base_zero_cell_61/S
+ sky130_rom_krom_rom_base_one_cell_205/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_190 wl_0_25 sky130_rom_krom_rom_base_one_cell_377/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_692 wl_0_11 sky130_rom_krom_rom_base_one_cell_692/D
+ sky130_rom_krom_rom_base_one_cell_755/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_681 wl_0_11 sky130_rom_krom_rom_base_one_cell_681/D
+ sky130_rom_krom_rom_base_one_cell_750/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_670 wl_0_12 sky130_rom_krom_rom_base_one_cell_670/D
+ sky130_rom_krom_rom_base_one_cell_796/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_904 wl_0_4 sky130_rom_krom_rom_base_one_cell_883/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_915 wl_0_4 sky130_rom_krom_rom_base_one_cell_979/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_926 wl_0_4 sky130_rom_krom_rom_base_one_cell_953/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_937 wl_0_3 sky130_rom_krom_rom_base_one_cell_964/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_948 wl_0_3 sky130_rom_krom_rom_base_one_cell_978/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_959 wl_0_3 sky130_rom_krom_rom_base_one_cell_867/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_9 wl_0_31 sky130_rom_krom_rom_base_zero_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_767 wl_0_9 sky130_rom_krom_rom_base_one_cell_792/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_756 wl_0_9 sky130_rom_krom_rom_base_one_cell_784/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_789 wl_0_8 sky130_rom_krom_rom_base_one_cell_853/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_778 wl_0_8 sky130_rom_krom_rom_base_one_cell_810/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_745 wl_0_9 sky130_rom_krom_rom_base_one_cell_775/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_701 wl_0_11 sky130_rom_krom_rom_base_one_cell_799/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_734 wl_0_10 sky130_rom_krom_rom_base_one_cell_799/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_723 wl_0_10 sky130_rom_krom_rom_base_one_cell_820/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_712 wl_0_10 sky130_rom_krom_rom_base_one_cell_743/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_531 wl_0_16 sky130_rom_krom_rom_base_one_cell_573/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_520 wl_0_16 sky130_rom_krom_rom_base_one_cell_658/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_597 wl_0_14 sky130_rom_krom_rom_base_one_cell_630/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_586 wl_0_14 sky130_rom_krom_rom_base_one_cell_652/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_575 wl_0_15 sky130_rom_krom_rom_base_one_cell_704/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_564 wl_0_15 sky130_rom_krom_rom_base_one_cell_596/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_553 wl_0_15 sky130_rom_krom_rom_base_one_cell_626/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_542 wl_0_15 sky130_rom_krom_rom_base_one_cell_615/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_11 wl_0_31 sky130_rom_krom_rom_base_one_cell_22/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_22 wl_0_31 sky130_rom_krom_rom_base_one_cell_57/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_33 wl_0_30 sky130_rom_krom_rom_base_one_cell_72/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_44 wl_0_30 sky130_rom_krom_rom_base_one_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_55 wl_0_29 sky130_rom_krom_rom_base_zero_cell_96/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_66 wl_0_29 sky130_rom_krom_rom_base_zero_cell_66/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_77 wl_0_29 sky130_rom_krom_rom_base_zero_cell_77/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_88 wl_0_29 sky130_rom_krom_rom_base_zero_cell_88/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_99 wl_0_28 sky130_rom_krom_rom_base_one_cell_69/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_307 wl_0_24 sky130_rom_krom_rom_base_one_cell_307/D
+ sky130_rom_krom_rom_base_one_cell_414/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_318 wl_0_24 sky130_rom_krom_rom_base_one_cell_318/D
+ sky130_rom_krom_rom_base_one_cell_369/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_329 wl_0_23 sky130_rom_krom_rom_base_one_cell_329/D
+ sky130_rom_krom_rom_base_one_cell_386/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_350 wl_0_21 sky130_rom_krom_rom_base_one_cell_417/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_361 wl_0_21 sky130_rom_krom_rom_base_one_cell_427/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_372 wl_0_20 sky130_rom_krom_rom_base_one_cell_438/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_394 wl_0_20 sky130_rom_krom_rom_base_one_cell_453/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_383 wl_0_20 sky130_rom_krom_rom_base_one_cell_475/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_896 wl_0_5 sky130_rom_krom_rom_base_one_cell_896/D
+ sky130_rom_krom_rom_base_one_cell_920/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_885 wl_0_5 sky130_rom_krom_rom_base_one_cell_885/D
+ sky130_rom_krom_rom_base_one_cell_940/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_874 wl_0_5 sky130_rom_krom_rom_base_one_cell_874/D
+ sky130_rom_krom_rom_base_one_cell_995/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_863 wl_0_6 sky130_rom_krom_rom_base_one_cell_863/D
+ sky130_rom_krom_rom_base_one_cell_984/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_852 wl_0_6 sky130_rom_krom_rom_base_one_cell_852/D
+ sky130_rom_krom_rom_base_one_cell_889/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_841 wl_0_6 sky130_rom_krom_rom_base_one_cell_841/D
+ sky130_rom_krom_rom_base_one_cell_879/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_830 wl_0_7 sky130_rom_krom_rom_base_one_cell_830/D
+ sky130_rom_krom_rom_base_one_cell_869/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_104 wl_0_30 sky130_rom_krom_rom_base_one_cell_0/S
+ sky130_rom_krom_rom_base_zero_cell_51/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_115 wl_0_30 sky130_rom_krom_rom_base_one_cell_76/S
+ sky130_rom_krom_rom_base_zero_cell_68/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_126 wl_0_30 sky130_rom_krom_rom_base_one_cell_43/S
+ sky130_rom_krom_rom_base_zero_cell_81/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_137 wl_0_30 sky130_rom_krom_rom_base_one_cell_137/D
+ sky130_rom_krom_rom_base_zero_cell_92/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_148 wl_0_29 sky130_rom_krom_rom_base_one_cell_148/D
+ sky130_rom_krom_rom_base_one_cell_176/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_159 wl_0_29 sky130_rom_krom_rom_base_one_cell_159/D
+ sky130_rom_krom_rom_base_one_cell_368/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_180 wl_0_26 sky130_rom_krom_rom_base_one_cell_291/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_191 wl_0_25 sky130_rom_krom_rom_base_one_cell_348/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_693 wl_0_11 sky130_rom_krom_rom_base_one_cell_693/D
+ sky130_rom_krom_rom_base_one_cell_727/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_682 wl_0_11 sky130_rom_krom_rom_base_one_cell_682/D
+ sky130_rom_krom_rom_base_one_cell_719/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_671 wl_0_12 sky130_rom_krom_rom_base_one_cell_671/D
+ sky130_rom_krom_rom_base_one_cell_799/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_660 wl_0_12 sky130_rom_krom_rom_base_one_cell_660/D
+ sky130_rom_krom_rom_base_one_cell_690/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_905 wl_0_4 bl_0_39 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_916 wl_0_4 sky130_rom_krom_rom_base_one_cell_948/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_927 wl_0_4 sky130_rom_krom_rom_base_one_cell_867/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_938 wl_0_3 bl_0_44 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_949 wl_0_3 bl_0_22 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_490 wl_0_17 sky130_rom_krom_rom_base_one_cell_490/D
+ sky130_rom_krom_rom_base_one_cell_549/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_713 wl_0_10 sky130_rom_krom_rom_base_one_cell_745/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_702 wl_0_10 sky130_rom_krom_rom_base_one_cell_871/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_768 wl_0_9 sky130_rom_krom_rom_base_one_cell_793/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_757 wl_0_9 sky130_rom_krom_rom_base_one_cell_820/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_746 wl_0_9 sky130_rom_krom_rom_base_one_cell_812/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_779 wl_0_8 sky130_rom_krom_rom_base_one_cell_811/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_735 wl_0_9 sky130_rom_krom_rom_base_one_cell_871/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_724 wl_0_10 sky130_rom_krom_rom_base_one_cell_754/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_554 wl_0_15 sky130_rom_krom_rom_base_one_cell_590/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_543 wl_0_15 sky130_rom_krom_rom_base_one_cell_582/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_532 wl_0_16 sky130_rom_krom_rom_base_one_cell_601/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_521 wl_0_16 sky130_rom_krom_rom_base_one_cell_630/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_510 wl_0_16 sky130_rom_krom_rom_base_one_cell_620/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_598 wl_0_14 sky130_rom_krom_rom_base_one_cell_661/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_587 wl_0_14 sky130_rom_krom_rom_base_one_cell_623/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_576 wl_0_15 sky130_rom_krom_rom_base_one_cell_607/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_565 wl_0_15 sky130_rom_krom_rom_base_one_cell_634/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_12 wl_0_31 sky130_rom_krom_rom_base_one_cell_24/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_23 wl_0_31 sky130_rom_krom_rom_base_one_cell_58/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_34 wl_0_30 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_45 wl_0_30 sky130_rom_krom_rom_base_one_cell_91/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_56 wl_0_29 sky130_rom_krom_rom_base_one_cell_67/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_67 wl_0_29 sky130_rom_krom_rom_base_zero_cell_67/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_78 wl_0_29 sky130_rom_krom_rom_base_zero_cell_78/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_89 wl_0_29 sky130_rom_krom_rom_base_one_cell_55/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_308 wl_0_24 sky130_rom_krom_rom_base_one_cell_308/D
+ sky130_rom_krom_rom_base_one_cell_507/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_319 wl_0_24 sky130_rom_krom_rom_base_one_cell_319/D
+ sky130_rom_krom_rom_base_one_cell_370/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_340 wl_0_21 sky130_rom_krom_rom_base_one_cell_442/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_351 wl_0_21 sky130_rom_krom_rom_base_one_cell_447/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_362 wl_0_21 sky130_rom_krom_rom_base_one_cell_602/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_395 wl_0_20 sky130_rom_krom_rom_base_one_cell_488/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_384 wl_0_20 sky130_rom_krom_rom_base_one_cell_591/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_373 wl_0_20 sky130_rom_krom_rom_base_one_cell_466/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_831 wl_0_7 sky130_rom_krom_rom_base_one_cell_831/D
+ sky130_rom_krom_rom_base_one_cell_899/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_820 wl_0_7 sky130_rom_krom_rom_base_one_cell_820/D
+ sky130_rom_krom_rom_base_one_cell_855/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_897 wl_0_5 sky130_rom_krom_rom_base_one_cell_897/D
+ sky130_rom_krom_rom_base_one_cell_983/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_886 wl_0_5 sky130_rom_krom_rom_base_one_cell_886/D
+ sky130_rom_krom_rom_base_one_cell_912/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_875 wl_0_5 sky130_rom_krom_rom_base_one_cell_875/D
+ sky130_rom_krom_rom_base_one_cell_904/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_864 wl_0_6 sky130_rom_krom_rom_base_one_cell_864/D
+ sky130_rom_krom_rom_base_one_cell_985/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_853 wl_0_6 sky130_rom_krom_rom_base_one_cell_853/D
+ sky130_rom_krom_rom_base_one_cell_853/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_842 wl_0_6 sky130_rom_krom_rom_base_one_cell_842/D
+ sky130_rom_krom_rom_base_one_cell_881/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_105 wl_0_30 sky130_rom_krom_rom_base_one_cell_66/S
+ sky130_rom_krom_rom_base_zero_cell_96/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_116 wl_0_30 sky130_rom_krom_rom_base_one_cell_28/S
+ sky130_rom_krom_rom_base_zero_cell_70/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_127 wl_0_30 sky130_rom_krom_rom_base_one_cell_88/S
+ sky130_rom_krom_rom_base_zero_cell_82/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_138 wl_0_30 sky130_rom_krom_rom_base_one_cell_138/D
+ sky130_rom_krom_rom_base_zero_cell_93/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_149 wl_0_29 sky130_rom_krom_rom_base_one_cell_27/S
+ sky130_rom_krom_rom_base_one_cell_177/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_170 wl_0_26 sky130_rom_krom_rom_base_one_cell_282/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_181 wl_0_26 sky130_rom_krom_rom_base_one_cell_368/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_192 wl_0_25 sky130_rom_krom_rom_base_one_cell_297/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_672 wl_0_11 sky130_rom_krom_rom_base_one_cell_672/D
+ sky130_rom_krom_rom_base_one_cell_801/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_661 wl_0_12 sky130_rom_krom_rom_base_one_cell_661/D
+ sky130_rom_krom_rom_base_one_cell_724/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_650 wl_0_12 sky130_rom_krom_rom_base_one_cell_650/D
+ sky130_rom_krom_rom_base_one_cell_712/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_694 wl_0_11 sky130_rom_krom_rom_base_one_cell_694/D
+ sky130_rom_krom_rom_base_one_cell_728/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_683 wl_0_11 sky130_rom_krom_rom_base_one_cell_683/D
+ sky130_rom_krom_rom_base_one_cell_720/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_906 wl_0_4 sky130_rom_krom_rom_base_one_cell_940/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_917 wl_0_4 sky130_rom_krom_rom_base_one_cell_949/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_928 wl_0_4 sky130_rom_krom_rom_base_one_cell_954/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_939 wl_0_3 sky130_rom_krom_rom_base_one_cell_882/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_491 wl_0_17 sky130_rom_krom_rom_base_one_cell_491/D
+ sky130_rom_krom_rom_base_one_cell_521/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_480 wl_0_18 sky130_rom_krom_rom_base_one_cell_480/D
+ sky130_rom_krom_rom_base_one_cell_512/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_747 wl_0_9 sky130_rom_krom_rom_base_one_cell_884/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_736 wl_0_9 sky130_rom_krom_rom_base_one_cell_801/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_725 wl_0_10 sky130_rom_krom_rom_base_one_cell_755/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_714 wl_0_10 sky130_rom_krom_rom_base_one_cell_812/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_703 wl_0_10 sky130_rom_krom_rom_base_one_cell_737/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_769 wl_0_9 sky130_rom_krom_rom_base_one_cell_795/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_758 wl_0_9 sky130_rom_krom_rom_base_one_cell_821/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_588 wl_0_14 sky130_rom_krom_rom_base_one_cell_624/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_577 wl_0_14 sky130_rom_krom_rom_base_one_cell_613/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_566 wl_0_15 sky130_rom_krom_rom_base_one_cell_636/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_555 wl_0_15 sky130_rom_krom_rom_base_one_cell_655/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_544 wl_0_15 sky130_rom_krom_rom_base_one_cell_616/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_533 wl_0_16 sky130_rom_krom_rom_base_one_cell_639/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_522 wl_0_16 sky130_rom_krom_rom_base_one_cell_568/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_511 wl_0_16 sky130_rom_krom_rom_base_one_cell_587/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_500 wl_0_17 sky130_rom_krom_rom_base_one_cell_704/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_599 wl_0_14 sky130_rom_krom_rom_base_one_cell_631/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_13 wl_0_31 sky130_rom_krom_rom_base_one_cell_26/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_24 wl_0_30 sky130_rom_krom_rom_base_one_cell_1/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_35 wl_0_30 sky130_rom_krom_rom_base_zero_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_46 wl_0_30 sky130_rom_krom_rom_base_one_cell_95/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_57 wl_0_29 sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_68 wl_0_29 sky130_rom_krom_rom_base_zero_cell_68/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_79 wl_0_29 sky130_rom_krom_rom_base_zero_cell_79/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_309 wl_0_24 sky130_rom_krom_rom_base_one_cell_309/D
+ sky130_rom_krom_rom_base_one_cell_357/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_330 wl_0_22 sky130_rom_krom_rom_base_one_cell_602/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_341 wl_0_21 sky130_rom_krom_rom_base_one_cell_499/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_352 wl_0_21 sky130_rom_krom_rom_base_one_cell_478/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_363 wl_0_21 sky130_rom_krom_rom_base_one_cell_603/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_396 wl_0_20 sky130_rom_krom_rom_base_one_cell_454/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_385 wl_0_20 sky130_rom_krom_rom_base_one_cell_447/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_374 wl_0_20 sky130_rom_krom_rom_base_one_cell_440/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_854 wl_0_6 sky130_rom_krom_rom_base_one_cell_854/D
+ sky130_rom_krom_rom_base_one_cell_890/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_843 wl_0_6 sky130_rom_krom_rom_base_one_cell_843/D
+ sky130_rom_krom_rom_base_one_cell_882/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_832 wl_0_7 sky130_rom_krom_rom_base_one_cell_832/D
+ sky130_rom_krom_rom_base_one_cell_870/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_821 wl_0_7 sky130_rom_krom_rom_base_one_cell_821/D
+ sky130_rom_krom_rom_base_one_cell_856/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_810 wl_0_7 sky130_rom_krom_rom_base_one_cell_810/D
+ sky130_rom_krom_rom_base_one_cell_842/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_898 wl_0_5 sky130_rom_krom_rom_base_one_cell_898/D
+ sky130_rom_krom_rom_base_one_cell_953/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_887 wl_0_5 sky130_rom_krom_rom_base_one_cell_887/D
+ sky130_rom_krom_rom_base_one_cell_915/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_876 wl_0_5 sky130_rom_krom_rom_base_one_cell_876/D
+ bl_0_55 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_865 wl_0_6 sky130_rom_krom_rom_base_one_cell_865/D
+ sky130_rom_krom_rom_base_one_cell_921/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_106 wl_0_30 sky130_rom_krom_rom_base_one_cell_68/S
+ sky130_rom_krom_rom_base_zero_cell_58/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_117 wl_0_30 sky130_rom_krom_rom_base_one_cell_29/S
+ sky130_rom_krom_rom_base_one_cell_150/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_128 wl_0_30 sky130_rom_krom_rom_base_one_cell_89/S
+ sky130_rom_krom_rom_base_one_cell_154/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_139 wl_0_30 sky130_rom_krom_rom_base_one_cell_139/D
+ sky130_rom_krom_rom_base_one_cell_160/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_160 wl_0_26 sky130_rom_krom_rom_base_one_cell_268/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_171 wl_0_26 sky130_rom_krom_rom_base_one_cell_284/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_182 wl_0_26 sky130_rom_krom_rom_base_one_cell_318/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_193 wl_0_25 sky130_rom_krom_rom_base_one_cell_298/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_695 wl_0_11 sky130_rom_krom_rom_base_one_cell_695/D
+ sky130_rom_krom_rom_base_one_cell_756/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_684 wl_0_11 sky130_rom_krom_rom_base_one_cell_684/D
+ sky130_rom_krom_rom_base_one_cell_722/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_673 wl_0_11 sky130_rom_krom_rom_base_one_cell_673/D
+ sky130_rom_krom_rom_base_one_cell_738/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_662 wl_0_12 sky130_rom_krom_rom_base_one_cell_662/D
+ sky130_rom_krom_rom_base_one_cell_691/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_651 wl_0_12 sky130_rom_krom_rom_base_one_cell_651/D
+ sky130_rom_krom_rom_base_one_cell_812/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_640 wl_0_13 sky130_rom_krom_rom_base_one_cell_640/D
+ sky130_rom_krom_rom_base_one_cell_670/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_907 wl_0_4 sky130_rom_krom_rom_base_one_cell_941/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_918 wl_0_4 sky130_rom_krom_rom_base_one_cell_950/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_929 wl_0_4 sky130_rom_krom_rom_base_one_cell_870/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_492 wl_0_17 sky130_rom_krom_rom_base_one_cell_492/D
+ sky130_rom_krom_rom_base_one_cell_578/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_481 wl_0_18 sky130_rom_krom_rom_base_one_cell_481/D
+ sky130_rom_krom_rom_base_one_cell_544/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_470 wl_0_18 sky130_rom_krom_rom_base_one_cell_470/D
+ sky130_rom_krom_rom_base_one_cell_501/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_759 wl_0_9 sky130_rom_krom_rom_base_one_cell_785/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_748 wl_0_9 sky130_rom_krom_rom_base_one_cell_780/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_737 wl_0_9 sky130_rom_krom_rom_base_one_cell_765/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_726 wl_0_10 sky130_rom_krom_rom_base_one_cell_756/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_715 wl_0_10 sky130_rom_krom_rom_base_one_cell_884/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_704 wl_0_10 sky130_rom_krom_rom_base_one_cell_801/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_589 wl_0_14 sky130_rom_krom_rom_base_one_cell_625/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_578 wl_0_14 sky130_rom_krom_rom_base_one_cell_708/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_567 wl_0_15 sky130_rom_krom_rom_base_one_cell_637/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_556 wl_0_15 sky130_rom_krom_rom_base_one_cell_685/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_545 wl_0_15 sky130_rom_krom_rom_base_one_cell_583/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_534 wl_0_16 sky130_rom_krom_rom_base_one_cell_602/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_523 wl_0_16 sky130_rom_krom_rom_base_one_cell_595/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_512 wl_0_16 sky130_rom_krom_rom_base_one_cell_622/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_501 wl_0_17 sky130_rom_krom_rom_base_one_cell_548/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_14 wl_0_31 sky130_rom_krom_rom_base_one_cell_27/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_25 wl_0_30 sky130_rom_krom_rom_base_one_cell_64/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_36 wl_0_30 sky130_rom_krom_rom_base_one_cell_74/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_47 wl_0_30 sky130_rom_krom_rom_base_one_cell_97/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_58 wl_0_29 sky130_rom_krom_rom_base_zero_cell_58/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_69 wl_0_29 sky130_rom_krom_rom_base_one_cell_26/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_320 wl_0_22 sky130_rom_krom_rom_base_one_cell_420/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_331 wl_0_22 sky130_rom_krom_rom_base_one_cell_429/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_342 wl_0_21 sky130_rom_krom_rom_base_one_cell_411/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_353 wl_0_21 sky130_rom_krom_rom_base_one_cell_418/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_364 wl_0_21 sky130_rom_krom_rom_base_one_cell_429/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_397 wl_0_20 sky130_rom_krom_rom_base_one_cell_602/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_386 wl_0_20 sky130_rom_krom_rom_base_one_cell_477/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_375 wl_0_20 sky130_rom_krom_rom_base_one_cell_587/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_888 wl_0_5 sky130_rom_krom_rom_base_one_cell_888/D
+ sky130_rom_krom_rom_base_one_cell_916/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_877 wl_0_5 sky130_rom_krom_rom_base_one_cell_877/D
+ sky130_rom_krom_rom_base_one_cell_964/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_866 wl_0_6 sky130_rom_krom_rom_base_one_cell_866/D
+ sky130_rom_krom_rom_base_one_cell_898/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_855 wl_0_6 sky130_rom_krom_rom_base_one_cell_855/D
+ sky130_rom_krom_rom_base_one_cell_918/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_844 wl_0_6 sky130_rom_krom_rom_base_one_cell_844/D
+ sky130_rom_krom_rom_base_one_cell_910/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_833 wl_0_7 sky130_rom_krom_rom_base_one_cell_833/D
+ sky130_rom_krom_rom_base_one_cell_925/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_822 wl_0_7 sky130_rom_krom_rom_base_one_cell_822/D
+ sky130_rom_krom_rom_base_one_cell_857/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_811 wl_0_7 sky130_rom_krom_rom_base_one_cell_811/D
+ sky130_rom_krom_rom_base_one_cell_843/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_800 wl_0_7 sky130_rom_krom_rom_base_one_cell_800/D
+ sky130_rom_krom_rom_base_one_cell_834/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_899 wl_0_5 sky130_rom_krom_rom_base_one_cell_899/D
+ sky130_rom_krom_rom_base_one_cell_923/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_107 wl_0_30 sky130_rom_krom_rom_base_one_cell_70/S
+ sky130_rom_krom_rom_base_zero_cell_60/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_118 wl_0_30 sky130_rom_krom_rom_base_one_cell_77/S
+ sky130_rom_krom_rom_base_one_cell_151/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_129 wl_0_30 sky130_rom_krom_rom_base_one_cell_90/S
+ sky130_rom_krom_rom_base_zero_cell_83/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_150 wl_0_26 sky130_rom_krom_rom_base_one_cell_263/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_161 wl_0_26 sky130_rom_krom_rom_base_one_cell_269/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_172 wl_0_26 sky130_rom_krom_rom_base_one_cell_285/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_183 wl_0_26 sky130_rom_krom_rom_base_one_cell_319/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_194 wl_0_25 sky130_rom_krom_rom_base_one_cell_299/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_696 wl_0_11 sky130_rom_krom_rom_base_one_cell_696/D
+ sky130_rom_krom_rom_base_one_cell_730/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_685 wl_0_11 sky130_rom_krom_rom_base_one_cell_685/D
+ sky130_rom_krom_rom_base_one_cell_816/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_674 wl_0_11 sky130_rom_krom_rom_base_one_cell_674/D
+ sky130_rom_krom_rom_base_one_cell_709/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_663 wl_0_12 sky130_rom_krom_rom_base_one_cell_663/D
+ sky130_rom_krom_rom_base_one_cell_692/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_652 wl_0_12 sky130_rom_krom_rom_base_one_cell_652/D
+ sky130_rom_krom_rom_base_one_cell_679/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_641 wl_0_13 sky130_rom_krom_rom_base_one_cell_641/D
+ sky130_rom_krom_rom_base_one_cell_703/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_630 wl_0_13 sky130_rom_krom_rom_base_one_cell_630/D
+ sky130_rom_krom_rom_base_one_cell_660/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_908 wl_0_4 sky130_rom_krom_rom_base_one_cell_942/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_919 wl_0_4 sky130_rom_krom_rom_base_one_cell_980/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_493 wl_0_17 sky130_rom_krom_rom_base_one_cell_493/D
+ sky130_rom_krom_rom_base_one_cell_553/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_482 wl_0_18 sky130_rom_krom_rom_base_one_cell_482/D
+ sky130_rom_krom_rom_base_one_cell_514/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_471 wl_0_18 sky130_rom_krom_rom_base_one_cell_471/D
+ sky130_rom_krom_rom_base_one_cell_535/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_460 wl_0_18 sky130_rom_krom_rom_base_one_cell_460/D
+ sky130_rom_krom_rom_base_one_cell_493/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_290 wl_0_25 sky130_rom_krom_rom_base_one_cell_290/D
+ sky130_rom_krom_rom_base_one_cell_396/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_749 wl_0_9 sky130_rom_krom_rom_base_one_cell_886/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_738 wl_0_9 sky130_rom_krom_rom_base_one_cell_766/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_727 wl_0_10 sky130_rom_krom_rom_base_one_cell_789/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_716 wl_0_10 sky130_rom_krom_rom_base_one_cell_750/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_705 wl_0_10 sky130_rom_krom_rom_base_one_cell_765/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_513 wl_0_16 sky130_rom_krom_rom_base_one_cell_561/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_502 wl_0_17 sky130_rom_krom_rom_base_one_cell_607/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_579 wl_0_14 sky130_rom_krom_rom_base_one_cell_615/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_568 wl_0_15 sky130_rom_krom_rom_base_one_cell_598/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_557 wl_0_15 sky130_rom_krom_rom_base_one_cell_591/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_546 wl_0_15 sky130_rom_krom_rom_base_one_cell_620/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_535 wl_0_16 sky130_rom_krom_rom_base_one_cell_603/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_524 wl_0_16 sky130_rom_krom_rom_base_one_cell_569/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_15 wl_0_31 sky130_rom_krom_rom_base_one_cell_28/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_26 wl_0_30 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_37 wl_0_30 sky130_rom_krom_rom_base_one_cell_75/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_48 wl_0_30 sky130_rom_krom_rom_base_one_cell_55/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_59 wl_0_29 sky130_rom_krom_rom_base_one_cell_69/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_310 wl_0_22 sky130_rom_krom_rom_base_one_cell_412/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_321 wl_0_22 sky130_rom_krom_rom_base_one_cell_391/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_332 wl_0_21 sky130_rom_krom_rom_base_one_cell_522/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_343 wl_0_21 sky130_rom_krom_rom_base_one_cell_470/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_354 wl_0_21 sky130_rom_krom_rom_base_one_cell_630/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_398 wl_0_20 sky130_rom_krom_rom_base_one_cell_603/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_387 wl_0_20 sky130_rom_krom_rom_base_one_cell_478/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_376 wl_0_20 sky130_rom_krom_rom_base_one_cell_468/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_365 wl_0_21 sky130_rom_krom_rom_base_one_cell_431/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_889 wl_0_5 sky130_rom_krom_rom_base_one_cell_889/D
+ sky130_rom_krom_rom_base_one_cell_917/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_878 wl_0_5 sky130_rom_krom_rom_base_one_cell_878/D
+ sky130_rom_krom_rom_base_one_cell_935/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_867 wl_0_6 sky130_rom_krom_rom_base_one_cell_867/D
+ sky130_rom_krom_rom_base_one_cell_867/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_856 wl_0_6 sky130_rom_krom_rom_base_one_cell_856/D
+ sky130_rom_krom_rom_base_one_cell_978/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_845 wl_0_6 sky130_rom_krom_rom_base_one_cell_845/D
+ bl_0_39 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_834 wl_0_6 sky130_rom_krom_rom_base_one_cell_834/D
+ sky130_rom_krom_rom_base_one_cell_872/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_823 wl_0_7 sky130_rom_krom_rom_base_one_cell_823/D
+ sky130_rom_krom_rom_base_one_cell_858/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_812 wl_0_7 sky130_rom_krom_rom_base_one_cell_812/D
+ sky130_rom_krom_rom_base_one_cell_844/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_801 wl_0_7 sky130_rom_krom_rom_base_one_cell_801/D
+ sky130_rom_krom_rom_base_one_cell_903/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_108 wl_0_30 sky130_rom_krom_rom_base_one_cell_71/S
+ sky130_rom_krom_rom_base_zero_cell_61/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_119 wl_0_30 sky130_rom_krom_rom_base_one_cell_81/S
+ sky130_rom_krom_rom_base_zero_cell_74/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_140 wl_0_27 sky130_rom_krom_rom_base_one_cell_286/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_151 wl_0_26 sky130_rom_krom_rom_base_one_cell_373/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_162 wl_0_26 sky130_rom_krom_rom_base_one_cell_301/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_173 wl_0_26 sky130_rom_krom_rom_base_one_cell_286/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_184 wl_0_26 sky130_rom_krom_rom_base_one_cell_344/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_195 wl_0_25 sky130_rom_krom_rom_base_one_cell_323/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_620 wl_0_13 sky130_rom_krom_rom_base_one_cell_620/D
+ sky130_rom_krom_rom_base_one_cell_650/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_697 wl_0_11 sky130_rom_krom_rom_base_one_cell_697/D
+ sky130_rom_krom_rom_base_one_cell_731/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_686 wl_0_11 sky130_rom_krom_rom_base_one_cell_686/D
+ sky130_rom_krom_rom_base_one_cell_723/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_675 wl_0_11 sky130_rom_krom_rom_base_one_cell_675/D
+ sky130_rom_krom_rom_base_one_cell_710/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_664 wl_0_12 sky130_rom_krom_rom_base_one_cell_664/D
+ sky130_rom_krom_rom_base_one_cell_694/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_653 wl_0_12 sky130_rom_krom_rom_base_one_cell_653/D
+ sky130_rom_krom_rom_base_one_cell_718/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_642 wl_0_13 sky130_rom_krom_rom_base_one_cell_642/D
+ sky130_rom_krom_rom_base_one_cell_671/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_631 wl_0_13 sky130_rom_krom_rom_base_one_cell_631/D
+ sky130_rom_krom_rom_base_one_cell_754/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_909 wl_0_4 sky130_rom_krom_rom_base_one_cell_943/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_472 wl_0_18 sky130_rom_krom_rom_base_one_cell_472/D
+ sky130_rom_krom_rom_base_one_cell_502/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_461 wl_0_18 sky130_rom_krom_rom_base_one_cell_461/D
+ sky130_rom_krom_rom_base_one_cell_494/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_450 wl_0_19 sky130_rom_krom_rom_base_one_cell_450/D
+ sky130_rom_krom_rom_base_one_cell_513/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_494 wl_0_17 sky130_rom_krom_rom_base_one_cell_494/D
+ sky130_rom_krom_rom_base_one_cell_525/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_483 wl_0_18 sky130_rom_krom_rom_base_one_cell_483/D
+ sky130_rom_krom_rom_base_one_cell_546/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_280 wl_0_25 sky130_rom_krom_rom_base_one_cell_280/D
+ sky130_rom_krom_rom_base_one_cell_310/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_291 wl_0_25 sky130_rom_krom_rom_base_one_cell_291/D
+ sky130_rom_krom_rom_base_one_cell_398/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_739 wl_0_9 sky130_rom_krom_rom_base_one_cell_769/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_728 wl_0_10 sky130_rom_krom_rom_base_one_cell_792/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_717 wl_0_10 sky130_rom_krom_rom_base_one_cell_816/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_706 wl_0_10 sky130_rom_krom_rom_base_one_cell_738/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_536 wl_0_16 sky130_rom_krom_rom_base_one_cell_604/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_525 wl_0_16 sky130_rom_krom_rom_base_one_cell_570/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_514 wl_0_16 sky130_rom_krom_rom_base_one_cell_626/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_503 wl_0_16 sky130_rom_krom_rom_base_one_cell_549/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_569 wl_0_15 sky130_rom_krom_rom_base_one_cell_601/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_558 wl_0_15 sky130_rom_krom_rom_base_one_cell_628/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_547 wl_0_15 sky130_rom_krom_rom_base_one_cell_587/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_16 wl_0_31 sky130_rom_krom_rom_base_one_cell_29/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_27 wl_0_30 sky130_rom_krom_rom_base_one_cell_65/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_38 wl_0_30 sky130_rom_krom_rom_base_one_cell_26/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_49 wl_0_30 sky130_rom_krom_rom_base_one_cell_57/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_300 wl_0_22 sky130_rom_krom_rom_base_one_cell_377/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_311 wl_0_22 sky130_rom_krom_rom_base_one_cell_443/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_322 wl_0_22 sky130_rom_krom_rom_base_one_cell_423/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_333 wl_0_21 sky130_rom_krom_rom_base_one_cell_403/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_344 wl_0_21 sky130_rom_krom_rom_base_one_cell_412/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_355 wl_0_21 sky130_rom_krom_rom_base_one_cell_419/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_388 wl_0_20 sky130_rom_krom_rom_base_one_cell_630/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_377 wl_0_20 sky130_rom_krom_rom_base_one_cell_442/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_366 wl_0_20 sky130_rom_krom_rom_base_one_cell_491/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_399 wl_0_19 sky130_rom_krom_rom_base_one_cell_491/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_813 wl_0_7 sky130_rom_krom_rom_base_one_cell_813/D
+ sky130_rom_krom_rom_base_one_cell_846/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_802 wl_0_7 sky130_rom_krom_rom_base_one_cell_802/D
+ sky130_rom_krom_rom_base_one_cell_873/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_879 wl_0_5 sky130_rom_krom_rom_base_one_cell_879/D
+ sky130_rom_krom_rom_base_one_cell_936/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_868 wl_0_6 sky130_rom_krom_rom_base_one_cell_868/D
+ sky130_rom_krom_rom_base_one_cell_922/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_857 wl_0_6 sky130_rom_krom_rom_base_one_cell_857/D
+ sky130_rom_krom_rom_base_one_cell_891/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_846 wl_0_6 sky130_rom_krom_rom_base_one_cell_846/D
+ sky130_rom_krom_rom_base_one_cell_885/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_835 wl_0_6 sky130_rom_krom_rom_base_one_cell_835/D
+ sky130_rom_krom_rom_base_one_cell_874/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_824 wl_0_7 sky130_rom_krom_rom_base_one_cell_824/D
+ sky130_rom_krom_rom_base_one_cell_861/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_109 wl_0_30 sky130_rom_krom_rom_base_zero_cell_6/S
+ sky130_rom_krom_rom_base_zero_cell_62/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_130 wl_0_27 sky130_rom_krom_rom_base_one_cell_240/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_141 wl_0_27 sky130_rom_krom_rom_base_zero_cell_83/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_152 wl_0_26 sky130_rom_krom_rom_base_one_cell_294/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_163 wl_0_26 sky130_rom_krom_rom_base_one_cell_271/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_174 wl_0_26 sky130_rom_krom_rom_base_zero_cell_83/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_185 wl_0_25 sky130_rom_krom_rom_base_one_cell_373/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_196 wl_0_25 sky130_rom_krom_rom_base_one_cell_301/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_654 wl_0_12 sky130_rom_krom_rom_base_one_cell_654/D
+ sky130_rom_krom_rom_base_one_cell_721/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_643 wl_0_12 sky130_rom_krom_rom_base_one_cell_643/D
+ sky130_rom_krom_rom_base_one_cell_871/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_632 wl_0_13 sky130_rom_krom_rom_base_one_cell_632/D
+ sky130_rom_krom_rom_base_one_cell_663/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_621 wl_0_13 sky130_rom_krom_rom_base_one_cell_621/D
+ sky130_rom_krom_rom_base_one_cell_676/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_610 wl_0_13 sky130_rom_krom_rom_base_one_cell_610/D
+ sky130_rom_krom_rom_base_one_cell_644/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_698 wl_0_11 sky130_rom_krom_rom_base_one_cell_698/D
+ sky130_rom_krom_rom_base_one_cell_732/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_687 wl_0_11 sky130_rom_krom_rom_base_one_cell_687/D
+ sky130_rom_krom_rom_base_one_cell_888/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_676 wl_0_11 sky130_rom_krom_rom_base_one_cell_676/D
+ sky130_rom_krom_rom_base_one_cell_745/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_665 wl_0_12 sky130_rom_krom_rom_base_one_cell_665/D
+ sky130_rom_krom_rom_base_one_cell_695/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_495 wl_0_17 sky130_rom_krom_rom_base_one_cell_495/D
+ sky130_rom_krom_rom_base_one_cell_554/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_484 wl_0_18 sky130_rom_krom_rom_base_one_cell_484/D
+ sky130_rom_krom_rom_base_one_cell_637/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_473 wl_0_18 sky130_rom_krom_rom_base_one_cell_473/D
+ sky130_rom_krom_rom_base_one_cell_503/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_462 wl_0_18 sky130_rom_krom_rom_base_one_cell_462/D
+ sky130_rom_krom_rom_base_one_cell_495/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_451 wl_0_19 sky130_rom_krom_rom_base_one_cell_451/D
+ sky130_rom_krom_rom_base_one_cell_484/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_440 wl_0_19 sky130_rom_krom_rom_base_one_cell_440/D
+ sky130_rom_krom_rom_base_one_cell_558/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_729 wl_0_10 sky130_rom_krom_rom_base_one_cell_793/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_718 wl_0_10 sky130_rom_krom_rom_base_one_cell_817/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_707 wl_0_10 sky130_rom_krom_rom_base_one_cell_770/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_270 wl_0_25 sky130_rom_krom_rom_base_one_cell_270/D
+ sky130_rom_krom_rom_base_one_cell_302/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_281 wl_0_25 sky130_rom_krom_rom_base_one_cell_281/D
+ sky130_rom_krom_rom_base_one_cell_332/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_292 wl_0_25 sky130_rom_krom_rom_base_one_cell_292/D
+ sky130_rom_krom_rom_base_one_cell_342/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_559 wl_0_15 sky130_rom_krom_rom_base_one_cell_658/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_548 wl_0_15 sky130_rom_krom_rom_base_one_cell_677/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_537 wl_0_16 sky130_rom_krom_rom_base_one_cell_704/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_526 wl_0_16 sky130_rom_krom_rom_base_one_cell_636/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_515 wl_0_16 sky130_rom_krom_rom_base_one_cell_563/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_504 wl_0_16 sky130_rom_krom_rom_base_one_cell_578/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_17 wl_0_31 sky130_rom_krom_rom_base_one_cell_35/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_28 wl_0_30 sky130_rom_krom_rom_base_one_cell_67/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_39 wl_0_30 sky130_rom_krom_rom_base_one_cell_27/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_301 wl_0_22 sky130_rom_krom_rom_base_one_cell_407/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_312 wl_0_22 sky130_rom_krom_rom_base_one_cell_414/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_323 wl_0_22 sky130_rom_krom_rom_base_one_cell_424/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_334 wl_0_21 sky130_rom_krom_rom_base_one_cell_435/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_345 wl_0_21 sky130_rom_krom_rom_base_one_cell_443/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_356 wl_0_21 sky130_rom_krom_rom_base_one_cell_420/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_389 wl_0_20 sky130_rom_krom_rom_base_one_cell_479/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_378 wl_0_20 sky130_rom_krom_rom_base_one_cell_499/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_367 wl_0_20 sky130_rom_krom_rom_base_one_cell_522/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_836 wl_0_6 sky130_rom_krom_rom_base_one_cell_836/D
+ sky130_rom_krom_rom_base_one_cell_876/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_825 wl_0_7 sky130_rom_krom_rom_base_one_cell_825/D
+ sky130_rom_krom_rom_base_one_cell_896/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_814 wl_0_7 sky130_rom_krom_rom_base_one_cell_814/D
+ sky130_rom_krom_rom_base_one_cell_848/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_803 wl_0_7 sky130_rom_krom_rom_base_one_cell_803/D
+ sky130_rom_krom_rom_base_one_cell_962/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_890 wl_0_5 sky130_rom_krom_rom_base_one_cell_925/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_869 wl_0_6 sky130_rom_krom_rom_base_one_cell_869/D
+ sky130_rom_krom_rom_base_one_cell_954/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_858 wl_0_6 sky130_rom_krom_rom_base_one_cell_858/D
+ sky130_rom_krom_rom_base_one_cell_892/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_847 wl_0_6 sky130_rom_krom_rom_base_one_cell_847/D
+ sky130_rom_krom_rom_base_one_cell_913/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_120 wl_0_28 sky130_rom_krom_rom_base_one_cell_57/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_131 wl_0_27 sky130_rom_krom_rom_base_zero_cell_66/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_142 wl_0_27 sky130_rom_krom_rom_base_one_cell_256/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_153 wl_0_26 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_164 wl_0_26 sky130_rom_krom_rom_base_one_cell_273/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_175 wl_0_26 sky130_rom_krom_rom_base_one_cell_316/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_186 wl_0_25 sky130_rom_krom_rom_base_one_cell_294/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_197 wl_0_25 sky130_rom_krom_rom_base_one_cell_304/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_688 wl_0_11 sky130_rom_krom_rom_base_one_cell_688/D
+ sky130_rom_krom_rom_base_one_cell_852/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_677 wl_0_11 sky130_rom_krom_rom_base_one_cell_677/D
+ sky130_rom_krom_rom_base_one_cell_714/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_666 wl_0_12 sky130_rom_krom_rom_base_one_cell_666/D
+ sky130_rom_krom_rom_base_one_cell_789/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_655 wl_0_12 sky130_rom_krom_rom_base_one_cell_655/D
+ sky130_rom_krom_rom_base_one_cell_684/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_644 wl_0_12 sky130_rom_krom_rom_base_one_cell_644/D
+ sky130_rom_krom_rom_base_one_cell_672/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_600 wl_0_14 sky130_rom_krom_rom_base_one_cell_600/D
+ sky130_rom_krom_rom_base_one_cell_733/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_633 wl_0_13 sky130_rom_krom_rom_base_one_cell_633/D
+ sky130_rom_krom_rom_base_one_cell_693/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_622 wl_0_13 sky130_rom_krom_rom_base_one_cell_622/D
+ sky130_rom_krom_rom_base_one_cell_715/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_611 wl_0_13 sky130_rom_krom_rom_base_one_cell_611/D
+ sky130_rom_krom_rom_base_one_cell_765/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_699 wl_0_11 sky130_rom_krom_rom_base_one_cell_699/D
+ sky130_rom_krom_rom_base_one_cell_793/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_496 wl_0_17 sky130_rom_krom_rom_base_one_cell_496/D
+ sky130_rom_krom_rom_base_one_cell_527/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_485 wl_0_18 sky130_rom_krom_rom_base_one_cell_485/D
+ sky130_rom_krom_rom_base_one_cell_516/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_474 wl_0_18 sky130_rom_krom_rom_base_one_cell_474/D
+ sky130_rom_krom_rom_base_one_cell_506/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_463 wl_0_18 sky130_rom_krom_rom_base_one_cell_463/D
+ sky130_rom_krom_rom_base_one_cell_615/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_452 wl_0_19 sky130_rom_krom_rom_base_one_cell_452/D
+ sky130_rom_krom_rom_base_one_cell_487/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_441 wl_0_19 sky130_rom_krom_rom_base_one_cell_441/D
+ sky130_rom_krom_rom_base_one_cell_497/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_430 wl_0_20 sky130_rom_krom_rom_base_one_cell_430/D
+ sky130_rom_krom_rom_base_one_cell_456/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_719 wl_0_10 sky130_rom_krom_rom_base_one_cell_888/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_708 wl_0_10 sky130_rom_krom_rom_base_one_cell_771/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_260 wl_0_26 sky130_rom_krom_rom_base_one_cell_57/S
+ sky130_rom_krom_rom_base_one_cell_292/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_271 wl_0_25 sky130_rom_krom_rom_base_one_cell_271/D
+ sky130_rom_krom_rom_base_one_cell_303/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_282 wl_0_25 sky130_rom_krom_rom_base_one_cell_282/D
+ sky130_rom_krom_rom_base_one_cell_334/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_293 wl_0_25 sky130_rom_krom_rom_base_one_cell_293/D
+ sky130_rom_krom_rom_base_one_cell_367/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_549 wl_0_15 sky130_rom_krom_rom_base_one_cell_622/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_538 wl_0_16 sky130_rom_krom_rom_base_one_cell_607/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_527 wl_0_16 sky130_rom_krom_rom_base_one_cell_637/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_516 wl_0_16 sky130_rom_krom_rom_base_one_cell_655/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_505 wl_0_16 sky130_rom_krom_rom_base_one_cell_553/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_18 wl_0_31 sky130_rom_krom_rom_base_one_cell_37/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_29 wl_0_30 sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_302 wl_0_22 sky130_rom_krom_rom_base_one_cell_438/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_313 wl_0_22 sky130_rom_krom_rom_base_one_cell_386/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_324 wl_0_22 sky130_rom_krom_rom_base_one_cell_425/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_335 wl_0_21 sky130_rom_krom_rom_base_one_cell_406/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_346 wl_0_21 sky130_rom_krom_rom_base_one_cell_414/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_357 wl_0_21 sky130_rom_krom_rom_base_one_cell_422/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_379 wl_0_20 sky130_rom_krom_rom_base_one_cell_470/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_368 wl_0_20 sky130_rom_krom_rom_base_one_cell_492/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_859 wl_0_6 sky130_rom_krom_rom_base_one_cell_859/D
+ sky130_rom_krom_rom_base_one_cell_893/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_848 wl_0_6 sky130_rom_krom_rom_base_one_cell_848/D
+ sky130_rom_krom_rom_base_one_cell_942/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_837 wl_0_6 sky130_rom_krom_rom_base_one_cell_837/D
+ sky130_rom_krom_rom_base_one_cell_906/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_826 wl_0_7 sky130_rom_krom_rom_base_one_cell_826/D
+ sky130_rom_krom_rom_base_one_cell_897/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_815 wl_0_7 sky130_rom_krom_rom_base_one_cell_815/D
+ sky130_rom_krom_rom_base_one_cell_914/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_804 wl_0_7 sky130_rom_krom_rom_base_one_cell_804/D
+ sky130_rom_krom_rom_base_one_cell_963/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_880 wl_0_5 sky130_rom_krom_rom_base_one_cell_919/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_891 wl_0_4 sky130_rom_krom_rom_base_one_cell_927/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_110 wl_0_28 sky130_rom_krom_rom_base_zero_cell_74/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_121 wl_0_28 sky130_rom_krom_rom_base_one_cell_368/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_132 wl_0_27 sky130_rom_krom_rom_base_one_cell_273/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_143 wl_0_27 sky130_rom_krom_rom_base_one_cell_258/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_154 wl_0_26 sky130_rom_krom_rom_base_zero_cell_96/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_165 wl_0_26 sky130_rom_krom_rom_base_one_cell_275/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_176 wl_0_26 sky130_rom_krom_rom_base_one_cell_288/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_187 wl_0_25 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_198 wl_0_25 sky130_rom_krom_rom_base_one_cell_305/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_689 wl_0_11 sky130_rom_krom_rom_base_one_cell_689/D
+ sky130_rom_krom_rom_base_one_cell_784/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_678 wl_0_11 sky130_rom_krom_rom_base_one_cell_678/D
+ sky130_rom_krom_rom_base_one_cell_716/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_667 wl_0_12 sky130_rom_krom_rom_base_one_cell_667/D
+ sky130_rom_krom_rom_base_one_cell_698/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_656 wl_0_12 sky130_rom_krom_rom_base_one_cell_656/D
+ sky130_rom_krom_rom_base_one_cell_686/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_645 wl_0_12 sky130_rom_krom_rom_base_one_cell_645/D
+ sky130_rom_krom_rom_base_one_cell_673/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_601 wl_0_14 sky130_rom_krom_rom_base_one_cell_601/D
+ sky130_rom_krom_rom_base_one_cell_699/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_634 wl_0_13 sky130_rom_krom_rom_base_one_cell_634/D
+ sky130_rom_krom_rom_base_one_cell_729/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_623 wl_0_13 sky130_rom_krom_rom_base_one_cell_623/D
+ sky130_rom_krom_rom_base_one_cell_680/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_612 wl_0_13 sky130_rom_krom_rom_base_one_cell_612/D
+ sky130_rom_krom_rom_base_one_cell_645/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_420 wl_0_20 sky130_rom_krom_rom_base_one_cell_420/D
+ sky130_rom_krom_rom_base_one_cell_481/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_497 wl_0_17 sky130_rom_krom_rom_base_one_cell_497/D
+ sky130_rom_krom_rom_base_one_cell_620/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_486 wl_0_18 sky130_rom_krom_rom_base_one_cell_486/D
+ sky130_rom_krom_rom_base_one_cell_517/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_475 wl_0_18 sky130_rom_krom_rom_base_one_cell_475/D
+ sky130_rom_krom_rom_base_one_cell_508/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_464 wl_0_18 sky130_rom_krom_rom_base_one_cell_464/D
+ sky130_rom_krom_rom_base_one_cell_526/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_453 wl_0_19 sky130_rom_krom_rom_base_one_cell_453/D
+ sky130_rom_krom_rom_base_one_cell_573/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_442 wl_0_19 sky130_rom_krom_rom_base_one_cell_442/D
+ sky130_rom_krom_rom_base_one_cell_469/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_431 wl_0_20 sky130_rom_krom_rom_base_one_cell_431/D
+ sky130_rom_krom_rom_base_one_cell_457/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_250 wl_0_26 sky130_rom_krom_rom_base_zero_cell_74/S
+ sky130_rom_krom_rom_base_one_cell_279/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_261 wl_0_26 sky130_rom_krom_rom_base_one_cell_261/D
+ sky130_rom_krom_rom_base_one_cell_293/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_272 wl_0_25 sky130_rom_krom_rom_base_one_cell_272/D
+ sky130_rom_krom_rom_base_one_cell_325/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_709 wl_0_10 sky130_rom_krom_rom_base_one_cell_807/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_294 wl_0_24 sky130_rom_krom_rom_base_one_cell_294/D
+ sky130_rom_krom_rom_base_one_cell_345/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_283 wl_0_25 sky130_rom_krom_rom_base_one_cell_283/D
+ sky130_rom_krom_rom_base_one_cell_313/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_539 wl_0_15 sky130_rom_krom_rom_base_one_cell_578/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_528 wl_0_16 sky130_rom_krom_rom_base_one_cell_598/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_517 wl_0_16 sky130_rom_krom_rom_base_one_cell_591/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_506 wl_0_16 sky130_rom_krom_rom_base_one_cell_554/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_19 wl_0_31 sky130_rom_krom_rom_base_one_cell_43/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_303 wl_0_22 sky130_rom_krom_rom_base_one_cell_379/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_314 wl_0_22 sky130_rom_krom_rom_base_one_cell_507/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_325 wl_0_22 sky130_rom_krom_rom_base_one_cell_392/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_336 wl_0_21 sky130_rom_krom_rom_base_one_cell_407/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_347 wl_0_21 sky130_rom_krom_rom_base_one_cell_444/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_358 wl_0_21 sky130_rom_krom_rom_base_one_cell_423/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_369 wl_0_20 sky130_rom_krom_rom_base_one_cell_434/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_881 wl_0_5 sky130_rom_krom_rom_base_one_cell_982/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_892 wl_0_4 sky130_rom_krom_rom_base_one_cell_962/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_870 wl_0_5 sky130_rom_krom_rom_base_one_cell_913/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_849 wl_0_6 sky130_rom_krom_rom_base_one_cell_849/D
+ sky130_rom_krom_rom_base_one_cell_943/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_838 wl_0_6 sky130_rom_krom_rom_base_one_cell_838/D
+ sky130_rom_krom_rom_base_one_cell_909/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_827 wl_0_7 sky130_rom_krom_rom_base_one_cell_827/D
+ sky130_rom_krom_rom_base_one_cell_986/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_816 wl_0_7 sky130_rom_krom_rom_base_one_cell_816/D
+ sky130_rom_krom_rom_base_one_cell_849/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_805 wl_0_7 sky130_rom_krom_rom_base_one_cell_805/D
+ sky130_rom_krom_rom_base_one_cell_837/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_100 wl_0_28 sky130_rom_krom_rom_base_one_cell_72/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_111 wl_0_28 sky130_rom_krom_rom_base_one_cell_251/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_122 wl_0_28 sky130_rom_krom_rom_base_one_cell_344/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_133 wl_0_27 sky130_rom_krom_rom_base_one_cell_243/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_144 wl_0_27 sky130_rom_krom_rom_base_one_cell_290/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_155 wl_0_26 sky130_rom_krom_rom_base_one_cell_376/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_166 wl_0_26 sky130_rom_krom_rom_base_one_cell_277/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_177 wl_0_26 sky130_rom_krom_rom_base_one_cell_289/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_188 wl_0_25 sky130_rom_krom_rom_base_one_cell_320/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_199 wl_0_25 sky130_rom_krom_rom_base_one_cell_328/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_602 wl_0_14 sky130_rom_krom_rom_base_one_cell_602/D
+ sky130_rom_krom_rom_base_one_cell_669/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_679 wl_0_11 sky130_rom_krom_rom_base_one_cell_679/D
+ sky130_rom_krom_rom_base_one_cell_717/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_668 wl_0_12 sky130_rom_krom_rom_base_one_cell_668/D
+ sky130_rom_krom_rom_base_one_cell_792/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_657 wl_0_12 sky130_rom_krom_rom_base_one_cell_657/D
+ sky130_rom_krom_rom_base_one_cell_688/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_646 wl_0_12 sky130_rom_krom_rom_base_one_cell_646/D
+ sky130_rom_krom_rom_base_one_cell_770/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_635 wl_0_13 sky130_rom_krom_rom_base_one_cell_635/D
+ sky130_rom_krom_rom_base_one_cell_665/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_624 wl_0_13 sky130_rom_krom_rom_base_one_cell_624/D
+ sky130_rom_krom_rom_base_one_cell_681/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_613 wl_0_13 sky130_rom_krom_rom_base_one_cell_613/D
+ sky130_rom_krom_rom_base_one_cell_707/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_454 wl_0_19 sky130_rom_krom_rom_base_one_cell_454/D
+ sky130_rom_krom_rom_base_one_cell_489/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_443 wl_0_19 sky130_rom_krom_rom_base_one_cell_443/D
+ sky130_rom_krom_rom_base_one_cell_472/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_432 wl_0_20 sky130_rom_krom_rom_base_one_cell_432/D
+ sky130_rom_krom_rom_base_one_cell_458/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_421 wl_0_20 sky130_rom_krom_rom_base_one_cell_421/D
+ sky130_rom_krom_rom_base_one_cell_450/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_410 wl_0_20 sky130_rom_krom_rom_base_one_cell_410/D
+ sky130_rom_krom_rom_base_one_cell_441/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_498 wl_0_17 sky130_rom_krom_rom_base_one_cell_498/D
+ sky130_rom_krom_rom_base_one_cell_532/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_487 wl_0_18 sky130_rom_krom_rom_base_one_cell_487/D
+ sky130_rom_krom_rom_base_one_cell_518/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_476 wl_0_18 sky130_rom_krom_rom_base_one_cell_476/D
+ sky130_rom_krom_rom_base_one_cell_510/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_465 wl_0_18 sky130_rom_krom_rom_base_one_cell_465/D
+ sky130_rom_krom_rom_base_one_cell_496/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_240 wl_0_26 sky130_rom_krom_rom_base_one_cell_240/D
+ sky130_rom_krom_rom_base_one_cell_270/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_251 wl_0_26 sky130_rom_krom_rom_base_one_cell_251/D
+ sky130_rom_krom_rom_base_one_cell_311/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_262 wl_0_26 sky130_rom_krom_rom_base_one_cell_262/D
+ sky130_rom_krom_rom_base_one_cell_343/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_295 wl_0_24 sky130_rom_krom_rom_base_one_cell_295/D
+ sky130_rom_krom_rom_base_one_cell_321/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_273 wl_0_25 sky130_rom_krom_rom_base_one_cell_273/D
+ sky130_rom_krom_rom_base_one_cell_327/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_284 wl_0_25 sky130_rom_krom_rom_base_one_cell_284/D
+ sky130_rom_krom_rom_base_one_cell_314/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_518 wl_0_16 sky130_rom_krom_rom_base_one_cell_564/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_507 wl_0_16 sky130_rom_krom_rom_base_one_cell_615/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_529 wl_0_16 sky130_rom_krom_rom_base_one_cell_571/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_304 wl_0_22 sky130_rom_krom_rom_base_one_cell_381/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_315 wl_0_22 sky130_rom_krom_rom_base_one_cell_475/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_326 wl_0_22 sky130_rom_krom_rom_base_one_cell_393/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_337 wl_0_21 sky130_rom_krom_rom_base_one_cell_438/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_348 wl_0_21 sky130_rom_krom_rom_base_one_cell_507/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_359 wl_0_21 sky130_rom_krom_rom_base_one_cell_424/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_882 wl_0_5 sky130_rom_krom_rom_base_one_cell_984/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_893 wl_0_4 sky130_rom_krom_rom_base_one_cell_995/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_871 wl_0_5 sky130_rom_krom_rom_base_one_cell_942/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_860 wl_0_5 sky130_rom_krom_rom_base_one_cell_905/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_839 wl_0_6 sky130_rom_krom_rom_base_one_cell_839/D
+ sky130_rom_krom_rom_base_one_cell_933/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_828 wl_0_7 sky130_rom_krom_rom_base_one_cell_828/D
+ sky130_rom_krom_rom_base_one_cell_867/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_817 wl_0_7 sky130_rom_krom_rom_base_one_cell_817/D
+ sky130_rom_krom_rom_base_one_cell_850/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_806 wl_0_7 sky130_rom_krom_rom_base_one_cell_806/D
+ sky130_rom_krom_rom_base_one_cell_877/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_101 wl_0_28 sky130_rom_krom_rom_base_zero_cell_65/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_112 wl_0_28 sky130_rom_krom_rom_base_one_cell_281/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_123 wl_0_27 sky130_rom_krom_rom_base_one_cell_294/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_134 wl_0_27 sky130_rom_krom_rom_base_one_cell_80/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_145 wl_0_27 sky130_rom_krom_rom_base_one_cell_57/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_156 wl_0_26 sky130_rom_krom_rom_base_one_cell_297/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_167 wl_0_26 sky130_rom_krom_rom_base_one_cell_80/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_178 wl_0_26 sky130_rom_krom_rom_base_one_cell_290/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_189 wl_0_25 sky130_rom_krom_rom_base_one_cell_376/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_603 wl_0_14 sky130_rom_krom_rom_base_one_cell_603/D
+ sky130_rom_krom_rom_base_one_cell_702/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_636 wl_0_13 sky130_rom_krom_rom_base_one_cell_636/D
+ sky130_rom_krom_rom_base_one_cell_666/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_625 wl_0_13 sky130_rom_krom_rom_base_one_cell_625/D
+ sky130_rom_krom_rom_base_one_cell_653/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_614 wl_0_13 sky130_rom_krom_rom_base_one_cell_614/D
+ sky130_rom_krom_rom_base_one_cell_674/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_690 wl_0_11 sky130_rom_krom_rom_base_one_cell_721/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_669 wl_0_12 sky130_rom_krom_rom_base_one_cell_669/D
+ sky130_rom_krom_rom_base_one_cell_701/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_658 wl_0_12 sky130_rom_krom_rom_base_one_cell_658/D
+ sky130_rom_krom_rom_base_one_cell_753/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_647 wl_0_12 sky130_rom_krom_rom_base_one_cell_647/D
+ sky130_rom_krom_rom_base_one_cell_711/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_400 wl_0_21 sky130_rom_krom_rom_base_one_cell_400/D
+ sky130_rom_krom_rom_base_one_cell_430/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_488 wl_0_18 sky130_rom_krom_rom_base_one_cell_488/D
+ sky130_rom_krom_rom_base_one_cell_519/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_477 wl_0_18 sky130_rom_krom_rom_base_one_cell_477/D
+ sky130_rom_krom_rom_base_one_cell_511/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_466 wl_0_18 sky130_rom_krom_rom_base_one_cell_466/D
+ sky130_rom_krom_rom_base_one_cell_528/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_455 wl_0_19 sky130_rom_krom_rom_base_one_cell_455/D
+ sky130_rom_krom_rom_base_one_cell_604/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_444 wl_0_19 sky130_rom_krom_rom_base_one_cell_444/D
+ sky130_rom_krom_rom_base_one_cell_504/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_433 wl_0_19 sky130_rom_krom_rom_base_one_cell_433/D
+ sky130_rom_krom_rom_base_one_cell_459/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_422 wl_0_20 sky130_rom_krom_rom_base_one_cell_422/D
+ sky130_rom_krom_rom_base_one_cell_482/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_411 wl_0_20 sky130_rom_krom_rom_base_one_cell_411/D
+ sky130_rom_krom_rom_base_one_cell_500/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_499 wl_0_17 sky130_rom_krom_rom_base_one_cell_499/D
+ sky130_rom_krom_rom_base_one_cell_622/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_230 wl_0_27 sky130_rom_krom_rom_base_one_cell_230/D
+ sky130_rom_krom_rom_base_one_cell_341/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_241 wl_0_26 sky130_rom_krom_rom_base_zero_cell_66/S
+ sky130_rom_krom_rom_base_one_cell_272/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_252 wl_0_26 sky130_rom_krom_rom_base_one_cell_252/D
+ sky130_rom_krom_rom_base_one_cell_360/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_263 wl_0_25 sky130_rom_krom_rom_base_one_cell_263/D
+ sky130_rom_krom_rom_base_one_cell_372/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_296 wl_0_24 sky130_rom_krom_rom_base_one_cell_296/D
+ sky130_rom_krom_rom_base_one_cell_347/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_274 wl_0_25 sky130_rom_krom_rom_base_one_cell_274/D
+ sky130_rom_krom_rom_base_one_cell_306/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_285 wl_0_25 sky130_rom_krom_rom_base_one_cell_285/D
+ sky130_rom_krom_rom_base_one_cell_420/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_519 wl_0_16 sky130_rom_krom_rom_base_one_cell_565/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_508 wl_0_16 sky130_rom_krom_rom_base_one_cell_583/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_305 wl_0_22 sky130_rom_krom_rom_base_one_cell_382/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_316 wl_0_22 sky130_rom_krom_rom_base_one_cell_387/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_327 wl_0_22 sky130_rom_krom_rom_base_one_cell_395/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_338 wl_0_21 sky130_rom_krom_rom_base_one_cell_440/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_349 wl_0_21 sky130_rom_krom_rom_base_one_cell_475/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_818 wl_0_7 sky130_rom_krom_rom_base_one_cell_818/D
+ sky130_rom_krom_rom_base_one_cell_851/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_807 wl_0_7 sky130_rom_krom_rom_base_one_cell_807/D
+ sky130_rom_krom_rom_base_one_cell_908/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_883 wl_0_5 sky130_rom_krom_rom_base_one_cell_985/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_894 wl_0_4 sky130_rom_krom_rom_base_one_cell_963/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_872 wl_0_5 sky130_rom_krom_rom_base_one_cell_914/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_861 wl_0_5 sky130_rom_krom_rom_base_one_cell_906/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_850 wl_0_6 sky130_rom_krom_rom_base_one_cell_919/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_829 wl_0_7 sky130_rom_krom_rom_base_one_cell_829/D
+ sky130_rom_krom_rom_base_one_cell_868/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_102 wl_0_28 sky130_rom_krom_rom_base_one_cell_240/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_113 wl_0_28 sky130_rom_krom_rom_base_zero_cell_76/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_124 wl_0_27 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_135 wl_0_27 sky130_rom_krom_rom_base_zero_cell_74/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_146 wl_0_27 sky130_rom_krom_rom_base_one_cell_261/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_157 wl_0_26 sky130_rom_krom_rom_base_one_cell_266/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_168 wl_0_26 sky130_rom_krom_rom_base_one_cell_280/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_179 wl_0_26 sky130_rom_krom_rom_base_one_cell_341/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_659 wl_0_12 sky130_rom_krom_rom_base_one_cell_659/D
+ sky130_rom_krom_rom_base_one_cell_689/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_648 wl_0_12 sky130_rom_krom_rom_base_one_cell_648/D
+ sky130_rom_krom_rom_base_one_cell_773/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_604 wl_0_14 sky130_rom_krom_rom_base_one_cell_604/D
+ sky130_rom_krom_rom_base_one_cell_640/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_637 wl_0_13 sky130_rom_krom_rom_base_one_cell_637/D
+ sky130_rom_krom_rom_base_one_cell_696/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_626 wl_0_13 sky130_rom_krom_rom_base_one_cell_626/D
+ sky130_rom_krom_rom_base_one_cell_682/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_615 wl_0_13 sky130_rom_krom_rom_base_one_cell_615/D
+ sky130_rom_krom_rom_base_one_cell_646/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_691 wl_0_11 sky130_rom_krom_rom_base_one_cell_817/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_680 wl_0_11 sky130_rom_krom_rom_base_one_cell_711/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_489 wl_0_18 sky130_rom_krom_rom_base_one_cell_489/D
+ sky130_rom_krom_rom_base_one_cell_639/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_478 wl_0_18 sky130_rom_krom_rom_base_one_cell_478/D
+ sky130_rom_krom_rom_base_one_cell_658/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_467 wl_0_18 sky130_rom_krom_rom_base_one_cell_467/D
+ sky130_rom_krom_rom_base_one_cell_529/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_456 wl_0_19 sky130_rom_krom_rom_base_one_cell_456/D
+ sky130_rom_krom_rom_base_one_cell_704/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_445 wl_0_19 sky130_rom_krom_rom_base_one_cell_445/D
+ sky130_rom_krom_rom_base_one_cell_505/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_434 wl_0_19 sky130_rom_krom_rom_base_one_cell_434/D
+ sky130_rom_krom_rom_base_one_cell_460/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_423 wl_0_20 sky130_rom_krom_rom_base_one_cell_423/D
+ sky130_rom_krom_rom_base_one_cell_515/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_412 wl_0_20 sky130_rom_krom_rom_base_one_cell_412/D
+ sky130_rom_krom_rom_base_one_cell_471/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_401 wl_0_21 sky130_rom_krom_rom_base_one_cell_401/D
+ sky130_rom_krom_rom_base_one_cell_432/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_990 wl_0_1 sky130_rom_krom_rom_base_one_cell_990/D
+ sky130_rom_krom_rom_base_one_cell_990/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_220 wl_0_27 sky130_rom_krom_rom_base_one_cell_220/D
+ sky130_rom_krom_rom_base_one_cell_253/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_231 wl_0_27 sky130_rom_krom_rom_base_zero_cell_90/S
+ sky130_rom_krom_rom_base_one_cell_291/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_242 wl_0_26 sky130_rom_krom_rom_base_one_cell_242/D
+ sky130_rom_krom_rom_base_one_cell_304/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_253 wl_0_26 sky130_rom_krom_rom_base_one_cell_253/D
+ sky130_rom_krom_rom_base_one_cell_312/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_264 wl_0_25 sky130_rom_krom_rom_base_zero_cell_96/S
+ sky130_rom_krom_rom_base_one_cell_295/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_297 wl_0_24 sky130_rom_krom_rom_base_one_cell_297/D
+ sky130_rom_krom_rom_base_one_cell_322/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_275 wl_0_25 sky130_rom_krom_rom_base_one_cell_275/D
+ sky130_rom_krom_rom_base_one_cell_355/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_286 wl_0_25 sky130_rom_krom_rom_base_one_cell_286/D
+ sky130_rom_krom_rom_base_one_cell_337/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_509 wl_0_16 sky130_rom_krom_rom_base_one_cell_558/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_306 wl_0_22 sky130_rom_krom_rom_base_one_cell_442/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_317 wl_0_22 sky130_rom_krom_rom_base_one_cell_478/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_328 wl_0_22 sky130_rom_krom_rom_base_one_cell_396/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_339 wl_0_21 sky130_rom_krom_rom_base_one_cell_410/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_840 wl_0_6 sky130_rom_krom_rom_base_one_cell_878/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_819 wl_0_7 sky130_rom_krom_rom_base_one_cell_819/D
+ sky130_rom_krom_rom_base_one_cell_854/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_808 wl_0_7 sky130_rom_krom_rom_base_one_cell_808/D
+ sky130_rom_krom_rom_base_one_cell_839/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_884 wl_0_5 sky130_rom_krom_rom_base_one_cell_986/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_895 wl_0_4 bl_0_55 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_873 wl_0_5 sky130_rom_krom_rom_base_one_cell_943/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_862 wl_0_5 sky130_rom_krom_rom_base_one_cell_907/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_851 wl_0_6 sky130_rom_krom_rom_base_one_cell_896/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_103 wl_0_28 sky130_rom_krom_rom_base_zero_cell_66/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_114 wl_0_28 sky130_rom_krom_rom_base_one_cell_286/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_125 wl_0_27 sky130_rom_krom_rom_base_zero_cell_96/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_136 wl_0_27 sky130_rom_krom_rom_base_one_cell_280/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_147 wl_0_27 sky130_rom_krom_rom_base_one_cell_368/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_158 wl_0_26 sky130_rom_krom_rom_base_one_cell_323/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_169 wl_0_26 sky130_rom_krom_rom_base_one_cell_281/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_692 wl_0_11 sky130_rom_krom_rom_base_one_cell_753/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_681 wl_0_11 sky130_rom_krom_rom_base_one_cell_807/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_670 wl_0_12 sky130_rom_krom_rom_base_one_cell_704/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_649 wl_0_12 sky130_rom_krom_rom_base_one_cell_649/D
+ sky130_rom_krom_rom_base_one_cell_743/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_605 wl_0_14 sky130_rom_krom_rom_base_one_cell_605/D
+ sky130_rom_krom_rom_base_one_cell_641/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_638 wl_0_13 sky130_rom_krom_rom_base_one_cell_638/D
+ sky130_rom_krom_rom_base_one_cell_667/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_627 wl_0_13 sky130_rom_krom_rom_base_one_cell_627/D
+ sky130_rom_krom_rom_base_one_cell_817/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_616 wl_0_13 sky130_rom_krom_rom_base_one_cell_616/D
+ sky130_rom_krom_rom_base_one_cell_675/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_402 wl_0_20 sky130_rom_krom_rom_base_one_cell_402/D
+ sky130_rom_krom_rom_base_one_cell_433/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_479 wl_0_18 sky130_rom_krom_rom_base_one_cell_479/D
+ sky130_rom_krom_rom_base_one_cell_542/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_468 wl_0_18 sky130_rom_krom_rom_base_one_cell_468/D
+ sky130_rom_krom_rom_base_one_cell_531/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_457 wl_0_19 sky130_rom_krom_rom_base_one_cell_457/D
+ sky130_rom_krom_rom_base_one_cell_548/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_446 wl_0_19 sky130_rom_krom_rom_base_one_cell_446/D
+ sky130_rom_krom_rom_base_one_cell_509/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_435 wl_0_19 sky130_rom_krom_rom_base_one_cell_435/D
+ sky130_rom_krom_rom_base_one_cell_461/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_424 wl_0_20 sky130_rom_krom_rom_base_one_cell_424/D
+ sky130_rom_krom_rom_base_one_cell_483/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_413 wl_0_20 sky130_rom_krom_rom_base_one_cell_413/D
+ sky130_rom_krom_rom_base_one_cell_473/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_980 wl_0_2 sky130_rom_krom_rom_base_one_cell_980/D
+ sky130_rom_krom_rom_base_one_cell_980/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_991 wl_0_1 sky130_rom_krom_rom_base_one_cell_991/D
+ bl_0_62 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_210 wl_0_27 sky130_rom_krom_rom_base_one_cell_210/D
+ sky130_rom_krom_rom_base_one_cell_242/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_221 wl_0_27 sky130_rom_krom_rom_base_one_cell_221/D
+ sky130_rom_krom_rom_base_one_cell_282/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_232 wl_0_27 sky130_rom_krom_rom_base_one_cell_232/D
+ sky130_rom_krom_rom_base_one_cell_318/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_243 wl_0_26 sky130_rom_krom_rom_base_one_cell_243/D
+ sky130_rom_krom_rom_base_one_cell_305/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_254 wl_0_26 sky130_rom_krom_rom_base_one_cell_254/D
+ sky130_rom_krom_rom_base_one_cell_283/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_265 wl_0_25 sky130_rom_krom_rom_base_one_cell_265/D
+ sky130_rom_krom_rom_base_one_cell_296/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_298 wl_0_24 sky130_rom_krom_rom_base_one_cell_298/D
+ sky130_rom_krom_rom_base_one_cell_349/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_276 wl_0_25 sky130_rom_krom_rom_base_one_cell_276/D
+ sky130_rom_krom_rom_base_one_cell_329/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_287 wl_0_25 sky130_rom_krom_rom_base_one_cell_287/D
+ sky130_rom_krom_rom_base_one_cell_338/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_307 wl_0_22 sky130_rom_krom_rom_base_one_cell_499/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_318 wl_0_22 sky130_rom_krom_rom_base_one_cell_419/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_329 wl_0_22 sky130_rom_krom_rom_base_one_cell_398/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_874 wl_0_5 sky130_rom_krom_rom_base_one_cell_945/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_863 wl_0_5 sky130_rom_krom_rom_base_one_cell_908/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_852 wl_0_6 sky130_rom_krom_rom_base_one_cell_897/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_841 wl_0_6 sky130_rom_krom_rom_base_one_cell_880/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_830 wl_0_6 sky130_rom_krom_rom_base_one_cell_871/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_809 wl_0_7 sky130_rom_krom_rom_base_one_cell_809/D
+ sky130_rom_krom_rom_base_one_cell_840/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_885 wl_0_5 sky130_rom_krom_rom_base_one_cell_921/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_896 wl_0_4 sky130_rom_krom_rom_base_one_cell_964/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_104 wl_0_28 sky130_rom_krom_rom_base_zero_cell_68/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_115 wl_0_28 sky130_rom_krom_rom_base_zero_cell_83/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_126 wl_0_27 sky130_rom_krom_rom_base_one_cell_376/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_137 wl_0_27 sky130_rom_krom_rom_base_one_cell_251/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_148 wl_0_27 sky130_rom_krom_rom_base_one_cell_262/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_159 wl_0_26 sky130_rom_krom_rom_base_one_cell_267/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_693 wl_0_11 sky130_rom_krom_rom_base_one_cell_724/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_682 wl_0_11 sky130_rom_krom_rom_base_one_cell_773/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_671 wl_0_12 sky130_rom_krom_rom_base_one_cell_705/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_660 wl_0_12 sky130_rom_krom_rom_base_one_cell_726/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_606 wl_0_14 sky130_rom_krom_rom_base_one_cell_606/D
+ sky130_rom_krom_rom_base_one_cell_705/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_639 wl_0_13 sky130_rom_krom_rom_base_one_cell_639/D
+ sky130_rom_krom_rom_base_one_cell_700/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_628 wl_0_13 sky130_rom_krom_rom_base_one_cell_628/D
+ sky130_rom_krom_rom_base_one_cell_656/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_617 wl_0_13 sky130_rom_krom_rom_base_one_cell_617/D
+ sky130_rom_krom_rom_base_one_cell_807/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_436 wl_0_19 sky130_rom_krom_rom_base_one_cell_436/D
+ sky130_rom_krom_rom_base_one_cell_464/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_425 wl_0_20 sky130_rom_krom_rom_base_one_cell_425/D
+ sky130_rom_krom_rom_base_one_cell_570/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_414 wl_0_20 sky130_rom_krom_rom_base_one_cell_414/D
+ sky130_rom_krom_rom_base_one_cell_537/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_403 wl_0_20 sky130_rom_krom_rom_base_one_cell_403/D
+ sky130_rom_krom_rom_base_one_cell_523/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_490 wl_0_17 sky130_rom_krom_rom_base_one_cell_544/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_469 wl_0_18 sky130_rom_krom_rom_base_one_cell_469/D
+ sky130_rom_krom_rom_base_one_cell_498/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_458 wl_0_19 sky130_rom_krom_rom_base_one_cell_458/D
+ sky130_rom_krom_rom_base_one_cell_607/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_447 wl_0_19 sky130_rom_krom_rom_base_one_cell_447/D
+ sky130_rom_krom_rom_base_one_cell_476/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_970 wl_0_2 sky130_rom_krom_rom_base_one_cell_970/D
+ bl_0_32 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_981 wl_0_2 sky130_rom_krom_rom_base_one_cell_981/D
+ bl_0_15 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_992 wl_0_1 sky130_rom_krom_rom_base_one_cell_992/D
+ sky130_rom_krom_rom_base_one_cell_992/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_200 wl_0_27 sky130_rom_krom_rom_base_one_cell_7/S
+ sky130_rom_krom_rom_base_one_cell_235/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_211 wl_0_27 sky130_rom_krom_rom_base_zero_cell_68/S
+ sky130_rom_krom_rom_base_one_cell_244/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_222 wl_0_27 sky130_rom_krom_rom_base_one_cell_222/D
+ sky130_rom_krom_rom_base_one_cell_254/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_233 wl_0_27 sky130_rom_krom_rom_base_one_cell_233/D
+ sky130_rom_krom_rom_base_one_cell_319/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_244 wl_0_26 sky130_rom_krom_rom_base_one_cell_244/D
+ sky130_rom_krom_rom_base_one_cell_274/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_255 wl_0_26 sky130_rom_krom_rom_base_one_cell_255/D
+ sky130_rom_krom_rom_base_one_cell_391/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_266 wl_0_25 sky130_rom_krom_rom_base_one_cell_266/D
+ sky130_rom_krom_rom_base_one_cell_379/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_277 wl_0_25 sky130_rom_krom_rom_base_one_cell_277/D
+ sky130_rom_krom_rom_base_one_cell_330/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_299 wl_0_24 sky130_rom_krom_rom_base_one_cell_299/D
+ sky130_rom_krom_rom_base_one_cell_438/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_288 wl_0_25 sky130_rom_krom_rom_base_one_cell_288/D
+ sky130_rom_krom_rom_base_one_cell_395/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_308 wl_0_22 sky130_rom_krom_rom_base_one_cell_411/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_319 wl_0_22 sky130_rom_krom_rom_base_one_cell_390/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_886 wl_0_5 sky130_rom_krom_rom_base_one_cell_867/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_897 wl_0_4 sky130_rom_krom_rom_base_one_cell_933/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_875 wl_0_5 sky130_rom_krom_rom_base_one_cell_853/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_864 wl_0_5 sky130_rom_krom_rom_base_one_cell_909/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_853 wl_0_6 sky130_rom_krom_rom_base_one_cell_986/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_842 wl_0_6 sky130_rom_krom_rom_base_one_cell_883/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_831 wl_0_6 sky130_rom_krom_rom_base_one_cell_903/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_820 wl_0_7 sky130_rom_krom_rom_base_one_cell_948/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_105 wl_0_28 sky130_rom_krom_rom_base_one_cell_26/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_116 wl_0_28 sky130_rom_krom_rom_base_one_cell_258/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_127 wl_0_27 sky130_rom_krom_rom_base_one_cell_69/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_138 wl_0_27 sky130_rom_krom_rom_base_one_cell_281/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_149 wl_0_27 sky130_rom_krom_rom_base_one_cell_344/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_607 wl_0_14 sky130_rom_krom_rom_base_one_cell_607/D
+ sky130_rom_krom_rom_base_one_cell_642/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_618 wl_0_13 sky130_rom_krom_rom_base_one_cell_618/D
+ sky130_rom_krom_rom_base_one_cell_648/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_694 wl_0_11 sky130_rom_krom_rom_base_one_cell_754/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_683 wl_0_11 sky130_rom_krom_rom_base_one_cell_742/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_672 wl_0_11 sky130_rom_krom_rom_base_one_cell_871/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_661 wl_0_12 sky130_rom_krom_rom_base_one_cell_693/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_650 wl_0_12 sky130_rom_krom_rom_base_one_cell_715/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_629 wl_0_13 sky130_rom_krom_rom_base_one_cell_629/D
+ sky130_rom_krom_rom_base_one_cell_687/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_459 wl_0_18 sky130_rom_krom_rom_base_one_cell_459/D
+ sky130_rom_krom_rom_base_one_cell_490/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_448 wl_0_19 sky130_rom_krom_rom_base_one_cell_448/D
+ sky130_rom_krom_rom_base_one_cell_543/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_437 wl_0_19 sky130_rom_krom_rom_base_one_cell_437/D
+ sky130_rom_krom_rom_base_one_cell_465/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_426 wl_0_20 sky130_rom_krom_rom_base_one_cell_426/D
+ sky130_rom_krom_rom_base_one_cell_636/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_415 wl_0_20 sky130_rom_krom_rom_base_one_cell_415/D
+ sky130_rom_krom_rom_base_one_cell_445/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_404 wl_0_20 sky130_rom_krom_rom_base_one_cell_404/D
+ sky130_rom_krom_rom_base_one_cell_524/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_491 wl_0_17 sky130_rom_krom_rom_base_one_cell_546/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_480 wl_0_17 sky130_rom_krom_rom_base_one_cell_587/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_960 wl_0_2 sky130_rom_krom_rom_base_one_cell_960/D
+ sky130_rom_krom_rom_base_one_cell_992/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_971 wl_0_2 sky130_rom_krom_rom_base_one_cell_971/D
+ sky130_rom_krom_rom_base_one_cell_971/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_982 wl_0_2 sky130_rom_krom_rom_base_one_cell_982/D
+ bl_0_13 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_993 wl_0_1 sky130_rom_krom_rom_base_one_cell_993/D
+ sky130_rom_krom_rom_base_one_cell_993/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_201 wl_0_27 sky130_rom_krom_rom_base_one_cell_201/D
+ sky130_rom_krom_rom_base_one_cell_236/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_212 wl_0_27 sky130_rom_krom_rom_base_one_cell_26/S
+ sky130_rom_krom_rom_base_one_cell_245/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_223 wl_0_27 sky130_rom_krom_rom_base_one_cell_223/D
+ sky130_rom_krom_rom_base_one_cell_284/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_234 wl_0_26 sky130_rom_krom_rom_base_one_cell_234/D
+ sky130_rom_krom_rom_base_one_cell_320/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_245 wl_0_26 sky130_rom_krom_rom_base_one_cell_245/D
+ sky130_rom_krom_rom_base_one_cell_328/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_256 wl_0_26 sky130_rom_krom_rom_base_one_cell_256/D
+ sky130_rom_krom_rom_base_one_cell_287/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_267 wl_0_25 sky130_rom_krom_rom_base_one_cell_267/D
+ sky130_rom_krom_rom_base_one_cell_381/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_278 wl_0_25 sky130_rom_krom_rom_base_one_cell_80/S
+ sky130_rom_krom_rom_base_one_cell_387/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_289 wl_0_25 sky130_rom_krom_rom_base_one_cell_289/D
+ sky130_rom_krom_rom_base_one_cell_317/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_790 wl_0_8 sky130_rom_krom_rom_base_one_cell_790/D
+ sky130_rom_krom_rom_base_one_cell_826/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_309 wl_0_22 sky130_rom_krom_rom_base_one_cell_470/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_887 wl_0_5 sky130_rom_krom_rom_base_one_cell_922/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_898 wl_0_4 sky130_rom_krom_rom_base_one_cell_934/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_876 wl_0_5 sky130_rom_krom_rom_base_one_cell_918/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_865 wl_0_5 sky130_rom_krom_rom_base_one_cell_933/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_854 wl_0_6 sky130_rom_krom_rom_base_one_cell_899/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_843 wl_0_6 sky130_rom_krom_rom_base_one_cell_884/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_832 wl_0_6 sky130_rom_krom_rom_base_one_cell_873/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_821 wl_0_7 sky130_rom_krom_rom_base_one_cell_919/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_810 wl_0_7 sky130_rom_krom_rom_base_one_cell_883/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_106 wl_0_28 sky130_rom_krom_rom_base_one_cell_215/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_117 wl_0_28 sky130_rom_krom_rom_base_one_cell_229/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_128 wl_0_27 sky130_rom_krom_rom_base_one_cell_323/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_139 wl_0_27 sky130_rom_krom_rom_base_one_cell_255/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_640 wl_0_12 sky130_rom_krom_rom_base_one_cell_707/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_619 wl_0_13 sky130_rom_krom_rom_base_one_cell_619/D
+ sky130_rom_krom_rom_base_one_cell_649/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_608 wl_0_13 sky130_rom_krom_rom_base_one_cell_608/D
+ sky130_rom_krom_rom_base_one_cell_643/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_695 wl_0_11 sky130_rom_krom_rom_base_one_cell_726/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_684 wl_0_11 sky130_rom_krom_rom_base_one_cell_743/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_673 wl_0_11 sky130_rom_krom_rom_base_one_cell_737/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_662 wl_0_12 sky130_rom_krom_rom_base_one_cell_729/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_651 wl_0_12 sky130_rom_krom_rom_base_one_cell_678/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_481 wl_0_17 sky130_rom_krom_rom_base_one_cell_531/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_470 wl_0_17 sky130_rom_krom_rom_base_one_cell_522/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_449 wl_0_19 sky130_rom_krom_rom_base_one_cell_449/D
+ sky130_rom_krom_rom_base_one_cell_480/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_438 wl_0_19 sky130_rom_krom_rom_base_one_cell_438/D
+ sky130_rom_krom_rom_base_one_cell_583/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_427 wl_0_20 sky130_rom_krom_rom_base_one_cell_427/D
+ sky130_rom_krom_rom_base_one_cell_452/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_416 wl_0_20 sky130_rom_krom_rom_base_one_cell_416/D
+ sky130_rom_krom_rom_base_one_cell_474/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_405 wl_0_20 sky130_rom_krom_rom_base_one_cell_405/D
+ sky130_rom_krom_rom_base_one_cell_462/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_492 wl_0_17 sky130_rom_krom_rom_base_one_cell_570/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_950 wl_0_3 sky130_rom_krom_rom_base_one_cell_950/D
+ bl_0_17 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_961 wl_0_2 sky130_rom_krom_rom_base_one_cell_961/D
+ sky130_rom_krom_rom_base_one_cell_993/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_972 wl_0_2 sky130_rom_krom_rom_base_one_cell_972/D
+ sky130_rom_krom_rom_base_one_cell_972/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_983 wl_0_2 sky130_rom_krom_rom_base_one_cell_983/D
+ sky130_rom_krom_rom_base_one_cell_983/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_994 wl_0_1 sky130_rom_krom_rom_base_one_cell_994/D
+ bl_0_59 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_202 wl_0_27 sky130_rom_krom_rom_base_one_cell_202/D
+ sky130_rom_krom_rom_base_one_cell_237/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_213 wl_0_27 sky130_rom_krom_rom_base_one_cell_213/D
+ sky130_rom_krom_rom_base_one_cell_246/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_224 wl_0_27 sky130_rom_krom_rom_base_one_cell_224/D
+ sky130_rom_krom_rom_base_one_cell_285/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_235 wl_0_26 sky130_rom_krom_rom_base_one_cell_235/D
+ sky130_rom_krom_rom_base_one_cell_265/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_246 wl_0_26 sky130_rom_krom_rom_base_one_cell_246/D
+ sky130_rom_krom_rom_base_one_cell_307/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_257 wl_0_26 sky130_rom_krom_rom_base_one_cell_257/D
+ sky130_rom_krom_rom_base_one_cell_339/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_268 wl_0_25 sky130_rom_krom_rom_base_one_cell_268/D
+ sky130_rom_krom_rom_base_one_cell_351/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_279 wl_0_25 sky130_rom_krom_rom_base_one_cell_279/D
+ sky130_rom_krom_rom_base_one_cell_309/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_90 wl_0_31 sky130_rom_krom_rom_base_one_cell_90/D
+ sky130_rom_krom_rom_base_one_cell_90/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_791 wl_0_8 sky130_rom_krom_rom_base_one_cell_791/D
+ sky130_rom_krom_rom_base_one_cell_863/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_780 wl_0_8 sky130_rom_krom_rom_base_one_cell_780/D
+ sky130_rom_krom_rom_base_one_cell_941/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_822 wl_0_7 sky130_rom_krom_rom_base_one_cell_859/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_811 wl_0_7 sky130_rom_krom_rom_base_one_cell_845/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_800 wl_0_7 sky130_rom_krom_rom_base_one_cell_871/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_888 wl_0_5 sky130_rom_krom_rom_base_one_cell_954/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_899 wl_0_4 sky130_rom_krom_rom_base_one_cell_935/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_877 wl_0_5 sky130_rom_krom_rom_base_one_cell_978/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_866 wl_0_5 sky130_rom_krom_rom_base_one_cell_934/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_855 wl_0_6 sky130_rom_krom_rom_base_one_cell_900/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_844 wl_0_6 sky130_rom_krom_rom_base_one_cell_941/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_833 wl_0_6 sky130_rom_krom_rom_base_one_cell_962/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_107 wl_0_28 sky130_rom_krom_rom_base_one_cell_78/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_118 wl_0_28 sky130_rom_krom_rom_base_one_cell_290/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_129 wl_0_27 sky130_rom_krom_rom_base_one_cell_268/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_674 wl_0_11 sky130_rom_krom_rom_base_one_cell_765/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_663 wl_0_12 sky130_rom_krom_rom_base_one_cell_696/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_652 wl_0_12 sky130_rom_krom_rom_base_one_cell_680/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_641 wl_0_12 sky130_rom_krom_rom_base_one_cell_708/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_630 wl_0_13 sky130_rom_krom_rom_base_one_cell_668/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_609 wl_0_13 sky130_rom_krom_rom_base_one_cell_609/D
+ sky130_rom_krom_rom_base_one_cell_737/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_696 wl_0_11 sky130_rom_krom_rom_base_one_cell_729/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_685 wl_0_11 sky130_rom_krom_rom_base_one_cell_712/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_493 wl_0_17 sky130_rom_krom_rom_base_one_cell_636/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_482 wl_0_17 sky130_rom_krom_rom_base_one_cell_535/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_471 wl_0_17 sky130_rom_krom_rom_base_one_cell_523/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_460 wl_0_18 sky130_rom_krom_rom_base_one_cell_570/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_439 wl_0_19 sky130_rom_krom_rom_base_one_cell_439/D
+ sky130_rom_krom_rom_base_one_cell_467/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_428 wl_0_20 sky130_rom_krom_rom_base_one_cell_428/D
+ sky130_rom_krom_rom_base_one_cell_455/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_417 wl_0_20 sky130_rom_krom_rom_base_one_cell_417/D
+ sky130_rom_krom_rom_base_one_cell_446/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_406 wl_0_20 sky130_rom_krom_rom_base_one_cell_406/D
+ sky130_rom_krom_rom_base_one_cell_463/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_940 wl_0_3 sky130_rom_krom_rom_base_one_cell_940/D
+ bl_0_37 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_951 wl_0_3 sky130_rom_krom_rom_base_one_cell_951/D
+ sky130_rom_krom_rom_base_one_cell_981/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_962 wl_0_2 sky130_rom_krom_rom_base_one_cell_962/D
+ sky130_rom_krom_rom_base_one_cell_994/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_973 wl_0_2 sky130_rom_krom_rom_base_one_cell_973/D
+ sky130_rom_krom_rom_base_one_cell_973/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_984 wl_0_2 sky130_rom_krom_rom_base_one_cell_984/D
+ sky130_rom_krom_rom_base_one_cell_984/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_995 wl_0_1 sky130_rom_krom_rom_base_one_cell_995/D
+ sky130_rom_krom_rom_base_one_cell_995/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_203 wl_0_27 sky130_rom_krom_rom_base_zero_cell_98/S
+ sky130_rom_krom_rom_base_one_cell_297/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_214 wl_0_27 sky130_rom_krom_rom_base_one_cell_214/D
+ sky130_rom_krom_rom_base_one_cell_275/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_225 wl_0_27 sky130_rom_krom_rom_base_one_cell_225/D
+ sky130_rom_krom_rom_base_one_cell_257/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_236 wl_0_26 sky130_rom_krom_rom_base_one_cell_236/D
+ sky130_rom_krom_rom_base_one_cell_377/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_247 wl_0_26 sky130_rom_krom_rom_base_one_cell_247/D
+ sky130_rom_krom_rom_base_one_cell_356/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_258 wl_0_26 sky130_rom_krom_rom_base_one_cell_258/D
+ sky130_rom_krom_rom_base_one_cell_340/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_269 wl_0_25 sky130_rom_krom_rom_base_one_cell_269/D
+ sky130_rom_krom_rom_base_one_cell_300/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_290 wl_0_23 sky130_rom_krom_rom_base_one_cell_398/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_80 wl_0_31 sky130_rom_krom_rom_base_one_cell_80/D
+ sky130_rom_krom_rom_base_one_cell_80/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_91 wl_0_31 sky130_rom_krom_rom_base_one_cell_91/D
+ sky130_rom_krom_rom_base_one_cell_91/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_781 wl_0_8 sky130_rom_krom_rom_base_one_cell_781/D
+ sky130_rom_krom_rom_base_one_cell_847/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_770 wl_0_8 sky130_rom_krom_rom_base_one_cell_770/D
+ sky130_rom_krom_rom_base_one_cell_905/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_792 wl_0_8 sky130_rom_krom_rom_base_one_cell_792/D
+ sky130_rom_krom_rom_base_one_cell_864/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_856 wl_0_6 sky130_rom_krom_rom_base_one_cell_925/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_845 wl_0_6 sky130_rom_krom_rom_base_one_cell_886/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_834 wl_0_6 sky130_rom_krom_rom_base_one_cell_875/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_823 wl_0_7 sky130_rom_krom_rom_base_one_cell_860/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_812 wl_0_7 sky130_rom_krom_rom_base_one_cell_884/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_801 wl_0_7 sky130_rom_krom_rom_base_one_cell_835/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_889 wl_0_5 sky130_rom_krom_rom_base_one_cell_870/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_878 wl_0_5 sky130_rom_krom_rom_base_one_cell_979/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_867 wl_0_5 sky130_rom_krom_rom_base_one_cell_910/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_108 wl_0_28 sky130_rom_krom_rom_base_one_cell_79/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_119 wl_0_28 sky130_rom_krom_rom_base_zero_cell_90/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_697 wl_0_11 sky130_rom_krom_rom_base_one_cell_789/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_686 wl_0_11 sky130_rom_krom_rom_base_one_cell_713/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_675 wl_0_11 sky130_rom_krom_rom_base_one_cell_706/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_664 wl_0_12 sky130_rom_krom_rom_base_one_cell_697/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_653 wl_0_12 sky130_rom_krom_rom_base_one_cell_681/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_642 wl_0_12 sky130_rom_krom_rom_base_one_cell_674/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_631 wl_0_13 sky130_rom_krom_rom_base_one_cell_733/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_620 wl_0_13 sky130_rom_krom_rom_base_one_cell_655/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_418 wl_0_20 sky130_rom_krom_rom_base_one_cell_418/D
+ sky130_rom_krom_rom_base_one_cell_541/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_407 wl_0_20 sky130_rom_krom_rom_base_one_cell_407/D
+ sky130_rom_krom_rom_base_one_cell_436/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_494 wl_0_17 sky130_rom_krom_rom_base_one_cell_637/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_483 wl_0_17 sky130_rom_krom_rom_base_one_cell_537/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_472 wl_0_17 sky130_rom_krom_rom_base_one_cell_524/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_461 wl_0_18 sky130_rom_krom_rom_base_one_cell_636/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_450 wl_0_18 sky130_rom_krom_rom_base_one_cell_504/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_429 wl_0_20 sky130_rom_krom_rom_base_one_cell_429/D
+ sky130_rom_krom_rom_base_one_cell_520/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_930 wl_0_3 sky130_rom_krom_rom_base_one_cell_930/D
+ bl_0_52 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_941 wl_0_3 sky130_rom_krom_rom_base_one_cell_941/D
+ sky130_rom_krom_rom_base_one_cell_968/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_952 wl_0_3 sky130_rom_krom_rom_base_one_cell_952/D
+ sky130_rom_krom_rom_base_one_cell_952/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_963 wl_0_2 sky130_rom_krom_rom_base_one_cell_963/D
+ sky130_rom_krom_rom_base_one_cell_996/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_974 wl_0_2 sky130_rom_krom_rom_base_one_cell_974/D
+ sky130_rom_krom_rom_base_one_cell_974/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_985 wl_0_2 sky130_rom_krom_rom_base_one_cell_985/D
+ sky130_rom_krom_rom_base_one_cell_985/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_996 wl_0_1 sky130_rom_krom_rom_base_one_cell_996/D
+ bl_0_56 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_204 wl_0_27 sky130_rom_krom_rom_base_one_cell_204/D
+ sky130_rom_krom_rom_base_one_cell_239/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_215 wl_0_27 sky130_rom_krom_rom_base_one_cell_215/D
+ sky130_rom_krom_rom_base_one_cell_247/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_226 wl_0_27 sky130_rom_krom_rom_base_one_cell_226/D
+ sky130_rom_krom_rom_base_one_cell_316/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_237 wl_0_26 sky130_rom_krom_rom_base_one_cell_237/D
+ sky130_rom_krom_rom_base_one_cell_348/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_248 wl_0_26 sky130_rom_krom_rom_base_one_cell_248/D
+ sky130_rom_krom_rom_base_one_cell_276/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_259 wl_0_26 sky130_rom_krom_rom_base_one_cell_259/D
+ sky130_rom_krom_rom_base_one_cell_364/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1050 wl_0_0 sky130_rom_krom_rom_base_one_cell_1050/D
+ bl_0_18 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_280 wl_0_23 sky130_rom_krom_rom_base_one_cell_359/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_291 wl_0_23 sky130_rom_krom_rom_base_one_cell_367/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_70 wl_0_31 sky130_rom_krom_rom_base_one_cell_70/D
+ sky130_rom_krom_rom_base_one_cell_70/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_81 wl_0_31 sky130_rom_krom_rom_base_one_cell_81/D
+ sky130_rom_krom_rom_base_one_cell_81/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_92 wl_0_31 sky130_rom_krom_rom_base_one_cell_92/D
+ sky130_rom_krom_rom_base_one_cell_92/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_760 wl_0_9 sky130_rom_krom_rom_base_one_cell_760/D
+ sky130_rom_krom_rom_base_one_cell_828/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_793 wl_0_8 sky130_rom_krom_rom_base_one_cell_793/D
+ sky130_rom_krom_rom_base_one_cell_865/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_782 wl_0_8 sky130_rom_krom_rom_base_one_cell_782/D
+ sky130_rom_krom_rom_base_one_cell_814/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_771 wl_0_8 sky130_rom_krom_rom_base_one_cell_771/D
+ sky130_rom_krom_rom_base_one_cell_805/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_590 wl_0_14 sky130_rom_krom_rom_base_one_cell_590/D
+ sky130_rom_krom_rom_base_one_cell_683/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_879 wl_0_5 sky130_rom_krom_rom_base_one_cell_948/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_868 wl_0_5 bl_0_39 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_857 wl_0_5 sky130_rom_krom_rom_base_one_cell_903/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_846 wl_0_6 sky130_rom_krom_rom_base_one_cell_914/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_835 wl_0_6 sky130_rom_krom_rom_base_one_cell_963/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_824 wl_0_7 sky130_rom_krom_rom_base_one_cell_862/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_813 wl_0_7 sky130_rom_krom_rom_base_one_cell_941/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_802 wl_0_7 sky130_rom_krom_rom_base_one_cell_875/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_109 wl_0_28 sky130_rom_krom_rom_base_one_cell_80/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_698 wl_0_11 sky130_rom_krom_rom_base_one_cell_792/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_687 wl_0_11 sky130_rom_krom_rom_base_one_cell_715/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_676 wl_0_11 sky130_rom_krom_rom_base_one_cell_707/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_665 wl_0_12 sky130_rom_krom_rom_base_one_cell_733/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_654 wl_0_12 sky130_rom_krom_rom_base_one_cell_682/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_643 wl_0_12 sky130_rom_krom_rom_base_one_cell_771/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_632 wl_0_13 sky130_rom_krom_rom_base_one_cell_699/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_621 wl_0_13 sky130_rom_krom_rom_base_one_cell_685/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_610 wl_0_13 sky130_rom_krom_rom_base_one_cell_771/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_419 wl_0_20 sky130_rom_krom_rom_base_one_cell_419/D
+ sky130_rom_krom_rom_base_one_cell_448/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_408 wl_0_20 sky130_rom_krom_rom_base_one_cell_408/D
+ sky130_rom_krom_rom_base_one_cell_439/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_495 wl_0_17 sky130_rom_krom_rom_base_one_cell_573/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_484 wl_0_17 sky130_rom_krom_rom_base_one_cell_591/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_473 wl_0_17 sky130_rom_krom_rom_base_one_cell_615/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_462 wl_0_18 sky130_rom_krom_rom_base_one_cell_573/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_451 wl_0_18 sky130_rom_krom_rom_base_one_cell_505/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_440 wl_0_18 sky130_rom_krom_rom_base_one_cell_523/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_920 wl_0_4 sky130_rom_krom_rom_base_one_cell_920/D
+ sky130_rom_krom_rom_base_one_cell_952/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_931 wl_0_3 sky130_rom_krom_rom_base_one_cell_931/D
+ sky130_rom_krom_rom_base_one_cell_965/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_942 wl_0_3 sky130_rom_krom_rom_base_one_cell_942/D
+ sky130_rom_krom_rom_base_one_cell_942/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_953 wl_0_3 sky130_rom_krom_rom_base_one_cell_953/D
+ sky130_rom_krom_rom_base_one_cell_987/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_964 wl_0_2 sky130_rom_krom_rom_base_one_cell_964/D
+ sky130_rom_krom_rom_base_one_cell_998/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_975 wl_0_2 sky130_rom_krom_rom_base_one_cell_975/D
+ sky130_rom_krom_rom_base_one_cell_975/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_986 wl_0_2 sky130_rom_krom_rom_base_one_cell_986/D
+ sky130_rom_krom_rom_base_one_cell_986/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_997 wl_0_1 sky130_rom_krom_rom_base_one_cell_997/D
+ bl_0_54 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_205 wl_0_27 sky130_rom_krom_rom_base_one_cell_205/D
+ sky130_rom_krom_rom_base_one_cell_266/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_216 wl_0_27 sky130_rom_krom_rom_base_one_cell_216/D
+ sky130_rom_krom_rom_base_one_cell_248/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_227 wl_0_27 sky130_rom_krom_rom_base_one_cell_227/D
+ sky130_rom_krom_rom_base_one_cell_259/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_238 wl_0_26 sky130_rom_krom_rom_base_one_cell_69/S
+ sky130_rom_krom_rom_base_one_cell_298/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_249 wl_0_26 sky130_rom_krom_rom_base_one_cell_249/D
+ sky130_rom_krom_rom_base_one_cell_308/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_270 wl_0_23 sky130_rom_krom_rom_base_one_cell_382/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_281 wl_0_23 sky130_rom_krom_rom_base_one_cell_360/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1051 wl_0_0 sky130_rom_krom_rom_base_one_cell_1051/D
+ bl_0_14 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1040 wl_0_0 sky130_rom_krom_rom_base_one_cell_882/S
+ bl_0_42 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_292 wl_0_23 sky130_rom_krom_rom_base_one_cell_368/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_60 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_60/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_71 wl_0_31 sky130_rom_krom_rom_base_one_cell_71/D
+ sky130_rom_krom_rom_base_one_cell_71/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_82 wl_0_31 sky130_rom_krom_rom_base_one_cell_82/D
+ sky130_rom_krom_rom_base_one_cell_82/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_93 wl_0_31 sky130_rom_krom_rom_base_one_cell_93/D
+ sky130_rom_krom_rom_base_one_cell_93/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_761 wl_0_9 sky130_rom_krom_rom_base_one_cell_761/D
+ sky130_rom_krom_rom_base_one_cell_797/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_794 wl_0_8 sky130_rom_krom_rom_base_one_cell_794/D
+ sky130_rom_krom_rom_base_one_cell_866/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_783 wl_0_8 sky130_rom_krom_rom_base_one_cell_783/D
+ sky130_rom_krom_rom_base_one_cell_818/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_750 wl_0_9 sky130_rom_krom_rom_base_one_cell_750/D
+ sky130_rom_krom_rom_base_one_cell_779/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_772 wl_0_8 sky130_rom_krom_rom_base_one_cell_772/D
+ sky130_rom_krom_rom_base_one_cell_907/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1050 wl_0_0 bl_0_6 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_591 wl_0_14 sky130_rom_krom_rom_base_one_cell_591/D
+ sky130_rom_krom_rom_base_one_cell_627/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_580 wl_0_14 sky130_rom_krom_rom_base_one_cell_580/D
+ sky130_rom_krom_rom_base_one_cell_612/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_869 wl_0_5 sky130_rom_krom_rom_base_one_cell_941/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_858 wl_0_5 sky130_rom_krom_rom_base_one_cell_962/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_847 wl_0_6 sky130_rom_krom_rom_base_one_cell_888/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_836 wl_0_6 sky130_rom_krom_rom_base_one_cell_905/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_825 wl_0_7 sky130_rom_krom_rom_base_one_cell_863/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_814 wl_0_7 sky130_rom_krom_rom_base_one_cell_886/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_803 wl_0_7 sky130_rom_krom_rom_base_one_cell_836/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_600 wl_0_14 sky130_rom_krom_rom_base_one_cell_632/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_622 wl_0_13 sky130_rom_krom_rom_base_one_cell_657/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_611 wl_0_13 sky130_rom_krom_rom_base_one_cell_647/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_699 wl_0_11 sky130_rom_krom_rom_base_one_cell_733/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_688 wl_0_11 sky130_rom_krom_rom_base_one_cell_812/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_677 wl_0_11 sky130_rom_krom_rom_base_one_cell_708/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_666 wl_0_12 sky130_rom_krom_rom_base_one_cell_699/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_655 wl_0_12 sky130_rom_krom_rom_base_one_cell_683/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_644 wl_0_12 sky130_rom_krom_rom_base_one_cell_675/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_633 wl_0_13 sky130_rom_krom_rom_base_one_cell_669/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_463 wl_0_18 sky130_rom_krom_rom_base_one_cell_602/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_452 wl_0_18 sky130_rom_krom_rom_base_one_cell_507/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_441 wl_0_18 sky130_rom_krom_rom_base_one_cell_524/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_430 wl_0_19 sky130_rom_krom_rom_base_one_cell_636/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_409 wl_0_20 sky130_rom_krom_rom_base_one_cell_409/D
+ sky130_rom_krom_rom_base_one_cell_530/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_496 wl_0_17 sky130_rom_krom_rom_base_one_cell_639/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_485 wl_0_17 sky130_rom_krom_rom_base_one_cell_658/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_474 wl_0_17 sky130_rom_krom_rom_base_one_cell_526/D
+ gnd sky130_rom_krom_rom_base_zero_cell
.ends

.subckt sky130_rom_krom_pinv_dec_3 A Z vdd w_692_n79# gnd
X0 vdd A Z w_692_n79# sky130_fd_pr__pfet_01v8 ad=1.5p pd=10.6u as=1.5p ps=10.6u w=5u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.504p pd=3.96u as=0.504p ps=3.96u w=1.68u l=0.15u
.ends

.subckt sky130_rom_krom_rom_bitline_inverter in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7
+ in_8 in_9 in_10 in_11 in_12 in_13 in_14 in_15 in_16 in_17 in_18 in_20 in_21 in_22
+ in_23 in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34 in_35 in_36
+ in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45 in_46 in_47 in_48 in_49 in_50
+ in_51 in_52 in_53 in_54 in_55 in_56 in_57 in_58 in_59 in_60 in_61 in_62 in_63 out_0
+ out_1 out_2 out_3 out_4 out_5 out_6 out_7 out_8 out_9 out_10 out_11 out_12 out_13
+ out_14 out_15 out_16 out_17 out_18 out_20 out_21 out_22 out_23 out_24 out_25 out_26
+ out_27 out_28 out_29 out_30 out_31 out_32 out_33 out_34 out_35 out_36 out_37 out_38
+ out_39 out_40 out_41 out_42 out_43 out_44 out_45 out_46 out_47 out_48 out_49 out_50
+ out_51 out_52 out_53 out_54 out_55 out_56 out_57 out_58 out_59 out_60 out_61 out_62
+ out_63 gnd in_19 sky130_rom_krom_pinv_dec_3_9/w_692_n79# vdd out_19
Xsky130_rom_krom_pinv_dec_3_0 in_0 out_0 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_1 in_1 out_1 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_2 in_2 out_2 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_3 in_3 out_3 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_4 in_4 out_4 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_5 in_5 out_5 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_6 in_6 out_6 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_7 in_7 out_7 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_8 in_8 out_8 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_9 in_9 out_9 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_60 in_60 out_60 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_50 in_50 out_50 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_61 in_61 out_61 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_40 in_40 out_40 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_51 in_51 out_51 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_62 in_62 out_62 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_30 in_30 out_30 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_41 in_41 out_41 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_52 in_52 out_52 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_63 in_63 out_63 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_20 in_20 out_20 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_31 in_31 out_31 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_42 in_42 out_42 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_53 in_53 out_53 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_10 in_10 out_10 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_21 in_21 out_21 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_32 in_32 out_32 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_43 in_43 out_43 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_54 in_54 out_54 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_11 in_11 out_11 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_22 in_22 out_22 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_33 in_33 out_33 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_44 in_44 out_44 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_55 in_55 out_55 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_12 in_12 out_12 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_13 in_13 out_13 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_23 in_23 out_23 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_24 in_24 out_24 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_34 in_34 out_34 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_35 in_35 out_35 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_45 in_45 out_45 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_46 in_46 out_46 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_56 in_56 out_56 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_57 in_57 out_57 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_14 in_14 out_14 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_25 in_25 out_25 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_36 in_36 out_36 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_47 in_47 out_47 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_58 in_58 out_58 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_15 in_15 out_15 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_26 in_26 out_26 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_37 in_37 out_37 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_48 in_48 out_48 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_59 in_59 out_59 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_16 in_16 out_16 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_27 in_27 out_27 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_38 in_38 out_38 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_49 in_49 out_49 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_17 in_17 out_17 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_28 in_28 out_28 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_39 in_39 out_39 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_18 in_18 out_18 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_29 in_29 out_29 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_19 in_19 out_19 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
.ends

.subckt sky130_rom_krom_rom_address_control_array_0 A0_in A1_in A2_in A0_out A1_out
+ A2_out Abar0_out Abar1_out clk vdd vdd_uq0 vdd_uq1 gnd Abar2_out
Xsky130_rom_krom_rom_address_control_buf_0 A2_in A2_out Abar2_out clk vdd vdd_uq0
+ vdd_uq1 gnd sky130_rom_krom_rom_address_control_buf
Xsky130_rom_krom_rom_address_control_buf_2 A0_in A0_out Abar0_out clk vdd vdd_uq0
+ vdd_uq1 gnd sky130_rom_krom_rom_address_control_buf
Xsky130_rom_krom_rom_address_control_buf_1 A1_in A1_out Abar1_out clk vdd vdd_uq0
+ vdd_uq1 gnd sky130_rom_krom_rom_address_control_buf
.ends

.subckt sky130_rom_krom_rom_precharge_array_1 pre_bl0_out pre_bl2_out pre_bl3_out
+ pre_bl6_out pre_bl4_out vdd pre_bl7_out gate pre_bl5_out pre_bl1_out
Xsky130_rom_krom_precharge_cell_2 pre_bl5_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_3 pre_bl4_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_4 pre_bl3_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_5 pre_bl2_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_6 pre_bl1_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_7 pre_bl0_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_0 pre_bl7_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_1 pre_bl6_out gate vdd sky130_rom_krom_precharge_cell
.ends

.subckt sky130_rom_krom_rom_column_decode_array bl_0_0 bl_0_1 bl_0_2 bl_0_3 bl_0_4
+ bl_0_5 bl_0_6 bl_0_7 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 gnd wl_0_0 vdd precharge
Xsky130_rom_krom_rom_base_one_cell_30 wl_0_0 sky130_rom_krom_rom_base_one_cell_30/D
+ bl_0_1 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_20 wl_0_2 sky130_rom_krom_rom_base_one_cell_9/S
+ sky130_rom_krom_rom_base_one_cell_26/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_31 wl_0_0 sky130_rom_krom_rom_base_one_cell_31/D
+ bl_0_0 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_10 wl_0_5 sky130_rom_krom_rom_base_one_cell_4/S
+ sky130_rom_krom_rom_base_zero_cell_6/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_21 wl_0_2 sky130_rom_krom_rom_base_zero_cell_9/S
+ sky130_rom_krom_rom_base_one_cell_27/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_11 wl_0_5 sky130_rom_krom_rom_base_one_cell_6/S
+ sky130_rom_krom_rom_base_zero_cell_7/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_22 wl_0_2 sky130_rom_krom_rom_base_zero_cell_7/S
+ sky130_rom_krom_rom_base_one_cell_30/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_0 precharge gnd sky130_rom_krom_rom_base_one_cell_8/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_12 wl_0_4 sky130_rom_krom_rom_base_one_cell_1/S
+ sky130_rom_krom_rom_base_one_cell_17/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_23 wl_0_2 sky130_rom_krom_rom_base_one_cell_23/D
+ sky130_rom_krom_rom_base_one_cell_31/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1 precharge gnd sky130_rom_krom_rom_base_one_cell_1/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_13 wl_0_4 sky130_rom_krom_rom_base_one_cell_3/S
+ sky130_rom_krom_rom_base_zero_cell_9/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_24 wl_0_1 sky130_rom_krom_rom_base_one_cell_24/D
+ bl_0_7 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_2 precharge gnd sky130_rom_krom_rom_base_one_cell_9/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_0 wl_0_5 sky130_rom_krom_rom_base_one_cell_1/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_14 wl_0_4 sky130_rom_krom_rom_base_one_cell_5/S
+ sky130_rom_krom_rom_base_one_cell_19/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_25 wl_0_1 sky130_rom_krom_rom_base_one_cell_25/D
+ bl_0_6 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_3 precharge gnd sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1 wl_0_5 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_2 wl_0_5 sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_15 wl_0_4 sky130_rom_krom_rom_base_one_cell_7/S
+ sky130_rom_krom_rom_base_one_cell_23/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_26 wl_0_1 sky130_rom_krom_rom_base_one_cell_26/D
+ bl_0_5 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_4 precharge gnd sky130_rom_krom_rom_base_one_cell_4/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_3 wl_0_5 sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_16 wl_0_3 sky130_rom_krom_rom_base_one_cell_8/S
+ sky130_rom_krom_rom_base_one_cell_24/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_17 wl_0_3 sky130_rom_krom_rom_base_one_cell_17/D
+ sky130_rom_krom_rom_base_one_cell_25/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_28 wl_0_0 sky130_rom_krom_rom_base_one_cell_28/D
+ bl_0_3 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_27 wl_0_1 sky130_rom_krom_rom_base_one_cell_27/D
+ bl_0_4 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_5 precharge gnd sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_4 wl_0_4 sky130_rom_krom_rom_base_one_cell_8/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_18 wl_0_3 sky130_rom_krom_rom_base_zero_cell_6/S
+ sky130_rom_krom_rom_base_one_cell_28/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_29 wl_0_0 sky130_rom_krom_rom_base_one_cell_29/D
+ bl_0_2 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_7 precharge gnd sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_6 precharge gnd sky130_rom_krom_rom_base_one_cell_6/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_5 wl_0_4 sky130_rom_krom_rom_base_one_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_19 wl_0_3 sky130_rom_krom_rom_base_one_cell_19/D
+ sky130_rom_krom_rom_base_one_cell_29/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_8 wl_0_5 sky130_rom_krom_rom_base_one_cell_8/D
+ sky130_rom_krom_rom_base_one_cell_8/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_6 wl_0_4 sky130_rom_krom_rom_base_zero_cell_6/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_9 wl_0_5 sky130_rom_krom_rom_base_one_cell_9/D
+ sky130_rom_krom_rom_base_one_cell_9/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_7 wl_0_4 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_20 wl_0_0 bl_0_7 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_8 wl_0_3 sky130_rom_krom_rom_base_one_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_10 wl_0_3 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_21 wl_0_0 bl_0_6 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_9 wl_0_3 sky130_rom_krom_rom_base_zero_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_11 wl_0_3 sky130_rom_krom_rom_base_one_cell_23/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_22 wl_0_0 bl_0_5 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_12 wl_0_2 sky130_rom_krom_rom_base_one_cell_24/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_23 wl_0_0 bl_0_4 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_13 wl_0_2 sky130_rom_krom_rom_base_one_cell_25/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_14 wl_0_2 sky130_rom_krom_rom_base_one_cell_28/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_15 wl_0_2 sky130_rom_krom_rom_base_one_cell_29/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_16 wl_0_1 sky130_rom_krom_rom_base_one_cell_28/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_17 wl_0_1 sky130_rom_krom_rom_base_one_cell_29/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_18 wl_0_1 sky130_rom_krom_rom_base_one_cell_30/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_19 wl_0_1 sky130_rom_krom_rom_base_one_cell_31/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_precharge_array_1_0 bl_0_0 bl_0_2 bl_0_3 bl_0_6 bl_0_4 vdd bl_0_7
+ precharge bl_0_5 bl_0_1 sky130_rom_krom_rom_precharge_array_1
.ends

.subckt sky130_rom_krom_pinv_dec_2 A Z vdd gnd w_504_n45#
X0 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.222p pd=2.08u as=0.222p ps=2.08u w=0.74u l=0.15u
X1 vdd A Z w_504_n45# sky130_fd_pr__pfet_01v8 ad=0.9p pd=6.6u as=0.9p ps=6.6u w=3u l=0.15u
.ends

.subckt sky130_rom_krom_rom_column_decode_wordline_buffer in_0 in_1 in_2 in_3 in_4
+ in_6 in_7 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd in_5
Xsky130_rom_krom_pinv_dec_2_0 in_7 out_7 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_1 in_6 out_6 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_2 in_5 out_5 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_3 in_4 out_4 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_4 in_3 out_3 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_5 in_2 out_2 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_7 in_0 out_0 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_6 in_1 out_1 vdd gnd vdd sky130_rom_krom_pinv_dec_2
.ends

.subckt sky130_rom_krom_rom_column_decode A0 A1 A2 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6
+ wl_7 clk vdd_uq0 vdd_uq1 vdd_uq4 precharge vdd_uq2 vdd gnd
Xsky130_rom_krom_rom_address_control_array_0_0 A0 A1 A2 sky130_rom_krom_rom_column_decode_array_0/wl_0_5
+ sky130_rom_krom_rom_column_decode_array_0/wl_0_3 sky130_rom_krom_rom_column_decode_array_0/wl_0_1
+ sky130_rom_krom_rom_column_decode_array_0/wl_0_4 sky130_rom_krom_rom_column_decode_array_0/wl_0_2
+ clk vdd_uq1 vdd vdd_uq2 gnd sky130_rom_krom_rom_column_decode_array_0/wl_0_0 sky130_rom_krom_rom_address_control_array_0
Xsky130_rom_krom_rom_column_decode_array_0 sky130_rom_krom_rom_column_decode_array_0/bl_0_0
+ sky130_rom_krom_rom_column_decode_array_0/bl_0_1 sky130_rom_krom_rom_column_decode_array_0/bl_0_2
+ sky130_rom_krom_rom_column_decode_array_0/bl_0_3 sky130_rom_krom_rom_column_decode_array_0/bl_0_4
+ sky130_rom_krom_rom_column_decode_array_0/bl_0_5 sky130_rom_krom_rom_column_decode_array_0/bl_0_6
+ sky130_rom_krom_rom_column_decode_array_0/bl_0_7 sky130_rom_krom_rom_column_decode_array_0/wl_0_1
+ sky130_rom_krom_rom_column_decode_array_0/wl_0_2 sky130_rom_krom_rom_column_decode_array_0/wl_0_3
+ sky130_rom_krom_rom_column_decode_array_0/wl_0_4 sky130_rom_krom_rom_column_decode_array_0/wl_0_5
+ gnd sky130_rom_krom_rom_column_decode_array_0/wl_0_0 vdd_uq0 precharge sky130_rom_krom_rom_column_decode_array
Xsky130_rom_krom_rom_column_decode_wordline_buffer_0 sky130_rom_krom_rom_column_decode_array_0/bl_0_0
+ sky130_rom_krom_rom_column_decode_array_0/bl_0_1 sky130_rom_krom_rom_column_decode_array_0/bl_0_2
+ sky130_rom_krom_rom_column_decode_array_0/bl_0_3 sky130_rom_krom_rom_column_decode_array_0/bl_0_4
+ sky130_rom_krom_rom_column_decode_array_0/bl_0_6 sky130_rom_krom_rom_column_decode_array_0/bl_0_7
+ wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 vdd_uq4 gnd sky130_rom_krom_rom_column_decode_array_0/bl_0_5
+ sky130_rom_krom_rom_column_decode_wordline_buffer
.ends

.subckt sky130_rom_krom clk0 cs0 addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5]
+ addr0[6] addr0[7] dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6]
+ dout0[7] vccd1 vssd1
Xsky130_rom_krom_rom_row_decode_0 addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] sky130_rom_krom_rom_row_decode_0/wl_0
+ sky130_rom_krom_rom_row_decode_0/wl_1 sky130_rom_krom_rom_row_decode_0/wl_2 sky130_rom_krom_rom_row_decode_0/wl_3
+ sky130_rom_krom_rom_row_decode_0/wl_4 sky130_rom_krom_rom_row_decode_0/wl_6 sky130_rom_krom_rom_row_decode_0/wl_7
+ sky130_rom_krom_rom_row_decode_0/wl_8 sky130_rom_krom_rom_row_decode_0/wl_9 sky130_rom_krom_rom_row_decode_0/wl_10
+ sky130_rom_krom_rom_row_decode_0/wl_11 sky130_rom_krom_rom_row_decode_0/wl_12 sky130_rom_krom_rom_row_decode_0/wl_13
+ sky130_rom_krom_rom_row_decode_0/wl_14 sky130_rom_krom_rom_row_decode_0/wl_15 sky130_rom_krom_rom_row_decode_0/wl_16
+ sky130_rom_krom_rom_row_decode_0/wl_17 sky130_rom_krom_rom_row_decode_0/wl_18 sky130_rom_krom_rom_row_decode_0/wl_19
+ sky130_rom_krom_rom_row_decode_0/wl_20 sky130_rom_krom_rom_row_decode_0/wl_21 sky130_rom_krom_rom_row_decode_0/wl_22
+ sky130_rom_krom_rom_row_decode_0/wl_23 sky130_rom_krom_rom_row_decode_0/wl_24 sky130_rom_krom_rom_row_decode_0/wl_25
+ sky130_rom_krom_rom_row_decode_0/wl_26 sky130_rom_krom_rom_row_decode_0/wl_27 sky130_rom_krom_rom_row_decode_0/wl_28
+ sky130_rom_krom_rom_row_decode_0/wl_29 sky130_rom_krom_rom_row_decode_0/wl_30 sky130_rom_krom_rom_row_decode_0/wl_31
+ sky130_rom_krom_rom_row_decode_0/clk vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 sky130_rom_krom_rom_row_decode_0/wl_5
+ sky130_rom_krom_rom_row_decode_0/clk vssd1 sky130_rom_krom_rom_row_decode
Xsky130_rom_krom_rom_output_buffer_0 sky130_rom_krom_rom_output_buffer_0/in_0 sky130_rom_krom_rom_output_buffer_0/in_1
+ sky130_rom_krom_rom_output_buffer_0/in_2 sky130_rom_krom_rom_output_buffer_0/in_4
+ sky130_rom_krom_rom_output_buffer_0/in_5 sky130_rom_krom_rom_output_buffer_0/in_6
+ sky130_rom_krom_rom_output_buffer_0/in_7 dout0[0] dout0[1] dout0[2] dout0[3] dout0[4]
+ dout0[5] dout0[6] dout0[7] vssd1 vccd1 sky130_rom_krom_rom_output_buffer_0/in_3
+ sky130_rom_krom_rom_output_buffer
Xsky130_rom_krom_rom_control_logic_0 clk0 cs0 sky130_rom_krom_rom_column_decode_0/clk
+ sky130_rom_krom_rom_row_decode_0/clk vccd1 vssd1 sky130_rom_krom_rom_control_logic
Xsky130_rom_krom_rom_column_mux_array_0 sky130_rom_krom_rom_column_mux_array_0/bl_0
+ sky130_rom_krom_rom_column_mux_array_0/bl_1 sky130_rom_krom_rom_column_mux_array_0/bl_2
+ sky130_rom_krom_rom_column_mux_array_0/bl_3 sky130_rom_krom_rom_column_mux_array_0/bl_4
+ sky130_rom_krom_rom_column_mux_array_0/bl_5 sky130_rom_krom_rom_column_mux_array_0/bl_6
+ sky130_rom_krom_rom_column_mux_array_0/bl_8 sky130_rom_krom_rom_column_mux_array_0/bl_9
+ sky130_rom_krom_rom_column_mux_array_0/bl_11 sky130_rom_krom_rom_column_mux_array_0/bl_15
+ sky130_rom_krom_rom_column_mux_array_0/bl_16 sky130_rom_krom_rom_column_mux_array_0/bl_17
+ sky130_rom_krom_rom_column_mux_array_0/bl_18 sky130_rom_krom_rom_column_mux_array_0/bl_19
+ sky130_rom_krom_rom_column_mux_array_0/bl_22 sky130_rom_krom_rom_column_mux_array_0/bl_26
+ sky130_rom_krom_rom_column_mux_array_0/bl_27 sky130_rom_krom_rom_column_mux_array_0/bl_28
+ sky130_rom_krom_rom_column_mux_array_0/bl_29 sky130_rom_krom_rom_column_mux_array_0/bl_30
+ sky130_rom_krom_rom_column_mux_array_0/bl_37 sky130_rom_krom_rom_column_mux_array_0/bl_38
+ sky130_rom_krom_rom_column_mux_array_0/bl_39 sky130_rom_krom_rom_column_mux_array_0/bl_41
+ sky130_rom_krom_rom_column_mux_array_0/bl_48 sky130_rom_krom_rom_column_mux_array_0/bl_49
+ sky130_rom_krom_rom_column_mux_array_0/bl_52 sky130_rom_krom_rom_column_mux_array_0/bl_59
+ sky130_rom_krom_rom_column_mux_array_0/bl_62 sky130_rom_krom_rom_column_decode_0/wl_3
+ sky130_rom_krom_rom_column_decode_0/wl_4 sky130_rom_krom_rom_column_decode_0/wl_5
+ sky130_rom_krom_rom_output_buffer_0/in_0 sky130_rom_krom_rom_output_buffer_0/in_1
+ sky130_rom_krom_rom_output_buffer_0/in_2 sky130_rom_krom_rom_output_buffer_0/in_3
+ sky130_rom_krom_rom_output_buffer_0/in_4 sky130_rom_krom_rom_output_buffer_0/in_5
+ sky130_rom_krom_rom_output_buffer_0/in_6 sky130_rom_krom_rom_output_buffer_0/in_7
+ vssd1 sky130_rom_krom_rom_column_mux_array_0/bl_24 sky130_rom_krom_rom_column_mux_array_0/bl_35
+ sky130_rom_krom_rom_column_mux_array_0/bl_56 sky130_rom_krom_rom_column_mux_array_0/bl_33
+ sky130_rom_krom_rom_column_mux_array_0/bl_46 sky130_rom_krom_rom_column_mux_array_0/bl_14
+ sky130_rom_krom_rom_column_mux_array_0/bl_12 sky130_rom_krom_rom_column_mux_array_0/bl_25
+ sky130_rom_krom_rom_column_mux_array_0/bl_20 sky130_rom_krom_rom_column_mux_array_0/bl_23
+ sky130_rom_krom_rom_column_mux_array_0/bl_54 sky130_rom_krom_rom_column_mux_array_0/bl_36
+ sky130_rom_krom_rom_column_mux_array_0/bl_31 sky130_rom_krom_rom_column_mux_array_0/bl_44
+ sky130_rom_krom_rom_column_mux_array_0/bl_57 sky130_rom_krom_rom_column_mux_array_0/bl_47
+ sky130_rom_krom_rom_column_mux_array_0/bl_42 sky130_rom_krom_rom_column_mux_array_0/bl_60
+ sky130_rom_krom_rom_column_mux_array_0/bl_50 sky130_rom_krom_rom_column_mux_array_0/bl_63
+ sky130_rom_krom_rom_column_mux_array_0/bl_53 sky130_rom_krom_rom_column_mux_array_0/bl_7
+ sky130_rom_krom_rom_column_mux_array_0/bl_10 sky130_rom_krom_rom_column_mux_array_0/bl_13
+ sky130_rom_krom_rom_column_mux_array_0/bl_21 sky130_rom_krom_rom_column_mux_array_0/bl_34
+ sky130_rom_krom_rom_column_mux_array_0/bl_55 sky130_rom_krom_rom_column_mux_array_0/bl_32
+ sky130_rom_krom_rom_column_mux_array_0/bl_58 sky130_rom_krom_rom_column_mux_array_0/bl_45
+ sky130_rom_krom_rom_column_mux_array_0/bl_40 sky130_rom_krom_rom_column_mux_array_0/bl_43
+ sky130_rom_krom_rom_column_mux_array_0/bl_61 sky130_rom_krom_rom_column_mux_array_0/bl_51
+ sky130_rom_krom_rom_column_decode_0/wl_7 sky130_rom_krom_rom_column_decode_0/wl_0
+ sky130_rom_krom_rom_column_decode_0/wl_6 sky130_rom_krom_rom_column_decode_0/wl_2
+ sky130_rom_krom_rom_column_decode_0/wl_1 sky130_rom_krom_rom_column_mux_array
Xsky130_rom_krom_rom_base_array_0 sky130_rom_krom_rom_base_array_0/bl_0_0 sky130_rom_krom_rom_base_array_0/bl_0_1
+ sky130_rom_krom_rom_base_array_0/bl_0_2 sky130_rom_krom_rom_base_array_0/bl_0_3
+ sky130_rom_krom_rom_base_array_0/bl_0_4 sky130_rom_krom_rom_base_array_0/bl_0_5
+ sky130_rom_krom_rom_base_array_0/bl_0_6 sky130_rom_krom_rom_base_array_0/bl_0_7
+ sky130_rom_krom_rom_base_array_0/bl_0_8 sky130_rom_krom_rom_base_array_0/bl_0_9
+ sky130_rom_krom_rom_base_array_0/bl_0_10 sky130_rom_krom_rom_base_array_0/bl_0_11
+ sky130_rom_krom_rom_base_array_0/bl_0_12 sky130_rom_krom_rom_base_array_0/bl_0_13
+ sky130_rom_krom_rom_base_array_0/bl_0_14 sky130_rom_krom_rom_base_array_0/bl_0_15
+ sky130_rom_krom_rom_base_array_0/bl_0_16 sky130_rom_krom_rom_base_array_0/bl_0_17
+ sky130_rom_krom_rom_base_array_0/bl_0_18 sky130_rom_krom_rom_base_array_0/bl_0_19
+ sky130_rom_krom_rom_base_array_0/bl_0_20 sky130_rom_krom_rom_base_array_0/bl_0_21
+ sky130_rom_krom_rom_base_array_0/bl_0_22 sky130_rom_krom_rom_base_array_0/bl_0_23
+ sky130_rom_krom_rom_base_array_0/bl_0_24 sky130_rom_krom_rom_base_array_0/bl_0_25
+ sky130_rom_krom_rom_base_array_0/bl_0_26 sky130_rom_krom_rom_base_array_0/bl_0_27
+ sky130_rom_krom_rom_base_array_0/bl_0_28 sky130_rom_krom_rom_base_array_0/bl_0_29
+ sky130_rom_krom_rom_base_array_0/bl_0_30 sky130_rom_krom_rom_base_array_0/bl_0_31
+ sky130_rom_krom_rom_base_array_0/bl_0_32 sky130_rom_krom_rom_base_array_0/bl_0_33
+ sky130_rom_krom_rom_base_array_0/bl_0_34 sky130_rom_krom_rom_base_array_0/bl_0_35
+ sky130_rom_krom_rom_base_array_0/bl_0_36 sky130_rom_krom_rom_base_array_0/bl_0_37
+ sky130_rom_krom_rom_base_array_0/bl_0_38 sky130_rom_krom_rom_base_array_0/bl_0_39
+ sky130_rom_krom_rom_base_array_0/bl_0_40 sky130_rom_krom_rom_base_array_0/bl_0_41
+ sky130_rom_krom_rom_base_array_0/bl_0_42 sky130_rom_krom_rom_base_array_0/bl_0_43
+ sky130_rom_krom_rom_base_array_0/bl_0_44 sky130_rom_krom_rom_base_array_0/bl_0_45
+ sky130_rom_krom_rom_base_array_0/bl_0_46 sky130_rom_krom_rom_base_array_0/bl_0_47
+ sky130_rom_krom_rom_base_array_0/bl_0_48 sky130_rom_krom_rom_base_array_0/bl_0_49
+ sky130_rom_krom_rom_base_array_0/bl_0_50 sky130_rom_krom_rom_base_array_0/bl_0_51
+ sky130_rom_krom_rom_base_array_0/bl_0_52 sky130_rom_krom_rom_base_array_0/bl_0_53
+ sky130_rom_krom_rom_base_array_0/bl_0_54 sky130_rom_krom_rom_base_array_0/bl_0_55
+ sky130_rom_krom_rom_base_array_0/bl_0_56 sky130_rom_krom_rom_base_array_0/bl_0_57
+ sky130_rom_krom_rom_base_array_0/bl_0_58 sky130_rom_krom_rom_base_array_0/bl_0_59
+ sky130_rom_krom_rom_base_array_0/bl_0_60 sky130_rom_krom_rom_base_array_0/bl_0_61
+ sky130_rom_krom_rom_base_array_0/bl_0_62 sky130_rom_krom_rom_base_array_0/bl_0_63
+ sky130_rom_krom_rom_row_decode_0/wl_1 sky130_rom_krom_rom_row_decode_0/wl_2 sky130_rom_krom_rom_row_decode_0/wl_3
+ sky130_rom_krom_rom_row_decode_0/wl_4 sky130_rom_krom_rom_row_decode_0/wl_5 sky130_rom_krom_rom_row_decode_0/wl_6
+ sky130_rom_krom_rom_row_decode_0/wl_7 sky130_rom_krom_rom_row_decode_0/wl_8 sky130_rom_krom_rom_row_decode_0/wl_9
+ sky130_rom_krom_rom_row_decode_0/wl_12 sky130_rom_krom_rom_row_decode_0/wl_15 sky130_rom_krom_rom_row_decode_0/wl_16
+ sky130_rom_krom_rom_row_decode_0/wl_17 sky130_rom_krom_rom_row_decode_0/wl_18 sky130_rom_krom_rom_row_decode_0/wl_19
+ sky130_rom_krom_rom_row_decode_0/wl_26 sky130_rom_krom_rom_row_decode_0/wl_27 sky130_rom_krom_rom_row_decode_0/wl_28
+ sky130_rom_krom_rom_row_decode_0/wl_31 vssd1 vssd1 sky130_rom_krom_rom_row_decode_0/wl_13
+ sky130_rom_krom_rom_row_decode_0/wl_22 sky130_rom_krom_rom_row_decode_0/wl_23 sky130_rom_krom_rom_row_decode_0/wl_14
+ sky130_rom_krom_rom_row_decode_0/wl_10 sky130_rom_krom_rom_row_decode_0/wl_24 sky130_rom_krom_rom_row_decode_0/wl_25
+ sky130_rom_krom_rom_row_decode_0/wl_20 sky130_rom_krom_rom_row_decode_0/wl_0 sky130_rom_krom_rom_row_decode_0/wl_21
+ sky130_rom_krom_rom_column_decode_0/clk sky130_rom_krom_rom_row_decode_0/wl_29 sky130_rom_krom_rom_row_decode_0/wl_11
+ sky130_rom_krom_rom_row_decode_0/wl_30 vccd1 sky130_rom_krom_rom_base_array
Xsky130_rom_krom_rom_bitline_inverter_0 sky130_rom_krom_rom_base_array_0/bl_0_0 sky130_rom_krom_rom_base_array_0/bl_0_1
+ sky130_rom_krom_rom_base_array_0/bl_0_2 sky130_rom_krom_rom_base_array_0/bl_0_3
+ sky130_rom_krom_rom_base_array_0/bl_0_4 sky130_rom_krom_rom_base_array_0/bl_0_5
+ sky130_rom_krom_rom_base_array_0/bl_0_6 sky130_rom_krom_rom_base_array_0/bl_0_7
+ sky130_rom_krom_rom_base_array_0/bl_0_8 sky130_rom_krom_rom_base_array_0/bl_0_9
+ sky130_rom_krom_rom_base_array_0/bl_0_10 sky130_rom_krom_rom_base_array_0/bl_0_11
+ sky130_rom_krom_rom_base_array_0/bl_0_12 sky130_rom_krom_rom_base_array_0/bl_0_13
+ sky130_rom_krom_rom_base_array_0/bl_0_14 sky130_rom_krom_rom_base_array_0/bl_0_15
+ sky130_rom_krom_rom_base_array_0/bl_0_16 sky130_rom_krom_rom_base_array_0/bl_0_17
+ sky130_rom_krom_rom_base_array_0/bl_0_18 sky130_rom_krom_rom_base_array_0/bl_0_20
+ sky130_rom_krom_rom_base_array_0/bl_0_21 sky130_rom_krom_rom_base_array_0/bl_0_22
+ sky130_rom_krom_rom_base_array_0/bl_0_23 sky130_rom_krom_rom_base_array_0/bl_0_24
+ sky130_rom_krom_rom_base_array_0/bl_0_25 sky130_rom_krom_rom_base_array_0/bl_0_26
+ sky130_rom_krom_rom_base_array_0/bl_0_27 sky130_rom_krom_rom_base_array_0/bl_0_28
+ sky130_rom_krom_rom_base_array_0/bl_0_29 sky130_rom_krom_rom_base_array_0/bl_0_30
+ sky130_rom_krom_rom_base_array_0/bl_0_31 sky130_rom_krom_rom_base_array_0/bl_0_32
+ sky130_rom_krom_rom_base_array_0/bl_0_33 sky130_rom_krom_rom_base_array_0/bl_0_34
+ sky130_rom_krom_rom_base_array_0/bl_0_35 sky130_rom_krom_rom_base_array_0/bl_0_36
+ sky130_rom_krom_rom_base_array_0/bl_0_37 sky130_rom_krom_rom_base_array_0/bl_0_38
+ sky130_rom_krom_rom_base_array_0/bl_0_39 sky130_rom_krom_rom_base_array_0/bl_0_40
+ sky130_rom_krom_rom_base_array_0/bl_0_41 sky130_rom_krom_rom_base_array_0/bl_0_42
+ sky130_rom_krom_rom_base_array_0/bl_0_43 sky130_rom_krom_rom_base_array_0/bl_0_44
+ sky130_rom_krom_rom_base_array_0/bl_0_45 sky130_rom_krom_rom_base_array_0/bl_0_46
+ sky130_rom_krom_rom_base_array_0/bl_0_47 sky130_rom_krom_rom_base_array_0/bl_0_48
+ sky130_rom_krom_rom_base_array_0/bl_0_49 sky130_rom_krom_rom_base_array_0/bl_0_50
+ sky130_rom_krom_rom_base_array_0/bl_0_51 sky130_rom_krom_rom_base_array_0/bl_0_52
+ sky130_rom_krom_rom_base_array_0/bl_0_53 sky130_rom_krom_rom_base_array_0/bl_0_54
+ sky130_rom_krom_rom_base_array_0/bl_0_55 sky130_rom_krom_rom_base_array_0/bl_0_56
+ sky130_rom_krom_rom_base_array_0/bl_0_57 sky130_rom_krom_rom_base_array_0/bl_0_58
+ sky130_rom_krom_rom_base_array_0/bl_0_59 sky130_rom_krom_rom_base_array_0/bl_0_60
+ sky130_rom_krom_rom_base_array_0/bl_0_61 sky130_rom_krom_rom_base_array_0/bl_0_62
+ sky130_rom_krom_rom_base_array_0/bl_0_63 sky130_rom_krom_rom_column_mux_array_0/bl_0
+ sky130_rom_krom_rom_column_mux_array_0/bl_1 sky130_rom_krom_rom_column_mux_array_0/bl_2
+ sky130_rom_krom_rom_column_mux_array_0/bl_3 sky130_rom_krom_rom_column_mux_array_0/bl_4
+ sky130_rom_krom_rom_column_mux_array_0/bl_5 sky130_rom_krom_rom_column_mux_array_0/bl_6
+ sky130_rom_krom_rom_column_mux_array_0/bl_7 sky130_rom_krom_rom_column_mux_array_0/bl_8
+ sky130_rom_krom_rom_column_mux_array_0/bl_9 sky130_rom_krom_rom_column_mux_array_0/bl_10
+ sky130_rom_krom_rom_column_mux_array_0/bl_11 sky130_rom_krom_rom_column_mux_array_0/bl_12
+ sky130_rom_krom_rom_column_mux_array_0/bl_13 sky130_rom_krom_rom_column_mux_array_0/bl_14
+ sky130_rom_krom_rom_column_mux_array_0/bl_15 sky130_rom_krom_rom_column_mux_array_0/bl_16
+ sky130_rom_krom_rom_column_mux_array_0/bl_17 sky130_rom_krom_rom_column_mux_array_0/bl_18
+ sky130_rom_krom_rom_column_mux_array_0/bl_20 sky130_rom_krom_rom_column_mux_array_0/bl_21
+ sky130_rom_krom_rom_column_mux_array_0/bl_22 sky130_rom_krom_rom_column_mux_array_0/bl_23
+ sky130_rom_krom_rom_column_mux_array_0/bl_24 sky130_rom_krom_rom_column_mux_array_0/bl_25
+ sky130_rom_krom_rom_column_mux_array_0/bl_26 sky130_rom_krom_rom_column_mux_array_0/bl_27
+ sky130_rom_krom_rom_column_mux_array_0/bl_28 sky130_rom_krom_rom_column_mux_array_0/bl_29
+ sky130_rom_krom_rom_column_mux_array_0/bl_30 sky130_rom_krom_rom_column_mux_array_0/bl_31
+ sky130_rom_krom_rom_column_mux_array_0/bl_32 sky130_rom_krom_rom_column_mux_array_0/bl_33
+ sky130_rom_krom_rom_column_mux_array_0/bl_34 sky130_rom_krom_rom_column_mux_array_0/bl_35
+ sky130_rom_krom_rom_column_mux_array_0/bl_36 sky130_rom_krom_rom_column_mux_array_0/bl_37
+ sky130_rom_krom_rom_column_mux_array_0/bl_38 sky130_rom_krom_rom_column_mux_array_0/bl_39
+ sky130_rom_krom_rom_column_mux_array_0/bl_40 sky130_rom_krom_rom_column_mux_array_0/bl_41
+ sky130_rom_krom_rom_column_mux_array_0/bl_42 sky130_rom_krom_rom_column_mux_array_0/bl_43
+ sky130_rom_krom_rom_column_mux_array_0/bl_44 sky130_rom_krom_rom_column_mux_array_0/bl_45
+ sky130_rom_krom_rom_column_mux_array_0/bl_46 sky130_rom_krom_rom_column_mux_array_0/bl_47
+ sky130_rom_krom_rom_column_mux_array_0/bl_48 sky130_rom_krom_rom_column_mux_array_0/bl_49
+ sky130_rom_krom_rom_column_mux_array_0/bl_50 sky130_rom_krom_rom_column_mux_array_0/bl_51
+ sky130_rom_krom_rom_column_mux_array_0/bl_52 sky130_rom_krom_rom_column_mux_array_0/bl_53
+ sky130_rom_krom_rom_column_mux_array_0/bl_54 sky130_rom_krom_rom_column_mux_array_0/bl_55
+ sky130_rom_krom_rom_column_mux_array_0/bl_56 sky130_rom_krom_rom_column_mux_array_0/bl_57
+ sky130_rom_krom_rom_column_mux_array_0/bl_58 sky130_rom_krom_rom_column_mux_array_0/bl_59
+ sky130_rom_krom_rom_column_mux_array_0/bl_60 sky130_rom_krom_rom_column_mux_array_0/bl_61
+ sky130_rom_krom_rom_column_mux_array_0/bl_62 sky130_rom_krom_rom_column_mux_array_0/bl_63
+ vssd1 sky130_rom_krom_rom_base_array_0/bl_0_19 vccd1 vccd1 sky130_rom_krom_rom_column_mux_array_0/bl_19
+ sky130_rom_krom_rom_bitline_inverter
Xsky130_rom_krom_rom_column_decode_0 addr0[0] addr0[1] addr0[2] sky130_rom_krom_rom_column_decode_0/wl_0
+ sky130_rom_krom_rom_column_decode_0/wl_1 sky130_rom_krom_rom_column_decode_0/wl_2
+ sky130_rom_krom_rom_column_decode_0/wl_3 sky130_rom_krom_rom_column_decode_0/wl_4
+ sky130_rom_krom_rom_column_decode_0/wl_5 sky130_rom_krom_rom_column_decode_0/wl_6
+ sky130_rom_krom_rom_column_decode_0/wl_7 sky130_rom_krom_rom_column_decode_0/clk
+ vccd1 vccd1 vccd1 sky130_rom_krom_rom_column_decode_0/clk vccd1 vccd1 vssd1 sky130_rom_krom_rom_column_decode
.ends

