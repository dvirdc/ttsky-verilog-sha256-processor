magic
tech sky130A
magscale 1 2
timestamp 1581320207
<< checkpaint >>
rect -1216 -1310 3060 3819
<< nwell >>
rect 1162 2106 1330 2274
rect 1162 1798 1330 1966
rect 1162 1490 1330 1658
rect 1162 1182 1330 1350
rect 1162 874 1330 1042
rect 1162 566 1330 734
rect 1162 258 1330 426
rect 1162 -50 1330 118
<< pwell >>
rect 263 2139 397 2241
rect 263 1831 397 1933
rect 263 1523 397 1625
rect 263 1215 397 1317
rect 263 907 397 1009
rect 263 599 397 701
rect 263 291 397 393
rect 263 -17 397 85
<< psubdiff >>
rect 289 2207 371 2215
rect 289 2173 313 2207
rect 347 2173 371 2207
rect 289 2165 371 2173
rect 289 1899 371 1907
rect 289 1865 313 1899
rect 347 1865 371 1899
rect 289 1857 371 1865
rect 289 1591 371 1599
rect 289 1557 313 1591
rect 347 1557 371 1591
rect 289 1549 371 1557
rect 289 1283 371 1291
rect 289 1249 313 1283
rect 347 1249 371 1283
rect 289 1241 371 1249
rect 289 975 371 983
rect 289 941 313 975
rect 347 941 371 975
rect 289 933 371 941
rect 289 667 371 675
rect 289 633 313 667
rect 347 633 371 667
rect 289 625 371 633
rect 289 359 371 367
rect 289 325 313 359
rect 347 325 371 359
rect 289 317 371 325
rect 289 51 371 59
rect 289 17 313 51
rect 347 17 371 51
rect 289 9 371 17
<< nsubdiff >>
rect 1205 2207 1287 2215
rect 1205 2173 1229 2207
rect 1263 2173 1287 2207
rect 1205 2165 1287 2173
rect 1205 1899 1287 1907
rect 1205 1865 1229 1899
rect 1263 1865 1287 1899
rect 1205 1857 1287 1865
rect 1205 1591 1287 1599
rect 1205 1557 1229 1591
rect 1263 1557 1287 1591
rect 1205 1549 1287 1557
rect 1205 1283 1287 1291
rect 1205 1249 1229 1283
rect 1263 1249 1287 1283
rect 1205 1241 1287 1249
rect 1205 975 1287 983
rect 1205 941 1229 975
rect 1263 941 1287 975
rect 1205 933 1287 941
rect 1205 667 1287 675
rect 1205 633 1229 667
rect 1263 633 1287 667
rect 1205 625 1287 633
rect 1205 359 1287 367
rect 1205 325 1229 359
rect 1263 325 1287 359
rect 1205 317 1287 325
rect 1205 51 1287 59
rect 1205 17 1229 51
rect 1263 17 1287 51
rect 1205 9 1287 17
<< psubdiffcont >>
rect 313 2173 347 2207
rect 313 1865 347 1899
rect 313 1557 347 1591
rect 313 1249 347 1283
rect 313 941 347 975
rect 313 633 347 667
rect 313 325 347 359
rect 313 17 347 51
<< nsubdiffcont >>
rect 1229 2173 1263 2207
rect 1229 1865 1263 1899
rect 1229 1557 1263 1591
rect 1229 1249 1263 1283
rect 1229 941 1263 975
rect 1229 633 1263 667
rect 1229 325 1263 359
rect 1229 17 1263 51
<< locali >>
rect 60 2311 94 2377
rect 1748 2294 1782 2361
rect 297 2173 313 2207
rect 347 2173 363 2207
rect 1213 2173 1229 2207
rect 1263 2173 1279 2207
rect 60 2003 94 2069
rect 1748 1986 1782 2053
rect 297 1865 313 1899
rect 347 1865 363 1899
rect 1213 1865 1229 1899
rect 1263 1865 1279 1899
rect 60 1695 94 1761
rect 1748 1678 1782 1745
rect 297 1557 313 1591
rect 347 1557 363 1591
rect 1213 1557 1229 1591
rect 1263 1557 1279 1591
rect 60 1387 94 1453
rect 1748 1370 1782 1437
rect 297 1249 313 1283
rect 347 1249 363 1283
rect 1213 1249 1229 1283
rect 1263 1249 1279 1283
rect 60 1079 94 1145
rect 1748 1062 1782 1129
rect 297 941 313 975
rect 347 941 363 975
rect 1213 941 1229 975
rect 1263 941 1279 975
rect 60 771 94 837
rect 1748 754 1782 821
rect 297 633 313 667
rect 347 633 363 667
rect 1213 633 1229 667
rect 1263 633 1279 667
rect 60 463 94 529
rect 1748 446 1782 513
rect 297 325 313 359
rect 347 325 363 359
rect 1213 325 1229 359
rect 1263 325 1279 359
rect 60 155 94 221
rect 1748 138 1782 205
rect 297 17 313 51
rect 347 17 363 51
rect 1213 17 1229 51
rect 1263 17 1279 51
<< viali >>
rect 313 2173 347 2207
rect 1229 2173 1263 2207
rect 313 1865 347 1899
rect 1229 1865 1263 1899
rect 313 1557 347 1591
rect 1229 1557 1263 1591
rect 313 1249 347 1283
rect 1229 1249 1263 1283
rect 313 941 347 975
rect 1229 941 1263 975
rect 313 633 347 667
rect 1229 633 1263 667
rect 313 325 347 359
rect 1229 325 1263 359
rect 313 17 347 51
rect 1229 17 1263 51
<< metal1 >>
rect 316 2219 344 2478
rect 1232 2219 1260 2478
rect 307 2207 353 2219
rect 307 2173 313 2207
rect 347 2173 353 2207
rect 307 2161 353 2173
rect 1223 2207 1269 2219
rect 1223 2173 1229 2207
rect 1263 2173 1269 2207
rect 1223 2161 1269 2173
rect 316 1911 344 2161
rect 1232 1911 1260 2161
rect 307 1899 353 1911
rect 307 1865 313 1899
rect 347 1865 353 1899
rect 307 1853 353 1865
rect 1223 1899 1269 1911
rect 1223 1865 1229 1899
rect 1263 1865 1269 1899
rect 1223 1853 1269 1865
rect 316 1603 344 1853
rect 1232 1603 1260 1853
rect 307 1591 353 1603
rect 307 1557 313 1591
rect 347 1557 353 1591
rect 307 1545 353 1557
rect 1223 1591 1269 1603
rect 1223 1557 1229 1591
rect 1263 1557 1269 1591
rect 1223 1545 1269 1557
rect 316 1295 344 1545
rect 1232 1295 1260 1545
rect 307 1283 353 1295
rect 307 1249 313 1283
rect 347 1249 353 1283
rect 307 1237 353 1249
rect 1223 1283 1269 1295
rect 1223 1249 1229 1283
rect 1263 1249 1269 1283
rect 1223 1237 1269 1249
rect 316 987 344 1237
rect 1232 987 1260 1237
rect 307 975 353 987
rect 307 941 313 975
rect 347 941 353 975
rect 307 929 353 941
rect 1223 975 1269 987
rect 1223 941 1229 975
rect 1263 941 1269 975
rect 1223 929 1269 941
rect 316 679 344 929
rect 1232 679 1260 929
rect 307 667 353 679
rect 307 633 313 667
rect 347 633 353 667
rect 307 621 353 633
rect 1223 667 1269 679
rect 1223 633 1229 667
rect 1263 633 1269 667
rect 1223 621 1269 633
rect 316 371 344 621
rect 1232 371 1260 621
rect 307 359 353 371
rect 307 325 313 359
rect 347 325 353 359
rect 307 313 353 325
rect 1223 359 1269 371
rect 1223 325 1229 359
rect 1263 325 1269 359
rect 1223 313 1269 325
rect 316 63 344 313
rect 1232 63 1260 313
rect 307 51 353 63
rect 307 17 313 51
rect 347 17 353 51
rect 307 5 353 17
rect 1223 51 1269 63
rect 1223 17 1229 51
rect 1263 17 1269 51
rect 1223 5 1269 17
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_0
timestamp 1581320207
transform 1 0 0 0 1 2260
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_1
timestamp 1581320207
transform 1 0 0 0 1 1952
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_2
timestamp 1581320207
transform 1 0 0 0 1 1644
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_3
timestamp 1581320207
transform 1 0 0 0 1 1336
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_4
timestamp 1581320207
transform 1 0 0 0 1 1028
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_5
timestamp 1581320207
transform 1 0 0 0 1 720
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_6
timestamp 1581320207
transform 1 0 0 0 1 412
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_7
timestamp 1581320207
transform 1 0 0 0 1 104
box 44 -50 1800 299
<< labels >>
rlabel locali s 77 188 77 188 4 in_0
port 2 nsew
rlabel locali s 1765 188 1765 188 4 out_0
port 3 nsew
rlabel locali s 77 496 77 496 4 in_1
port 4 nsew
rlabel locali s 1765 496 1765 496 4 out_1
port 5 nsew
rlabel locali s 77 804 77 804 4 in_2
port 6 nsew
rlabel locali s 1765 804 1765 804 4 out_2
port 7 nsew
rlabel locali s 77 1112 77 1112 4 in_3
port 8 nsew
rlabel locali s 1765 1112 1765 1112 4 out_3
port 9 nsew
rlabel locali s 77 1420 77 1420 4 in_4
port 10 nsew
rlabel locali s 1765 1420 1765 1420 4 out_4
port 11 nsew
rlabel locali s 77 1728 77 1728 4 in_5
port 12 nsew
rlabel locali s 1765 1728 1765 1728 4 out_5
port 13 nsew
rlabel locali s 77 2036 77 2036 4 in_6
port 14 nsew
rlabel locali s 1765 2036 1765 2036 4 out_6
port 15 nsew
rlabel locali s 77 2344 77 2344 4 in_7
port 16 nsew
rlabel locali s 1765 2344 1765 2344 4 out_7
port 17 nsew
rlabel metal1 s 316 6 344 34 4 gnd
port 19 nsew
rlabel metal1 s 316 2450 344 2478 4 gnd
port 19 nsew
rlabel metal1 s 1232 2450 1260 2478 4 vdd
port 21 nsew
rlabel metal1 s 1232 6 1260 34 4 vdd
port 21 nsew
<< properties >>
string FIXED_BBOX 1162 -50 1330 0
<< end >>
