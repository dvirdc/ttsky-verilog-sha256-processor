magic
tech sky130A
magscale 1 2
timestamp 1581320205
<< checkpaint >>
rect -1260 -1472 14424 1668
<< nwell >>
rect 0 -196 13164 408
<< poly >>
rect 60 65 90 240
rect 1692 65 1722 240
rect 3324 65 3354 240
rect 4956 65 4986 240
rect 6588 65 6618 240
rect 8220 65 8250 240
rect 9852 65 9882 240
rect 11484 65 11514 240
rect 13116 65 13146 240
rect 60 50 13146 65
rect 61 35 13146 50
<< locali >>
rect 35 -111 69 -95
rect 35 -161 69 -145
rect 239 -111 273 -95
rect 239 -161 273 -145
rect 443 -111 477 -95
rect 443 -161 477 -145
rect 647 -111 681 -95
rect 647 -161 681 -145
rect 851 -111 885 -95
rect 851 -161 885 -145
rect 1055 -111 1089 -95
rect 1055 -161 1089 -145
rect 1259 -111 1293 -95
rect 1259 -161 1293 -145
rect 1463 -111 1497 -95
rect 1463 -161 1497 -145
rect 1667 -111 1701 -95
rect 1667 -161 1701 -145
rect 1871 -111 1905 -95
rect 1871 -161 1905 -145
rect 2075 -111 2109 -95
rect 2075 -161 2109 -145
rect 2279 -111 2313 -95
rect 2279 -161 2313 -145
rect 2483 -111 2517 -95
rect 2483 -161 2517 -145
rect 2687 -111 2721 -95
rect 2687 -161 2721 -145
rect 2891 -111 2925 -95
rect 2891 -161 2925 -145
rect 3095 -111 3129 -95
rect 3095 -161 3129 -145
rect 3299 -111 3333 -95
rect 3299 -161 3333 -145
rect 3503 -111 3537 -95
rect 3503 -161 3537 -145
rect 3707 -111 3741 -95
rect 3707 -161 3741 -145
rect 3911 -111 3945 -95
rect 3911 -161 3945 -145
rect 4115 -111 4149 -95
rect 4115 -161 4149 -145
rect 4319 -111 4353 -95
rect 4319 -161 4353 -145
rect 4523 -111 4557 -95
rect 4523 -161 4557 -145
rect 4727 -111 4761 -95
rect 4727 -161 4761 -145
rect 4931 -111 4965 -95
rect 4931 -161 4965 -145
rect 5135 -111 5169 -95
rect 5135 -161 5169 -145
rect 5339 -111 5373 -95
rect 5339 -161 5373 -145
rect 5543 -111 5577 -95
rect 5543 -161 5577 -145
rect 5747 -111 5781 -95
rect 5747 -161 5781 -145
rect 5951 -111 5985 -95
rect 5951 -161 5985 -145
rect 6155 -111 6189 -95
rect 6155 -161 6189 -145
rect 6359 -111 6393 -95
rect 6359 -161 6393 -145
rect 6563 -111 6597 -95
rect 6563 -161 6597 -145
rect 6767 -111 6801 -95
rect 6767 -161 6801 -145
rect 6971 -111 7005 -95
rect 6971 -161 7005 -145
rect 7175 -111 7209 -95
rect 7175 -161 7209 -145
rect 7379 -111 7413 -95
rect 7379 -161 7413 -145
rect 7583 -111 7617 -95
rect 7583 -161 7617 -145
rect 7787 -111 7821 -95
rect 7787 -161 7821 -145
rect 7991 -111 8025 -95
rect 7991 -161 8025 -145
rect 8195 -111 8229 -95
rect 8195 -161 8229 -145
rect 8399 -111 8433 -95
rect 8399 -161 8433 -145
rect 8603 -111 8637 -95
rect 8603 -161 8637 -145
rect 8807 -111 8841 -95
rect 8807 -161 8841 -145
rect 9011 -111 9045 -95
rect 9011 -161 9045 -145
rect 9215 -111 9249 -95
rect 9215 -161 9249 -145
rect 9419 -111 9453 -95
rect 9419 -161 9453 -145
rect 9623 -111 9657 -95
rect 9623 -161 9657 -145
rect 9827 -111 9861 -95
rect 9827 -161 9861 -145
rect 10031 -111 10065 -95
rect 10031 -161 10065 -145
rect 10235 -111 10269 -95
rect 10235 -161 10269 -145
rect 10439 -111 10473 -95
rect 10439 -161 10473 -145
rect 10643 -111 10677 -95
rect 10643 -161 10677 -145
rect 10847 -111 10881 -95
rect 10847 -161 10881 -145
rect 11051 -111 11085 -95
rect 11051 -161 11085 -145
rect 11255 -111 11289 -95
rect 11255 -161 11289 -145
rect 11459 -111 11493 -95
rect 11459 -161 11493 -145
rect 11663 -111 11697 -95
rect 11663 -161 11697 -145
rect 11867 -111 11901 -95
rect 11867 -161 11901 -145
rect 12071 -111 12105 -95
rect 12071 -161 12105 -145
rect 12275 -111 12309 -95
rect 12275 -161 12309 -145
rect 12479 -111 12513 -95
rect 12479 -161 12513 -145
rect 12683 -111 12717 -95
rect 12683 -161 12717 -145
rect 12887 -111 12921 -95
rect 12887 -161 12921 -145
<< viali >>
rect 35 -145 69 -111
rect 239 -145 273 -111
rect 443 -145 477 -111
rect 647 -145 681 -111
rect 851 -145 885 -111
rect 1055 -145 1089 -111
rect 1259 -145 1293 -111
rect 1463 -145 1497 -111
rect 1667 -145 1701 -111
rect 1871 -145 1905 -111
rect 2075 -145 2109 -111
rect 2279 -145 2313 -111
rect 2483 -145 2517 -111
rect 2687 -145 2721 -111
rect 2891 -145 2925 -111
rect 3095 -145 3129 -111
rect 3299 -145 3333 -111
rect 3503 -145 3537 -111
rect 3707 -145 3741 -111
rect 3911 -145 3945 -111
rect 4115 -145 4149 -111
rect 4319 -145 4353 -111
rect 4523 -145 4557 -111
rect 4727 -145 4761 -111
rect 4931 -145 4965 -111
rect 5135 -145 5169 -111
rect 5339 -145 5373 -111
rect 5543 -145 5577 -111
rect 5747 -145 5781 -111
rect 5951 -145 5985 -111
rect 6155 -145 6189 -111
rect 6359 -145 6393 -111
rect 6563 -145 6597 -111
rect 6767 -145 6801 -111
rect 6971 -145 7005 -111
rect 7175 -145 7209 -111
rect 7379 -145 7413 -111
rect 7583 -145 7617 -111
rect 7787 -145 7821 -111
rect 7991 -145 8025 -111
rect 8195 -145 8229 -111
rect 8399 -145 8433 -111
rect 8603 -145 8637 -111
rect 8807 -145 8841 -111
rect 9011 -145 9045 -111
rect 9215 -145 9249 -111
rect 9419 -145 9453 -111
rect 9623 -145 9657 -111
rect 9827 -145 9861 -111
rect 10031 -145 10065 -111
rect 10235 -145 10269 -111
rect 10439 -145 10473 -111
rect 10643 -145 10677 -111
rect 10847 -145 10881 -111
rect 11051 -145 11085 -111
rect 11255 -145 11289 -111
rect 11459 -145 11493 -111
rect 11663 -145 11697 -111
rect 11867 -145 11901 -111
rect 12071 -145 12105 -111
rect 12275 -145 12309 -111
rect 12479 -145 12513 -111
rect 12683 -145 12717 -111
rect 12887 -145 12921 -111
<< metal1 >>
rect 122 86 150 114
rect 326 86 354 114
rect 530 86 558 114
rect 734 86 762 114
rect 938 86 966 114
rect 1142 86 1170 114
rect 1346 86 1374 114
rect 1550 86 1578 114
rect 1754 86 1782 114
rect 1958 86 1986 114
rect 2162 86 2190 114
rect 2366 86 2394 114
rect 2570 86 2598 114
rect 2774 86 2802 114
rect 2978 86 3006 114
rect 3182 86 3210 114
rect 3386 86 3414 114
rect 3590 86 3618 114
rect 3794 86 3822 114
rect 3998 86 4026 114
rect 4202 86 4230 114
rect 4406 86 4434 114
rect 4610 86 4638 114
rect 4814 86 4842 114
rect 5018 86 5046 114
rect 5222 86 5250 114
rect 5426 86 5454 114
rect 5630 86 5658 114
rect 5834 86 5862 114
rect 6038 86 6066 114
rect 6242 86 6270 114
rect 6446 86 6474 114
rect 6650 86 6678 114
rect 6854 86 6882 114
rect 7058 86 7086 114
rect 7262 86 7290 114
rect 7466 86 7494 114
rect 7670 86 7698 114
rect 7874 86 7902 114
rect 8078 86 8106 114
rect 8282 86 8310 114
rect 8486 86 8514 114
rect 8690 86 8718 114
rect 8894 86 8922 114
rect 9098 86 9126 114
rect 9302 86 9330 114
rect 9506 86 9534 114
rect 9710 86 9738 114
rect 9914 86 9942 114
rect 10118 86 10146 114
rect 10322 86 10350 114
rect 10526 86 10554 114
rect 10730 86 10758 114
rect 10934 86 10962 114
rect 11138 86 11166 114
rect 11342 86 11370 114
rect 11546 86 11574 114
rect 11750 86 11778 114
rect 11954 86 11982 114
rect 12158 86 12186 114
rect 12362 86 12390 114
rect 12566 86 12594 114
rect 12770 86 12798 114
rect 12974 86 13002 114
rect 20 -154 26 -102
rect 78 -154 84 -102
rect 224 -154 230 -102
rect 282 -154 288 -102
rect 428 -154 434 -102
rect 486 -154 492 -102
rect 632 -154 638 -102
rect 690 -154 696 -102
rect 836 -154 842 -102
rect 894 -154 900 -102
rect 1040 -154 1046 -102
rect 1098 -154 1104 -102
rect 1244 -154 1250 -102
rect 1302 -154 1308 -102
rect 1448 -154 1454 -102
rect 1506 -154 1512 -102
rect 1652 -154 1658 -102
rect 1710 -154 1716 -102
rect 1856 -154 1862 -102
rect 1914 -154 1920 -102
rect 2060 -154 2066 -102
rect 2118 -154 2124 -102
rect 2264 -154 2270 -102
rect 2322 -154 2328 -102
rect 2468 -154 2474 -102
rect 2526 -154 2532 -102
rect 2672 -154 2678 -102
rect 2730 -154 2736 -102
rect 2876 -154 2882 -102
rect 2934 -154 2940 -102
rect 3080 -154 3086 -102
rect 3138 -154 3144 -102
rect 3284 -154 3290 -102
rect 3342 -154 3348 -102
rect 3488 -154 3494 -102
rect 3546 -154 3552 -102
rect 3692 -154 3698 -102
rect 3750 -154 3756 -102
rect 3896 -154 3902 -102
rect 3954 -154 3960 -102
rect 4100 -154 4106 -102
rect 4158 -154 4164 -102
rect 4304 -154 4310 -102
rect 4362 -154 4368 -102
rect 4508 -154 4514 -102
rect 4566 -154 4572 -102
rect 4712 -154 4718 -102
rect 4770 -154 4776 -102
rect 4916 -154 4922 -102
rect 4974 -154 4980 -102
rect 5120 -154 5126 -102
rect 5178 -154 5184 -102
rect 5324 -154 5330 -102
rect 5382 -154 5388 -102
rect 5528 -154 5534 -102
rect 5586 -154 5592 -102
rect 5732 -154 5738 -102
rect 5790 -154 5796 -102
rect 5936 -154 5942 -102
rect 5994 -154 6000 -102
rect 6140 -154 6146 -102
rect 6198 -154 6204 -102
rect 6344 -154 6350 -102
rect 6402 -154 6408 -102
rect 6548 -154 6554 -102
rect 6606 -154 6612 -102
rect 6752 -154 6758 -102
rect 6810 -154 6816 -102
rect 6956 -154 6962 -102
rect 7014 -154 7020 -102
rect 7160 -154 7166 -102
rect 7218 -154 7224 -102
rect 7364 -154 7370 -102
rect 7422 -154 7428 -102
rect 7568 -154 7574 -102
rect 7626 -154 7632 -102
rect 7772 -154 7778 -102
rect 7830 -154 7836 -102
rect 7976 -154 7982 -102
rect 8034 -154 8040 -102
rect 8180 -154 8186 -102
rect 8238 -154 8244 -102
rect 8384 -154 8390 -102
rect 8442 -154 8448 -102
rect 8588 -154 8594 -102
rect 8646 -154 8652 -102
rect 8792 -154 8798 -102
rect 8850 -154 8856 -102
rect 8996 -154 9002 -102
rect 9054 -154 9060 -102
rect 9200 -154 9206 -102
rect 9258 -154 9264 -102
rect 9404 -154 9410 -102
rect 9462 -154 9468 -102
rect 9608 -154 9614 -102
rect 9666 -154 9672 -102
rect 9812 -154 9818 -102
rect 9870 -154 9876 -102
rect 10016 -154 10022 -102
rect 10074 -154 10080 -102
rect 10220 -154 10226 -102
rect 10278 -154 10284 -102
rect 10424 -154 10430 -102
rect 10482 -154 10488 -102
rect 10628 -154 10634 -102
rect 10686 -154 10692 -102
rect 10832 -154 10838 -102
rect 10890 -154 10896 -102
rect 11036 -154 11042 -102
rect 11094 -154 11100 -102
rect 11240 -154 11246 -102
rect 11298 -154 11304 -102
rect 11444 -154 11450 -102
rect 11502 -154 11508 -102
rect 11648 -154 11654 -102
rect 11706 -154 11712 -102
rect 11852 -154 11858 -102
rect 11910 -154 11916 -102
rect 12056 -154 12062 -102
rect 12114 -154 12120 -102
rect 12260 -154 12266 -102
rect 12318 -154 12324 -102
rect 12464 -154 12470 -102
rect 12522 -154 12528 -102
rect 12668 -154 12674 -102
rect 12726 -154 12732 -102
rect 12872 -154 12878 -102
rect 12930 -154 12936 -102
<< via1 >>
rect 26 -111 78 -102
rect 26 -145 35 -111
rect 35 -145 69 -111
rect 69 -145 78 -111
rect 26 -154 78 -145
rect 230 -111 282 -102
rect 230 -145 239 -111
rect 239 -145 273 -111
rect 273 -145 282 -111
rect 230 -154 282 -145
rect 434 -111 486 -102
rect 434 -145 443 -111
rect 443 -145 477 -111
rect 477 -145 486 -111
rect 434 -154 486 -145
rect 638 -111 690 -102
rect 638 -145 647 -111
rect 647 -145 681 -111
rect 681 -145 690 -111
rect 638 -154 690 -145
rect 842 -111 894 -102
rect 842 -145 851 -111
rect 851 -145 885 -111
rect 885 -145 894 -111
rect 842 -154 894 -145
rect 1046 -111 1098 -102
rect 1046 -145 1055 -111
rect 1055 -145 1089 -111
rect 1089 -145 1098 -111
rect 1046 -154 1098 -145
rect 1250 -111 1302 -102
rect 1250 -145 1259 -111
rect 1259 -145 1293 -111
rect 1293 -145 1302 -111
rect 1250 -154 1302 -145
rect 1454 -111 1506 -102
rect 1454 -145 1463 -111
rect 1463 -145 1497 -111
rect 1497 -145 1506 -111
rect 1454 -154 1506 -145
rect 1658 -111 1710 -102
rect 1658 -145 1667 -111
rect 1667 -145 1701 -111
rect 1701 -145 1710 -111
rect 1658 -154 1710 -145
rect 1862 -111 1914 -102
rect 1862 -145 1871 -111
rect 1871 -145 1905 -111
rect 1905 -145 1914 -111
rect 1862 -154 1914 -145
rect 2066 -111 2118 -102
rect 2066 -145 2075 -111
rect 2075 -145 2109 -111
rect 2109 -145 2118 -111
rect 2066 -154 2118 -145
rect 2270 -111 2322 -102
rect 2270 -145 2279 -111
rect 2279 -145 2313 -111
rect 2313 -145 2322 -111
rect 2270 -154 2322 -145
rect 2474 -111 2526 -102
rect 2474 -145 2483 -111
rect 2483 -145 2517 -111
rect 2517 -145 2526 -111
rect 2474 -154 2526 -145
rect 2678 -111 2730 -102
rect 2678 -145 2687 -111
rect 2687 -145 2721 -111
rect 2721 -145 2730 -111
rect 2678 -154 2730 -145
rect 2882 -111 2934 -102
rect 2882 -145 2891 -111
rect 2891 -145 2925 -111
rect 2925 -145 2934 -111
rect 2882 -154 2934 -145
rect 3086 -111 3138 -102
rect 3086 -145 3095 -111
rect 3095 -145 3129 -111
rect 3129 -145 3138 -111
rect 3086 -154 3138 -145
rect 3290 -111 3342 -102
rect 3290 -145 3299 -111
rect 3299 -145 3333 -111
rect 3333 -145 3342 -111
rect 3290 -154 3342 -145
rect 3494 -111 3546 -102
rect 3494 -145 3503 -111
rect 3503 -145 3537 -111
rect 3537 -145 3546 -111
rect 3494 -154 3546 -145
rect 3698 -111 3750 -102
rect 3698 -145 3707 -111
rect 3707 -145 3741 -111
rect 3741 -145 3750 -111
rect 3698 -154 3750 -145
rect 3902 -111 3954 -102
rect 3902 -145 3911 -111
rect 3911 -145 3945 -111
rect 3945 -145 3954 -111
rect 3902 -154 3954 -145
rect 4106 -111 4158 -102
rect 4106 -145 4115 -111
rect 4115 -145 4149 -111
rect 4149 -145 4158 -111
rect 4106 -154 4158 -145
rect 4310 -111 4362 -102
rect 4310 -145 4319 -111
rect 4319 -145 4353 -111
rect 4353 -145 4362 -111
rect 4310 -154 4362 -145
rect 4514 -111 4566 -102
rect 4514 -145 4523 -111
rect 4523 -145 4557 -111
rect 4557 -145 4566 -111
rect 4514 -154 4566 -145
rect 4718 -111 4770 -102
rect 4718 -145 4727 -111
rect 4727 -145 4761 -111
rect 4761 -145 4770 -111
rect 4718 -154 4770 -145
rect 4922 -111 4974 -102
rect 4922 -145 4931 -111
rect 4931 -145 4965 -111
rect 4965 -145 4974 -111
rect 4922 -154 4974 -145
rect 5126 -111 5178 -102
rect 5126 -145 5135 -111
rect 5135 -145 5169 -111
rect 5169 -145 5178 -111
rect 5126 -154 5178 -145
rect 5330 -111 5382 -102
rect 5330 -145 5339 -111
rect 5339 -145 5373 -111
rect 5373 -145 5382 -111
rect 5330 -154 5382 -145
rect 5534 -111 5586 -102
rect 5534 -145 5543 -111
rect 5543 -145 5577 -111
rect 5577 -145 5586 -111
rect 5534 -154 5586 -145
rect 5738 -111 5790 -102
rect 5738 -145 5747 -111
rect 5747 -145 5781 -111
rect 5781 -145 5790 -111
rect 5738 -154 5790 -145
rect 5942 -111 5994 -102
rect 5942 -145 5951 -111
rect 5951 -145 5985 -111
rect 5985 -145 5994 -111
rect 5942 -154 5994 -145
rect 6146 -111 6198 -102
rect 6146 -145 6155 -111
rect 6155 -145 6189 -111
rect 6189 -145 6198 -111
rect 6146 -154 6198 -145
rect 6350 -111 6402 -102
rect 6350 -145 6359 -111
rect 6359 -145 6393 -111
rect 6393 -145 6402 -111
rect 6350 -154 6402 -145
rect 6554 -111 6606 -102
rect 6554 -145 6563 -111
rect 6563 -145 6597 -111
rect 6597 -145 6606 -111
rect 6554 -154 6606 -145
rect 6758 -111 6810 -102
rect 6758 -145 6767 -111
rect 6767 -145 6801 -111
rect 6801 -145 6810 -111
rect 6758 -154 6810 -145
rect 6962 -111 7014 -102
rect 6962 -145 6971 -111
rect 6971 -145 7005 -111
rect 7005 -145 7014 -111
rect 6962 -154 7014 -145
rect 7166 -111 7218 -102
rect 7166 -145 7175 -111
rect 7175 -145 7209 -111
rect 7209 -145 7218 -111
rect 7166 -154 7218 -145
rect 7370 -111 7422 -102
rect 7370 -145 7379 -111
rect 7379 -145 7413 -111
rect 7413 -145 7422 -111
rect 7370 -154 7422 -145
rect 7574 -111 7626 -102
rect 7574 -145 7583 -111
rect 7583 -145 7617 -111
rect 7617 -145 7626 -111
rect 7574 -154 7626 -145
rect 7778 -111 7830 -102
rect 7778 -145 7787 -111
rect 7787 -145 7821 -111
rect 7821 -145 7830 -111
rect 7778 -154 7830 -145
rect 7982 -111 8034 -102
rect 7982 -145 7991 -111
rect 7991 -145 8025 -111
rect 8025 -145 8034 -111
rect 7982 -154 8034 -145
rect 8186 -111 8238 -102
rect 8186 -145 8195 -111
rect 8195 -145 8229 -111
rect 8229 -145 8238 -111
rect 8186 -154 8238 -145
rect 8390 -111 8442 -102
rect 8390 -145 8399 -111
rect 8399 -145 8433 -111
rect 8433 -145 8442 -111
rect 8390 -154 8442 -145
rect 8594 -111 8646 -102
rect 8594 -145 8603 -111
rect 8603 -145 8637 -111
rect 8637 -145 8646 -111
rect 8594 -154 8646 -145
rect 8798 -111 8850 -102
rect 8798 -145 8807 -111
rect 8807 -145 8841 -111
rect 8841 -145 8850 -111
rect 8798 -154 8850 -145
rect 9002 -111 9054 -102
rect 9002 -145 9011 -111
rect 9011 -145 9045 -111
rect 9045 -145 9054 -111
rect 9002 -154 9054 -145
rect 9206 -111 9258 -102
rect 9206 -145 9215 -111
rect 9215 -145 9249 -111
rect 9249 -145 9258 -111
rect 9206 -154 9258 -145
rect 9410 -111 9462 -102
rect 9410 -145 9419 -111
rect 9419 -145 9453 -111
rect 9453 -145 9462 -111
rect 9410 -154 9462 -145
rect 9614 -111 9666 -102
rect 9614 -145 9623 -111
rect 9623 -145 9657 -111
rect 9657 -145 9666 -111
rect 9614 -154 9666 -145
rect 9818 -111 9870 -102
rect 9818 -145 9827 -111
rect 9827 -145 9861 -111
rect 9861 -145 9870 -111
rect 9818 -154 9870 -145
rect 10022 -111 10074 -102
rect 10022 -145 10031 -111
rect 10031 -145 10065 -111
rect 10065 -145 10074 -111
rect 10022 -154 10074 -145
rect 10226 -111 10278 -102
rect 10226 -145 10235 -111
rect 10235 -145 10269 -111
rect 10269 -145 10278 -111
rect 10226 -154 10278 -145
rect 10430 -111 10482 -102
rect 10430 -145 10439 -111
rect 10439 -145 10473 -111
rect 10473 -145 10482 -111
rect 10430 -154 10482 -145
rect 10634 -111 10686 -102
rect 10634 -145 10643 -111
rect 10643 -145 10677 -111
rect 10677 -145 10686 -111
rect 10634 -154 10686 -145
rect 10838 -111 10890 -102
rect 10838 -145 10847 -111
rect 10847 -145 10881 -111
rect 10881 -145 10890 -111
rect 10838 -154 10890 -145
rect 11042 -111 11094 -102
rect 11042 -145 11051 -111
rect 11051 -145 11085 -111
rect 11085 -145 11094 -111
rect 11042 -154 11094 -145
rect 11246 -111 11298 -102
rect 11246 -145 11255 -111
rect 11255 -145 11289 -111
rect 11289 -145 11298 -111
rect 11246 -154 11298 -145
rect 11450 -111 11502 -102
rect 11450 -145 11459 -111
rect 11459 -145 11493 -111
rect 11493 -145 11502 -111
rect 11450 -154 11502 -145
rect 11654 -111 11706 -102
rect 11654 -145 11663 -111
rect 11663 -145 11697 -111
rect 11697 -145 11706 -111
rect 11654 -154 11706 -145
rect 11858 -111 11910 -102
rect 11858 -145 11867 -111
rect 11867 -145 11901 -111
rect 11901 -145 11910 -111
rect 11858 -154 11910 -145
rect 12062 -111 12114 -102
rect 12062 -145 12071 -111
rect 12071 -145 12105 -111
rect 12105 -145 12114 -111
rect 12062 -154 12114 -145
rect 12266 -111 12318 -102
rect 12266 -145 12275 -111
rect 12275 -145 12309 -111
rect 12309 -145 12318 -111
rect 12266 -154 12318 -145
rect 12470 -111 12522 -102
rect 12470 -145 12479 -111
rect 12479 -145 12513 -111
rect 12513 -145 12522 -111
rect 12470 -154 12522 -145
rect 12674 -111 12726 -102
rect 12674 -145 12683 -111
rect 12683 -145 12717 -111
rect 12717 -145 12726 -111
rect 12674 -154 12726 -145
rect 12878 -111 12930 -102
rect 12878 -145 12887 -111
rect 12887 -145 12921 -111
rect 12921 -145 12930 -111
rect 12878 -154 12930 -145
<< metal2 >>
rect 61 240 13145 268
rect 12 -102 13082 -96
rect 12 -154 26 -102
rect 78 -154 230 -102
rect 282 -154 434 -102
rect 486 -154 638 -102
rect 690 -154 842 -102
rect 894 -154 1046 -102
rect 1098 -154 1250 -102
rect 1302 -154 1454 -102
rect 1506 -154 1658 -102
rect 1710 -154 1862 -102
rect 1914 -154 2066 -102
rect 2118 -154 2270 -102
rect 2322 -154 2474 -102
rect 2526 -154 2678 -102
rect 2730 -154 2882 -102
rect 2934 -154 3086 -102
rect 3138 -154 3290 -102
rect 3342 -154 3494 -102
rect 3546 -154 3698 -102
rect 3750 -154 3902 -102
rect 3954 -154 4106 -102
rect 4158 -154 4310 -102
rect 4362 -154 4514 -102
rect 4566 -154 4718 -102
rect 4770 -154 4922 -102
rect 4974 -154 5126 -102
rect 5178 -154 5330 -102
rect 5382 -154 5534 -102
rect 5586 -154 5738 -102
rect 5790 -154 5942 -102
rect 5994 -154 6146 -102
rect 6198 -154 6350 -102
rect 6402 -154 6554 -102
rect 6606 -154 6758 -102
rect 6810 -154 6962 -102
rect 7014 -154 7166 -102
rect 7218 -154 7370 -102
rect 7422 -154 7574 -102
rect 7626 -154 7778 -102
rect 7830 -154 7982 -102
rect 8034 -154 8186 -102
rect 8238 -154 8390 -102
rect 8442 -154 8594 -102
rect 8646 -154 8798 -102
rect 8850 -154 9002 -102
rect 9054 -154 9206 -102
rect 9258 -154 9410 -102
rect 9462 -154 9614 -102
rect 9666 -154 9818 -102
rect 9870 -154 10022 -102
rect 10074 -154 10226 -102
rect 10278 -154 10430 -102
rect 10482 -154 10634 -102
rect 10686 -154 10838 -102
rect 10890 -154 11042 -102
rect 11094 -154 11246 -102
rect 11298 -154 11450 -102
rect 11502 -154 11654 -102
rect 11706 -154 11858 -102
rect 11910 -154 12062 -102
rect 12114 -154 12266 -102
rect 12318 -154 12470 -102
rect 12522 -154 12674 -102
rect 12726 -154 12878 -102
rect 12930 -154 13082 -102
rect 12 -160 13082 -154
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_0
timestamp 1581320205
transform 1 0 12852 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_1
timestamp 1581320205
transform 1 0 12648 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_2
timestamp 1581320205
transform 1 0 12444 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_3
timestamp 1581320205
transform 1 0 12240 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_4
timestamp 1581320205
transform 1 0 12036 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_5
timestamp 1581320205
transform 1 0 11832 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_6
timestamp 1581320205
transform 1 0 11628 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_7
timestamp 1581320205
transform 1 0 11424 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_8
timestamp 1581320205
transform 1 0 11220 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_9
timestamp 1581320205
transform 1 0 11016 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_10
timestamp 1581320205
transform 1 0 10812 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_11
timestamp 1581320205
transform 1 0 10608 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_12
timestamp 1581320205
transform 1 0 10404 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_13
timestamp 1581320205
transform 1 0 10200 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_14
timestamp 1581320205
transform 1 0 9996 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_15
timestamp 1581320205
transform 1 0 9792 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_16
timestamp 1581320205
transform 1 0 9588 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_17
timestamp 1581320205
transform 1 0 9384 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_18
timestamp 1581320205
transform 1 0 9180 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_19
timestamp 1581320205
transform 1 0 8976 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_20
timestamp 1581320205
transform 1 0 8772 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_21
timestamp 1581320205
transform 1 0 8568 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_22
timestamp 1581320205
transform 1 0 8364 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_23
timestamp 1581320205
transform 1 0 8160 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_24
timestamp 1581320205
transform 1 0 7956 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_25
timestamp 1581320205
transform 1 0 7752 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_26
timestamp 1581320205
transform 1 0 7548 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_27
timestamp 1581320205
transform 1 0 7344 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_28
timestamp 1581320205
transform 1 0 7140 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_29
timestamp 1581320205
transform 1 0 6936 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_30
timestamp 1581320205
transform 1 0 6732 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_31
timestamp 1581320205
transform 1 0 6528 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_32
timestamp 1581320205
transform 1 0 6324 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_33
timestamp 1581320205
transform 1 0 6120 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_34
timestamp 1581320205
transform 1 0 5916 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_35
timestamp 1581320205
transform 1 0 5712 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_36
timestamp 1581320205
transform 1 0 5508 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_37
timestamp 1581320205
transform 1 0 5304 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_38
timestamp 1581320205
transform 1 0 5100 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_39
timestamp 1581320205
transform 1 0 4896 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_40
timestamp 1581320205
transform 1 0 4692 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_41
timestamp 1581320205
transform 1 0 4488 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_42
timestamp 1581320205
transform 1 0 4284 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_43
timestamp 1581320205
transform 1 0 4080 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_44
timestamp 1581320205
transform 1 0 3876 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_45
timestamp 1581320205
transform 1 0 3672 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_46
timestamp 1581320205
transform 1 0 3468 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_47
timestamp 1581320205
transform 1 0 3264 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_48
timestamp 1581320205
transform 1 0 3060 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_49
timestamp 1581320205
transform 1 0 2856 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_50
timestamp 1581320205
transform 1 0 2652 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_51
timestamp 1581320205
transform 1 0 2448 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_52
timestamp 1581320205
transform 1 0 2244 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_53
timestamp 1581320205
transform 1 0 2040 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_54
timestamp 1581320205
transform 1 0 1836 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_55
timestamp 1581320205
transform 1 0 1632 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_56
timestamp 1581320205
transform 1 0 1428 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_57
timestamp 1581320205
transform 1 0 1224 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_58
timestamp 1581320205
transform 1 0 1020 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_59
timestamp 1581320205
transform 1 0 816 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_60
timestamp 1581320205
transform 1 0 612 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_61
timestamp 1581320205
transform 1 0 408 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_62
timestamp 1581320205
transform 1 0 204 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_63
timestamp 1581320205
transform 1 0 0 0 1 0
box 0 -212 232 184
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_0
timestamp 1581320205
transform 1 0 13098 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_1
timestamp 1581320205
transform 1 0 11466 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_2
timestamp 1581320205
transform 1 0 9834 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_3
timestamp 1581320205
transform 1 0 8202 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_4
timestamp 1581320205
transform 1 0 6570 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_5
timestamp 1581320205
transform 1 0 4938 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_6
timestamp 1581320205
transform 1 0 3306 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_7
timestamp 1581320205
transform 1 0 1674 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_8
timestamp 1581320205
transform 1 0 42 0 1 204
box 0 17 66 83
<< labels >>
rlabel nwell s 13164 408 13164 408 4 upper right
rlabel metal2 s 61 240 89 268 4 gate
port 3 nsew
rlabel metal2 s 13117 240 13145 268 4 precharge_r
port 5 nsew
rlabel metal1 s 122 86 150 114 4 pre_bl0_out
port 7 nsew
rlabel metal1 s 326 86 354 114 4 pre_bl1_out
port 9 nsew
rlabel metal1 s 530 86 558 114 4 pre_bl2_out
port 11 nsew
rlabel metal1 s 734 86 762 114 4 pre_bl3_out
port 13 nsew
rlabel metal1 s 938 86 966 114 4 pre_bl4_out
port 15 nsew
rlabel metal1 s 1142 86 1170 114 4 pre_bl5_out
port 17 nsew
rlabel metal1 s 1346 86 1374 114 4 pre_bl6_out
port 19 nsew
rlabel metal1 s 1550 86 1578 114 4 pre_bl7_out
port 21 nsew
rlabel metal1 s 1754 86 1782 114 4 pre_bl8_out
port 23 nsew
rlabel metal1 s 1958 86 1986 114 4 pre_bl9_out
port 25 nsew
rlabel metal1 s 2162 86 2190 114 4 pre_bl10_out
port 27 nsew
rlabel metal1 s 2366 86 2394 114 4 pre_bl11_out
port 29 nsew
rlabel metal1 s 2570 86 2598 114 4 pre_bl12_out
port 31 nsew
rlabel metal1 s 2774 86 2802 114 4 pre_bl13_out
port 33 nsew
rlabel metal1 s 2978 86 3006 114 4 pre_bl14_out
port 35 nsew
rlabel metal1 s 3182 86 3210 114 4 pre_bl15_out
port 37 nsew
rlabel metal1 s 3386 86 3414 114 4 pre_bl16_out
port 39 nsew
rlabel metal1 s 3590 86 3618 114 4 pre_bl17_out
port 41 nsew
rlabel metal1 s 3794 86 3822 114 4 pre_bl18_out
port 43 nsew
rlabel metal1 s 3998 86 4026 114 4 pre_bl19_out
port 45 nsew
rlabel metal1 s 4202 86 4230 114 4 pre_bl20_out
port 47 nsew
rlabel metal1 s 4406 86 4434 114 4 pre_bl21_out
port 49 nsew
rlabel metal1 s 4610 86 4638 114 4 pre_bl22_out
port 51 nsew
rlabel metal1 s 4814 86 4842 114 4 pre_bl23_out
port 53 nsew
rlabel metal1 s 5018 86 5046 114 4 pre_bl24_out
port 55 nsew
rlabel metal1 s 5222 86 5250 114 4 pre_bl25_out
port 57 nsew
rlabel metal1 s 5426 86 5454 114 4 pre_bl26_out
port 59 nsew
rlabel metal1 s 5630 86 5658 114 4 pre_bl27_out
port 61 nsew
rlabel metal1 s 5834 86 5862 114 4 pre_bl28_out
port 63 nsew
rlabel metal1 s 6038 86 6066 114 4 pre_bl29_out
port 65 nsew
rlabel metal1 s 6242 86 6270 114 4 pre_bl30_out
port 67 nsew
rlabel metal1 s 6446 86 6474 114 4 pre_bl31_out
port 69 nsew
rlabel metal1 s 6650 86 6678 114 4 pre_bl32_out
port 71 nsew
rlabel metal1 s 6854 86 6882 114 4 pre_bl33_out
port 73 nsew
rlabel metal1 s 7058 86 7086 114 4 pre_bl34_out
port 75 nsew
rlabel metal1 s 7262 86 7290 114 4 pre_bl35_out
port 77 nsew
rlabel metal1 s 7466 86 7494 114 4 pre_bl36_out
port 79 nsew
rlabel metal1 s 7670 86 7698 114 4 pre_bl37_out
port 81 nsew
rlabel metal1 s 7874 86 7902 114 4 pre_bl38_out
port 83 nsew
rlabel metal1 s 8078 86 8106 114 4 pre_bl39_out
port 85 nsew
rlabel metal1 s 8282 86 8310 114 4 pre_bl40_out
port 87 nsew
rlabel metal1 s 8486 86 8514 114 4 pre_bl41_out
port 89 nsew
rlabel metal1 s 8690 86 8718 114 4 pre_bl42_out
port 91 nsew
rlabel metal1 s 8894 86 8922 114 4 pre_bl43_out
port 93 nsew
rlabel metal1 s 9098 86 9126 114 4 pre_bl44_out
port 95 nsew
rlabel metal1 s 9302 86 9330 114 4 pre_bl45_out
port 97 nsew
rlabel metal1 s 9506 86 9534 114 4 pre_bl46_out
port 99 nsew
rlabel metal1 s 9710 86 9738 114 4 pre_bl47_out
port 101 nsew
rlabel metal1 s 9914 86 9942 114 4 pre_bl48_out
port 103 nsew
rlabel metal1 s 10118 86 10146 114 4 pre_bl49_out
port 105 nsew
rlabel metal1 s 10322 86 10350 114 4 pre_bl50_out
port 107 nsew
rlabel metal1 s 10526 86 10554 114 4 pre_bl51_out
port 109 nsew
rlabel metal1 s 10730 86 10758 114 4 pre_bl52_out
port 111 nsew
rlabel metal1 s 10934 86 10962 114 4 pre_bl53_out
port 113 nsew
rlabel metal1 s 11138 86 11166 114 4 pre_bl54_out
port 115 nsew
rlabel metal1 s 11342 86 11370 114 4 pre_bl55_out
port 117 nsew
rlabel metal1 s 11546 86 11574 114 4 pre_bl56_out
port 119 nsew
rlabel metal1 s 11750 86 11778 114 4 pre_bl57_out
port 121 nsew
rlabel metal1 s 11954 86 11982 114 4 pre_bl58_out
port 123 nsew
rlabel metal1 s 12158 86 12186 114 4 pre_bl59_out
port 125 nsew
rlabel metal1 s 12362 86 12390 114 4 pre_bl60_out
port 127 nsew
rlabel metal1 s 12566 86 12594 114 4 pre_bl61_out
port 129 nsew
rlabel metal1 s 12770 86 12798 114 4 pre_bl62_out
port 131 nsew
rlabel metal1 s 12974 86 13002 114 4 pre_bl63_out
port 133 nsew
rlabel metal2 s 12 -160 40 -96 4 vdd
port 135 nsew
<< properties >>
string FIXED_BBOX 12875 -161 12933 -160
<< end >>
