magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1296 -1277 2312 3436
<< nwell >>
rect -36 1017 1052 2176
<< pwell >>
rect 28 159 878 477
rect 28 25 982 159
<< scnmos >>
rect 114 51 144 451
rect 222 51 252 451
rect 330 51 360 451
rect 438 51 468 451
rect 546 51 576 451
rect 654 51 684 451
rect 762 51 792 451
<< scpmos >>
rect 114 1468 144 2068
rect 222 1468 252 2068
rect 330 1468 360 2068
rect 438 1468 468 2068
rect 546 1468 576 2068
rect 654 1468 684 2068
rect 762 1468 792 2068
<< ndiff >>
rect 54 268 114 451
rect 54 234 62 268
rect 96 234 114 268
rect 54 51 114 234
rect 144 268 222 451
rect 144 234 166 268
rect 200 234 222 268
rect 144 51 222 234
rect 252 268 330 451
rect 252 234 274 268
rect 308 234 330 268
rect 252 51 330 234
rect 360 268 438 451
rect 360 234 382 268
rect 416 234 438 268
rect 360 51 438 234
rect 468 268 546 451
rect 468 234 490 268
rect 524 234 546 268
rect 468 51 546 234
rect 576 268 654 451
rect 576 234 598 268
rect 632 234 654 268
rect 576 51 654 234
rect 684 268 762 451
rect 684 234 706 268
rect 740 234 762 268
rect 684 51 762 234
rect 792 268 852 451
rect 792 234 810 268
rect 844 234 852 268
rect 792 51 852 234
<< pdiff >>
rect 54 1785 114 2068
rect 54 1751 62 1785
rect 96 1751 114 1785
rect 54 1468 114 1751
rect 144 1785 222 2068
rect 144 1751 166 1785
rect 200 1751 222 1785
rect 144 1468 222 1751
rect 252 1785 330 2068
rect 252 1751 274 1785
rect 308 1751 330 1785
rect 252 1468 330 1751
rect 360 1785 438 2068
rect 360 1751 382 1785
rect 416 1751 438 1785
rect 360 1468 438 1751
rect 468 1785 546 2068
rect 468 1751 490 1785
rect 524 1751 546 1785
rect 468 1468 546 1751
rect 576 1785 654 2068
rect 576 1751 598 1785
rect 632 1751 654 1785
rect 576 1468 654 1751
rect 684 1785 762 2068
rect 684 1751 706 1785
rect 740 1751 762 1785
rect 684 1468 762 1751
rect 792 1785 852 2068
rect 792 1751 810 1785
rect 844 1751 852 1785
rect 792 1468 852 1751
<< ndiffc >>
rect 62 234 96 268
rect 166 234 200 268
rect 274 234 308 268
rect 382 234 416 268
rect 490 234 524 268
rect 598 234 632 268
rect 706 234 740 268
rect 810 234 844 268
<< pdiffc >>
rect 62 1751 96 1785
rect 166 1751 200 1785
rect 274 1751 308 1785
rect 382 1751 416 1785
rect 490 1751 524 1785
rect 598 1751 632 1785
rect 706 1751 740 1785
rect 810 1751 844 1785
<< psubdiff >>
rect 906 109 956 133
rect 906 75 914 109
rect 948 75 956 109
rect 906 51 956 75
<< nsubdiff >>
rect 906 2031 956 2055
rect 906 1997 914 2031
rect 948 1997 956 2031
rect 906 1973 956 1997
<< psubdiffcont >>
rect 914 75 948 109
<< nsubdiffcont >>
rect 914 1997 948 2031
<< poly >>
rect 114 2068 144 2094
rect 222 2068 252 2094
rect 330 2068 360 2094
rect 438 2068 468 2094
rect 546 2068 576 2094
rect 654 2068 684 2094
rect 762 2068 792 2094
rect 114 1442 144 1468
rect 222 1442 252 1468
rect 330 1442 360 1468
rect 438 1442 468 1468
rect 546 1442 576 1468
rect 654 1442 684 1468
rect 762 1442 792 1468
rect 114 1412 792 1442
rect 114 1042 144 1412
rect 48 1026 144 1042
rect 48 992 64 1026
rect 98 992 144 1026
rect 48 976 144 992
rect 114 507 144 976
rect 114 477 792 507
rect 114 451 144 477
rect 222 451 252 477
rect 330 451 360 477
rect 438 451 468 477
rect 546 451 576 477
rect 654 451 684 477
rect 762 451 792 477
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
rect 438 25 468 51
rect 546 25 576 51
rect 654 25 684 51
rect 762 25 792 51
<< polycont >>
rect 64 992 98 1026
<< locali >>
rect 0 2102 1016 2136
rect 62 1785 96 2102
rect 62 1735 96 1751
rect 166 1785 200 1801
rect 166 1701 200 1751
rect 274 1785 308 2102
rect 274 1735 308 1751
rect 382 1785 416 1801
rect 382 1701 416 1751
rect 490 1785 524 2102
rect 490 1735 524 1751
rect 598 1785 632 1801
rect 598 1701 632 1751
rect 706 1785 740 2102
rect 914 2031 948 2102
rect 914 1981 948 1997
rect 706 1735 740 1751
rect 810 1785 844 1801
rect 810 1701 844 1751
rect 166 1667 844 1701
rect 64 1026 98 1042
rect 64 976 98 992
rect 488 1026 522 1667
rect 488 992 539 1026
rect 488 352 522 992
rect 166 318 844 352
rect 62 268 96 284
rect 62 17 96 234
rect 166 268 200 318
rect 166 218 200 234
rect 274 268 308 284
rect 274 17 308 234
rect 382 268 416 318
rect 382 218 416 234
rect 490 268 524 284
rect 490 17 524 234
rect 598 268 632 318
rect 598 218 632 234
rect 706 268 740 284
rect 706 17 740 234
rect 810 268 844 318
rect 810 218 844 234
rect 914 109 948 125
rect 914 17 948 75
rect 0 -17 1016 17
<< labels >>
rlabel locali s 81 1009 81 1009 4 A
port 1 nsew
rlabel locali s 522 1009 522 1009 4 Z
port 2 nsew
rlabel locali s 508 0 508 0 4 gnd
port 3 nsew
rlabel locali s 508 2119 508 2119 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1016 1684
<< end >>
