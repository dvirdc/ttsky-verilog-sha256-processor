magic
tech sky130A
magscale 1 2
timestamp 1581479693
<< checkpaint >>
rect -1296 -1277 1772 3946
<< nwell >>
rect -36 1262 512 2686
<< pwell >>
rect 28 159 338 329
rect 28 25 442 159
<< scnmos >>
rect 114 51 144 303
rect 222 51 252 303
<< scpmos >>
rect 114 2178 144 2578
rect 222 2178 252 2578
<< ndiff >>
rect 54 194 114 303
rect 54 160 62 194
rect 96 160 114 194
rect 54 51 114 160
rect 144 194 222 303
rect 144 160 166 194
rect 200 160 222 194
rect 144 51 222 160
rect 252 194 312 303
rect 252 160 270 194
rect 304 160 312 194
rect 252 51 312 160
<< pdiff >>
rect 54 2395 114 2578
rect 54 2361 62 2395
rect 96 2361 114 2395
rect 54 2178 114 2361
rect 144 2395 222 2578
rect 144 2361 166 2395
rect 200 2361 222 2395
rect 144 2178 222 2361
rect 252 2395 312 2578
rect 252 2361 270 2395
rect 304 2361 312 2395
rect 252 2178 312 2361
<< ndiffc >>
rect 62 160 96 194
rect 166 160 200 194
rect 270 160 304 194
<< pdiffc >>
rect 62 2361 96 2395
rect 166 2361 200 2395
rect 270 2361 304 2395
<< psubdiff >>
rect 366 109 416 133
rect 366 75 374 109
rect 408 75 416 109
rect 366 51 416 75
<< nsubdiff >>
rect 366 2541 416 2565
rect 366 2507 374 2541
rect 408 2507 416 2541
rect 366 2483 416 2507
<< psubdiffcont >>
rect 374 75 408 109
<< nsubdiffcont >>
rect 374 2507 408 2541
<< poly >>
rect 114 2578 144 2604
rect 222 2578 252 2604
rect 114 2152 144 2178
rect 222 2152 252 2178
rect 114 2122 252 2152
rect 114 1310 144 2122
rect 48 1294 144 1310
rect 48 1260 64 1294
rect 98 1260 144 1294
rect 48 1244 144 1260
rect 114 359 144 1244
rect 114 329 252 359
rect 114 303 144 329
rect 222 303 252 329
rect 114 25 144 51
rect 222 25 252 51
<< polycont >>
rect 64 1260 98 1294
<< locali >>
rect 0 2612 476 2646
rect 62 2395 96 2612
rect 62 2345 96 2361
rect 166 2395 200 2411
rect 64 1294 98 1310
rect 64 1244 98 1260
rect 166 1294 200 2361
rect 270 2395 304 2612
rect 374 2541 408 2612
rect 374 2491 408 2507
rect 270 2345 304 2361
rect 166 1260 217 1294
rect 62 194 96 210
rect 62 17 96 160
rect 166 194 200 1260
rect 166 144 200 160
rect 270 194 304 210
rect 270 17 304 160
rect 374 109 408 125
rect 374 17 408 75
rect 0 -17 476 17
<< labels >>
rlabel locali s 81 1277 81 1277 4 A
port 1 nsew
rlabel locali s 200 1277 200 1277 4 Z
port 2 nsew
rlabel locali s 238 0 238 0 4 gnd
port 3 nsew
rlabel locali s 238 2629 238 2629 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 476 2294
<< end >>
