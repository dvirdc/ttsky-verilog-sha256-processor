magic
tech sky130A
magscale 1 2
timestamp 1581398725
<< checkpaint >>
rect -1216 -1310 6970 1559
<< locali >>
rect 60 51 94 117
rect 2506 51 2540 101
rect 2446 17 2540 51
rect 3275 17 5692 51
<< metal1 >>
rect 448 0 476 204
rect 1696 0 1724 204
rect 3294 0 3322 204
rect 4942 0 4970 204
use sky130_rom_krom_pinv_dec_0  sky130_rom_krom_pinv_dec_0_0
timestamp 1581398725
transform 1 0 0 0 1 0
box 44 -50 2464 299
use sky130_rom_krom_pinv_dec_1  sky130_rom_krom_pinv_dec_1_0
timestamp 1581398725
transform 1 0 2446 0 1 0
box 44 -50 3264 299
<< labels >>
rlabel locali s 4483 34 4483 34 4 Z
port 2 nsew
rlabel locali s 77 84 77 84 4 A
port 3 nsew
rlabel metal1 s 1696 0 1724 204 4 vdd
port 5 nsew
rlabel metal1 s 4942 0 4970 204 4 vdd
port 5 nsew
rlabel metal1 s 3294 0 3322 204 4 gnd
port 7 nsew
rlabel metal1 s 448 0 476 204 4 gnd
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 5692 204
<< end >>
