magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1266 -1344 2305 3164
<< poly >>
rect 0 1756 66 1772
rect 0 1722 16 1756
rect 50 1754 66 1756
rect 716 1756 782 1772
rect 716 1754 732 1756
rect 50 1724 732 1754
rect 50 1722 66 1724
rect 0 1706 66 1722
rect 716 1722 732 1724
rect 766 1722 782 1756
rect 716 1706 782 1722
rect 0 1552 66 1568
rect 0 1518 16 1552
rect 50 1550 66 1552
rect 716 1552 782 1568
rect 716 1550 732 1552
rect 50 1520 732 1550
rect 50 1518 66 1520
rect 0 1502 66 1518
rect 716 1518 732 1520
rect 766 1518 782 1552
rect 716 1502 782 1518
rect 0 1348 66 1364
rect 0 1314 16 1348
rect 50 1346 66 1348
rect 716 1348 782 1364
rect 716 1346 732 1348
rect 50 1316 732 1346
rect 50 1314 66 1316
rect 0 1298 66 1314
rect 716 1314 732 1316
rect 766 1314 782 1348
rect 716 1298 782 1314
rect 0 1144 66 1160
rect 0 1110 16 1144
rect 50 1142 66 1144
rect 716 1144 782 1160
rect 716 1142 732 1144
rect 50 1112 732 1142
rect 50 1110 66 1112
rect 0 1094 66 1110
rect 716 1110 732 1112
rect 766 1110 782 1144
rect 716 1094 782 1110
rect 0 940 66 956
rect 0 906 16 940
rect 50 938 66 940
rect 716 940 782 956
rect 716 938 732 940
rect 50 908 732 938
rect 50 906 66 908
rect 0 890 66 906
rect 716 906 732 908
rect 766 906 782 940
rect 716 890 782 906
<< polycont >>
rect 16 1722 50 1756
rect 732 1722 766 1756
rect 16 1518 50 1552
rect 732 1518 766 1552
rect 16 1314 50 1348
rect 732 1314 766 1348
rect 16 1110 50 1144
rect 732 1110 766 1144
rect 16 906 50 940
rect 732 906 766 940
<< locali >>
rect 16 1756 50 1772
rect 16 1706 50 1722
rect 732 1756 766 1772
rect 732 1706 766 1722
rect 28 1620 44 1654
rect 78 1620 94 1654
rect 744 1620 760 1654
rect 794 1620 810 1654
rect 16 1552 50 1568
rect 16 1502 50 1518
rect 732 1552 766 1568
rect 732 1502 766 1518
rect 28 1416 44 1450
rect 78 1416 94 1450
rect 744 1416 760 1450
rect 794 1416 810 1450
rect 16 1348 50 1364
rect 16 1298 50 1314
rect 732 1348 766 1364
rect 732 1298 766 1314
rect 28 1212 44 1246
rect 78 1212 94 1246
rect 744 1212 760 1246
rect 794 1212 810 1246
rect 16 1144 50 1160
rect 16 1094 50 1110
rect 732 1144 766 1160
rect 732 1094 766 1110
rect 28 1008 44 1042
rect 78 1008 94 1042
rect 744 1008 760 1042
rect 794 1008 810 1042
rect 16 940 50 956
rect 16 890 50 906
rect 732 940 766 956
rect 732 890 766 906
<< viali >>
rect 16 1722 50 1756
rect 732 1722 766 1756
rect 44 1620 78 1654
rect 760 1620 794 1654
rect 16 1518 50 1552
rect 732 1518 766 1552
rect 44 1416 78 1450
rect 760 1416 794 1450
rect 16 1314 50 1348
rect 732 1314 766 1348
rect 44 1212 78 1246
rect 760 1212 794 1246
rect 16 1110 50 1144
rect 732 1110 766 1144
rect 44 1008 78 1042
rect 760 1008 794 1042
rect 16 906 50 940
rect 732 906 766 940
<< metal1 >>
rect 29 1840 35 1892
rect 87 1880 93 1892
rect 745 1880 751 1892
rect 87 1852 751 1880
rect 87 1840 93 1852
rect 745 1840 751 1852
rect 803 1840 809 1892
rect 8 1765 59 1772
rect 724 1765 775 1772
rect 1 1713 7 1765
rect 59 1713 65 1765
rect 717 1713 723 1765
rect 775 1753 781 1765
rect 775 1725 1045 1753
rect 775 1713 781 1725
rect 8 1706 59 1713
rect 724 1706 775 1713
rect 35 1663 87 1669
rect 35 1605 87 1611
rect 751 1663 803 1669
rect 751 1605 803 1611
rect 8 1561 59 1568
rect 724 1561 775 1568
rect 1 1509 7 1561
rect 59 1509 65 1561
rect 717 1509 723 1561
rect 775 1509 781 1561
rect 8 1502 59 1509
rect 724 1502 775 1509
rect 35 1459 87 1465
rect 35 1401 87 1407
rect 751 1459 803 1465
rect 751 1401 803 1407
rect 8 1357 59 1364
rect 724 1357 775 1364
rect 1 1305 7 1357
rect 59 1305 65 1357
rect 717 1305 723 1357
rect 775 1305 781 1357
rect 8 1298 59 1305
rect 724 1298 775 1305
rect 35 1255 87 1261
rect 35 1197 87 1203
rect 751 1255 803 1261
rect 751 1197 803 1203
rect 8 1153 59 1160
rect 724 1153 775 1160
rect 1 1101 7 1153
rect 59 1101 65 1153
rect 717 1101 723 1153
rect 775 1101 781 1153
rect 8 1094 59 1101
rect 724 1094 775 1101
rect 35 1051 87 1057
rect 35 993 87 999
rect 751 1051 803 1057
rect 751 993 803 999
rect 8 949 59 956
rect 724 949 775 956
rect 1 897 7 949
rect 59 897 65 949
rect 717 897 723 949
rect 775 897 781 949
rect 8 890 59 897
rect 724 890 775 897
rect 232 -14 260 873
rect 436 -14 464 873
rect 640 -14 668 873
rect 1017 396 1045 1725
rect 791 368 1045 396
<< via1 >>
rect 35 1840 87 1892
rect 751 1840 803 1892
rect 7 1756 59 1765
rect 7 1722 16 1756
rect 16 1722 50 1756
rect 50 1722 59 1756
rect 7 1713 59 1722
rect 723 1756 775 1765
rect 723 1722 732 1756
rect 732 1722 766 1756
rect 766 1722 775 1756
rect 723 1713 775 1722
rect 35 1654 87 1663
rect 35 1620 44 1654
rect 44 1620 78 1654
rect 78 1620 87 1654
rect 35 1611 87 1620
rect 751 1654 803 1663
rect 751 1620 760 1654
rect 760 1620 794 1654
rect 794 1620 803 1654
rect 751 1611 803 1620
rect 7 1552 59 1561
rect 7 1518 16 1552
rect 16 1518 50 1552
rect 50 1518 59 1552
rect 7 1509 59 1518
rect 723 1552 775 1561
rect 723 1518 732 1552
rect 732 1518 766 1552
rect 766 1518 775 1552
rect 723 1509 775 1518
rect 35 1450 87 1459
rect 35 1416 44 1450
rect 44 1416 78 1450
rect 78 1416 87 1450
rect 35 1407 87 1416
rect 751 1450 803 1459
rect 751 1416 760 1450
rect 760 1416 794 1450
rect 794 1416 803 1450
rect 751 1407 803 1416
rect 7 1348 59 1357
rect 7 1314 16 1348
rect 16 1314 50 1348
rect 50 1314 59 1348
rect 7 1305 59 1314
rect 723 1348 775 1357
rect 723 1314 732 1348
rect 732 1314 766 1348
rect 766 1314 775 1348
rect 723 1305 775 1314
rect 35 1246 87 1255
rect 35 1212 44 1246
rect 44 1212 78 1246
rect 78 1212 87 1246
rect 35 1203 87 1212
rect 751 1246 803 1255
rect 751 1212 760 1246
rect 760 1212 794 1246
rect 794 1212 803 1246
rect 751 1203 803 1212
rect 7 1144 59 1153
rect 7 1110 16 1144
rect 16 1110 50 1144
rect 50 1110 59 1144
rect 7 1101 59 1110
rect 723 1144 775 1153
rect 723 1110 732 1144
rect 732 1110 766 1144
rect 766 1110 775 1144
rect 723 1101 775 1110
rect 35 1042 87 1051
rect 35 1008 44 1042
rect 44 1008 78 1042
rect 78 1008 87 1042
rect 35 999 87 1008
rect 751 1042 803 1051
rect 751 1008 760 1042
rect 760 1008 794 1042
rect 794 1008 803 1042
rect 751 999 803 1008
rect 7 940 59 949
rect 7 906 16 940
rect 16 906 50 940
rect 50 906 59 940
rect 7 897 59 906
rect 723 940 775 949
rect 723 906 732 940
rect 732 906 766 940
rect 766 906 775 940
rect 723 897 775 906
<< metal2 >>
rect 33 1895 89 1904
rect 33 1830 89 1839
rect 749 1895 805 1904
rect 749 1830 805 1839
rect 7 1765 59 1771
rect 1 1718 7 1761
rect 723 1765 775 1771
rect 59 1753 65 1761
rect 717 1753 723 1761
rect 59 1725 723 1753
rect 59 1718 65 1725
rect 717 1718 723 1725
rect 7 1707 59 1713
rect 775 1718 781 1761
rect 723 1707 775 1713
rect 24 1609 33 1665
rect 89 1609 98 1665
rect 740 1609 749 1665
rect 805 1609 814 1665
rect 7 1561 59 1567
rect 1 1514 7 1557
rect 723 1561 775 1567
rect 59 1549 65 1557
rect 717 1549 723 1557
rect 59 1521 723 1549
rect 59 1514 65 1521
rect 717 1514 723 1521
rect 7 1503 59 1509
rect 775 1514 781 1557
rect 723 1503 775 1509
rect 24 1405 33 1461
rect 89 1405 98 1461
rect 740 1405 749 1461
rect 805 1405 814 1461
rect 7 1357 59 1363
rect 1 1310 7 1353
rect 723 1357 775 1363
rect 59 1345 65 1353
rect 717 1345 723 1353
rect 59 1317 723 1345
rect 59 1310 65 1317
rect 717 1310 723 1317
rect 7 1299 59 1305
rect 775 1310 781 1353
rect 723 1299 775 1305
rect 24 1201 33 1257
rect 89 1201 98 1257
rect 740 1201 749 1257
rect 805 1201 814 1257
rect 7 1153 59 1159
rect 1 1106 7 1149
rect 723 1153 775 1159
rect 59 1141 65 1149
rect 717 1141 723 1149
rect 59 1113 723 1141
rect 59 1106 65 1113
rect 717 1106 723 1113
rect 7 1095 59 1101
rect 775 1106 781 1149
rect 723 1095 775 1101
rect 24 997 33 1053
rect 89 997 98 1053
rect 740 997 749 1053
rect 805 997 814 1053
rect 7 949 59 955
rect 1 902 7 945
rect 723 949 775 955
rect 59 937 65 945
rect 717 937 723 945
rect 59 909 723 937
rect 59 902 65 909
rect 717 902 723 909
rect 7 891 59 897
rect 775 902 781 945
rect 723 891 775 897
rect 61 368 89 396
rect 12 -32 40 32
<< via2 >>
rect 33 1892 89 1895
rect 33 1840 35 1892
rect 35 1840 87 1892
rect 87 1840 89 1892
rect 33 1839 89 1840
rect 749 1892 805 1895
rect 749 1840 751 1892
rect 751 1840 803 1892
rect 803 1840 805 1892
rect 749 1839 805 1840
rect 33 1663 89 1665
rect 33 1611 35 1663
rect 35 1611 87 1663
rect 87 1611 89 1663
rect 33 1609 89 1611
rect 749 1663 805 1665
rect 749 1611 751 1663
rect 751 1611 803 1663
rect 803 1611 805 1663
rect 749 1609 805 1611
rect 33 1459 89 1461
rect 33 1407 35 1459
rect 35 1407 87 1459
rect 87 1407 89 1459
rect 33 1405 89 1407
rect 749 1459 805 1461
rect 749 1407 751 1459
rect 751 1407 803 1459
rect 803 1407 805 1459
rect 749 1405 805 1407
rect 33 1255 89 1257
rect 33 1203 35 1255
rect 35 1203 87 1255
rect 87 1203 89 1255
rect 33 1201 89 1203
rect 749 1255 805 1257
rect 749 1203 751 1255
rect 751 1203 803 1255
rect 803 1203 805 1255
rect 749 1201 805 1203
rect 33 1051 89 1053
rect 33 999 35 1051
rect 35 999 87 1051
rect 87 999 89 1051
rect 33 997 89 999
rect 749 1051 805 1053
rect 749 999 751 1051
rect 751 999 803 1051
rect 803 999 805 1051
rect 749 997 805 999
<< metal3 >>
rect 28 1895 94 1900
rect 28 1839 33 1895
rect 89 1839 94 1895
rect 28 1834 94 1839
rect 744 1895 810 1900
rect 744 1839 749 1895
rect 805 1839 810 1895
rect 744 1834 810 1839
rect 31 1670 91 1834
rect 747 1670 807 1834
rect 28 1665 94 1670
rect 28 1609 33 1665
rect 89 1609 94 1665
rect 28 1604 94 1609
rect 744 1665 810 1670
rect 744 1609 749 1665
rect 805 1609 810 1665
rect 744 1604 810 1609
rect 31 1466 91 1604
rect 747 1466 807 1604
rect 28 1461 94 1466
rect 28 1405 33 1461
rect 89 1405 94 1461
rect 28 1400 94 1405
rect 744 1461 810 1466
rect 744 1405 749 1461
rect 805 1405 810 1461
rect 744 1400 810 1405
rect 31 1262 91 1400
rect 747 1262 807 1400
rect 28 1257 94 1262
rect 28 1201 33 1257
rect 89 1201 94 1257
rect 28 1196 94 1201
rect 744 1257 810 1262
rect 744 1201 749 1257
rect 805 1201 810 1257
rect 744 1196 810 1201
rect 31 1058 91 1196
rect 747 1058 807 1196
rect 28 1053 94 1058
rect 28 997 33 1053
rect 89 997 94 1053
rect 28 992 94 997
rect 744 1053 810 1058
rect 744 997 749 1053
rect 805 997 810 1053
rect 744 992 810 997
rect 31 978 91 992
rect 747 978 807 992
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_0
timestamp 1581321262
transform 1 0 512 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1
timestamp 1581321262
transform 1 0 308 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_2
timestamp 1581321262
transform 1 0 104 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_3
timestamp 1581321262
transform 1 0 308 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_4
timestamp 1581321262
transform 1 0 512 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_5
timestamp 1581321262
transform 1 0 104 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_6
timestamp 1581321262
transform 1 0 512 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_7
timestamp 1581321262
transform 1 0 308 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_8
timestamp 1581321262
transform 1 0 104 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_0
timestamp 1581321262
transform 1 0 512 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1
timestamp 1581321262
transform 1 0 104 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_2
timestamp 1581321262
transform 1 0 308 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_3
timestamp 1581321262
transform 1 0 308 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_4
timestamp 1581321262
transform 1 0 104 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_5
timestamp 1581321262
transform 1 0 512 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_0
timestamp 1581321264
transform 1 0 716 0 1 1485
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_1
timestamp 1581321264
transform 1 0 0 0 1 1485
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_2
timestamp 1581321264
transform 1 0 716 0 1 1281
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_3
timestamp 1581321264
transform 1 0 0 0 1 1281
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_4
timestamp 1581321264
transform 1 0 716 0 1 1077
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_5
timestamp 1581321264
transform 1 0 0 0 1 1077
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_6
timestamp 1581321264
transform 1 0 716 0 1 873
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_7
timestamp 1581321264
transform 1 0 0 0 1 873
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_2  sky130_rom_krom_rom_poly_tap_2_0
timestamp 1581321264
transform 1 0 716 0 1 1689
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_2  sky130_rom_krom_rom_poly_tap_2_1
timestamp 1581321264
transform 1 0 0 0 1 1689
box 0 17 66 83
use sky130_rom_krom_rom_precharge_array_1  sky130_rom_krom_rom_precharge_array_1_0
timestamp 1581321264
transform 1 0 0 0 1 128
box 0 -212 928 408
<< labels >>
rlabel metal2 s 61 368 89 396 4 precharge
port 3 nsew
rlabel metal2 s 19 909 47 937 4 wl_0_0
port 5 nsew
rlabel metal2 s 19 1113 47 1141 4 wl_0_1
port 7 nsew
rlabel metal2 s 19 1317 47 1345 4 wl_0_2
port 9 nsew
rlabel metal2 s 19 1521 47 1549 4 wl_0_3
port 11 nsew
rlabel metal1 s 232 -14 260 14 4 bl_0_0
port 13 nsew
rlabel metal1 s 436 -14 464 14 4 bl_0_1
port 15 nsew
rlabel metal1 s 640 -14 668 14 4 bl_0_2
port 17 nsew
rlabel metal1 s 1017 368 1045 396 4 precharge_r
port 19 nsew
rlabel metal3 s 747 978 807 1038 4 gnd
port 21 nsew
rlabel metal3 s 747 1836 807 1896 4 gnd
port 21 nsew
rlabel metal3 s 31 1836 91 1896 4 gnd
port 21 nsew
rlabel metal3 s 31 978 91 1038 4 gnd
port 21 nsew
rlabel metal2 s 12 -32 40 32 4 vdd
port 23 nsew
<< properties >>
string FIXED_BBOX 0 0 1045 870
<< end >>
