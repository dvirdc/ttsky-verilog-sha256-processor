magic
tech sky130A
magscale 1 2
timestamp 1581585458
<< checkpaint >>
rect -1296 -1289 7004 6546
<< locali >>
rect 2821 5240 2837 5274
rect 2871 5240 2887 5274
rect 64 3997 98 4013
rect 64 3947 98 3963
rect 4443 3925 4477 3959
rect 865 2611 881 2645
rect 915 2611 931 2645
rect 2126 2383 2160 2399
rect 2126 2333 2160 2349
rect 1501 1332 1535 1348
rect 64 1244 98 1310
rect 1501 1282 1535 1298
rect 2008 535 2042 551
rect 2008 485 2042 501
rect 1908 237 1942 303
rect 865 -17 881 17
rect 915 -17 931 17
<< viali >>
rect 2837 5240 2871 5274
rect 64 3963 98 3997
rect 881 2611 915 2645
rect 2126 2349 2160 2383
rect 1501 1298 1535 1332
rect 2008 501 2042 535
rect 881 -17 915 17
<< metal1 >>
rect 2831 5283 2877 5286
rect 2828 5274 2880 5283
rect 2828 5240 2837 5274
rect 2871 5240 2880 5274
rect 2828 5231 2880 5240
rect 2831 5228 2877 5231
rect 52 3997 110 4003
rect 52 3963 64 3997
rect 98 3963 110 3997
rect 52 3957 110 3963
rect 67 3882 95 3957
rect 67 3854 2157 3882
rect 875 2654 921 2657
rect 872 2645 924 2654
rect 872 2611 881 2645
rect 915 2611 924 2645
rect 872 2602 924 2611
rect 875 2599 921 2602
rect 2129 2389 2157 3854
rect 2114 2383 2172 2389
rect 2114 2349 2126 2383
rect 2160 2349 2172 2383
rect 2114 2343 2172 2349
rect 1489 1332 1547 1338
rect 1489 1298 1501 1332
rect 1535 1298 1547 1332
rect 1489 1292 1547 1298
rect 1504 532 1532 1292
rect 1996 535 2054 541
rect 1996 532 2008 535
rect 1504 504 2008 532
rect 1996 501 2008 504
rect 2042 501 2054 535
rect 1996 495 2054 501
rect 875 26 921 29
rect 872 17 924 26
rect 872 -17 881 17
rect 915 -17 924 17
rect 872 -26 924 -17
rect 875 -29 921 -26
use sky130_rom_krom_rom_clock_driver  sky130_rom_krom_rom_clock_driver_0
timestamp 1581585458
transform 1 0 0 0 1 0
box -36 -17 1832 2686
use sky130_rom_krom_rom_control_nand  sky130_rom_krom_rom_control_nand_0
timestamp 1581585458
transform 1 0 1796 0 1 0
box -36 -17 414 2686
use sky130_rom_krom_rom_precharge_driver  sky130_rom_krom_rom_precharge_driver_0
timestamp 1581585458
transform 1 0 0 0 -1 5257
box -36 -17 5744 2686
<< labels >>
rlabel locali s 81 1277 81 1277 4 clk_in
port 2 nsew
rlabel locali s 1518 1315 1518 1315 4 clk_out
port 3 nsew
rlabel locali s 4460 3942 4460 3942 4 prechrg
port 4 nsew
rlabel locali s 1925 270 1925 270 4 CS
port 5 nsew
rlabel metal1 s 872 -26 924 26 4 gnd
port 7 nsew
rlabel metal1 s 2828 5231 2880 5283 4 gnd
port 7 nsew
rlabel metal1 s 872 2602 924 2654 4 vdd
port 9 nsew
<< properties >>
string FIXED_BBOX 865 -29 931 0
<< end >>
