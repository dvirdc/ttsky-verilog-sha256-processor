magic
tech sky130A
magscale 1 2
timestamp 1581365180
<< checkpaint >>
rect -2756 -2756 63334 15012
<< locali >>
rect 7959 11882 7993 11898
rect 7959 11832 7993 11848
rect 7959 11678 7993 11694
rect 7959 11628 7993 11644
rect 7959 11474 7993 11490
rect 7959 11424 7993 11440
rect 7959 11270 7993 11286
rect 7959 11220 7993 11236
rect 7959 11066 7993 11082
rect 7959 11016 7993 11032
rect 7959 10862 7993 10878
rect 7959 10812 7993 10828
rect 7959 10658 7993 10674
rect 7959 10608 7993 10624
rect 7959 10454 7993 10470
rect 7959 10404 7993 10420
rect 8214 9329 8230 9363
rect 8264 9329 8280 9363
rect 8418 9329 8434 9363
rect 8468 9329 8484 9363
rect 8622 9329 8638 9363
rect 8672 9329 8688 9363
rect 8826 9329 8842 9363
rect 8876 9329 8892 9363
rect 9030 9329 9046 9363
rect 9080 9329 9096 9363
rect 9234 9329 9250 9363
rect 9284 9329 9300 9363
rect 9438 9329 9454 9363
rect 9488 9329 9504 9363
rect 9642 9329 9658 9363
rect 9692 9329 9708 9363
rect 9846 9329 9862 9363
rect 9896 9329 9912 9363
rect 10050 9329 10066 9363
rect 10100 9329 10116 9363
rect 10254 9329 10270 9363
rect 10304 9329 10320 9363
rect 10458 9329 10474 9363
rect 10508 9329 10524 9363
rect 10662 9329 10678 9363
rect 10712 9329 10728 9363
rect 10866 9329 10882 9363
rect 10916 9329 10932 9363
rect 11070 9329 11086 9363
rect 11120 9329 11136 9363
rect 11274 9329 11290 9363
rect 11324 9329 11340 9363
rect 11478 9329 11494 9363
rect 11528 9329 11544 9363
rect 11682 9329 11698 9363
rect 11732 9329 11748 9363
rect 11886 9329 11902 9363
rect 11936 9329 11952 9363
rect 12090 9329 12106 9363
rect 12140 9329 12156 9363
rect 12294 9329 12310 9363
rect 12344 9329 12360 9363
rect 12498 9329 12514 9363
rect 12548 9329 12564 9363
rect 12702 9329 12718 9363
rect 12752 9329 12768 9363
rect 12906 9329 12922 9363
rect 12956 9329 12972 9363
rect 13110 9329 13126 9363
rect 13160 9329 13176 9363
rect 13314 9329 13330 9363
rect 13364 9329 13380 9363
rect 13518 9329 13534 9363
rect 13568 9329 13584 9363
rect 13722 9329 13738 9363
rect 13772 9329 13788 9363
rect 13926 9329 13942 9363
rect 13976 9329 13992 9363
rect 14130 9329 14146 9363
rect 14180 9329 14196 9363
rect 14334 9329 14350 9363
rect 14384 9329 14400 9363
rect 14538 9329 14554 9363
rect 14588 9329 14604 9363
rect 14742 9329 14758 9363
rect 14792 9329 14808 9363
rect 14946 9329 14962 9363
rect 14996 9329 15012 9363
rect 15150 9329 15166 9363
rect 15200 9329 15216 9363
rect 15354 9329 15370 9363
rect 15404 9329 15420 9363
rect 15558 9329 15574 9363
rect 15608 9329 15624 9363
rect 15762 9329 15778 9363
rect 15812 9329 15828 9363
rect 15966 9329 15982 9363
rect 16016 9329 16032 9363
rect 16170 9329 16186 9363
rect 16220 9329 16236 9363
rect 16374 9329 16390 9363
rect 16424 9329 16440 9363
rect 16578 9329 16594 9363
rect 16628 9329 16644 9363
rect 16782 9329 16798 9363
rect 16832 9329 16848 9363
rect 16986 9329 17002 9363
rect 17036 9329 17052 9363
rect 17190 9329 17206 9363
rect 17240 9329 17256 9363
rect 17394 9329 17410 9363
rect 17444 9329 17460 9363
rect 17598 9329 17614 9363
rect 17648 9329 17664 9363
rect 17802 9329 17818 9363
rect 17852 9329 17868 9363
rect 18006 9329 18022 9363
rect 18056 9329 18072 9363
rect 18210 9329 18226 9363
rect 18260 9329 18276 9363
rect 18414 9329 18430 9363
rect 18464 9329 18480 9363
rect 18618 9329 18634 9363
rect 18668 9329 18684 9363
rect 18822 9329 18838 9363
rect 18872 9329 18888 9363
rect 19026 9329 19042 9363
rect 19076 9329 19092 9363
rect 19230 9329 19246 9363
rect 19280 9329 19296 9363
rect 19434 9329 19450 9363
rect 19484 9329 19500 9363
rect 19638 9329 19654 9363
rect 19688 9329 19704 9363
rect 19842 9329 19858 9363
rect 19892 9329 19908 9363
rect 20046 9329 20062 9363
rect 20096 9329 20112 9363
rect 20250 9329 20266 9363
rect 20300 9329 20316 9363
rect 20454 9329 20470 9363
rect 20504 9329 20520 9363
rect 20658 9329 20674 9363
rect 20708 9329 20724 9363
rect 20862 9329 20878 9363
rect 20912 9329 20928 9363
rect 21066 9329 21082 9363
rect 21116 9329 21132 9363
rect 21270 9329 21286 9363
rect 21320 9329 21336 9363
rect 21474 9329 21490 9363
rect 21524 9329 21540 9363
rect 21678 9329 21694 9363
rect 21728 9329 21744 9363
rect 21882 9329 21898 9363
rect 21932 9329 21948 9363
rect 22086 9329 22102 9363
rect 22136 9329 22152 9363
rect 22290 9329 22306 9363
rect 22340 9329 22356 9363
rect 22494 9329 22510 9363
rect 22544 9329 22560 9363
rect 22698 9329 22714 9363
rect 22748 9329 22764 9363
rect 22902 9329 22918 9363
rect 22952 9329 22968 9363
rect 23106 9329 23122 9363
rect 23156 9329 23172 9363
rect 23310 9329 23326 9363
rect 23360 9329 23376 9363
rect 23514 9329 23530 9363
rect 23564 9329 23580 9363
rect 23718 9329 23734 9363
rect 23768 9329 23784 9363
rect 23922 9329 23938 9363
rect 23972 9329 23988 9363
rect 24126 9329 24142 9363
rect 24176 9329 24192 9363
rect 24330 9329 24346 9363
rect 24380 9329 24396 9363
rect 24534 9329 24550 9363
rect 24584 9329 24600 9363
rect 24738 9329 24754 9363
rect 24788 9329 24804 9363
rect 24942 9329 24958 9363
rect 24992 9329 25008 9363
rect 25146 9329 25162 9363
rect 25196 9329 25212 9363
rect 25350 9329 25366 9363
rect 25400 9329 25416 9363
rect 25554 9329 25570 9363
rect 25604 9329 25620 9363
rect 25758 9329 25774 9363
rect 25808 9329 25824 9363
rect 25962 9329 25978 9363
rect 26012 9329 26028 9363
rect 26166 9329 26182 9363
rect 26216 9329 26232 9363
rect 26370 9329 26386 9363
rect 26420 9329 26436 9363
rect 26574 9329 26590 9363
rect 26624 9329 26640 9363
rect 26778 9329 26794 9363
rect 26828 9329 26844 9363
rect 26982 9329 26998 9363
rect 27032 9329 27048 9363
rect 27186 9329 27202 9363
rect 27236 9329 27252 9363
rect 27390 9329 27406 9363
rect 27440 9329 27456 9363
rect 27594 9329 27610 9363
rect 27644 9329 27660 9363
rect 27798 9329 27814 9363
rect 27848 9329 27864 9363
rect 28002 9329 28018 9363
rect 28052 9329 28068 9363
rect 28206 9329 28222 9363
rect 28256 9329 28272 9363
rect 28410 9329 28426 9363
rect 28460 9329 28476 9363
rect 28614 9329 28630 9363
rect 28664 9329 28680 9363
rect 28818 9329 28834 9363
rect 28868 9329 28884 9363
rect 29022 9329 29038 9363
rect 29072 9329 29088 9363
rect 29226 9329 29242 9363
rect 29276 9329 29292 9363
rect 29430 9329 29446 9363
rect 29480 9329 29496 9363
rect 29634 9329 29650 9363
rect 29684 9329 29700 9363
rect 29838 9329 29854 9363
rect 29888 9329 29904 9363
rect 30042 9329 30058 9363
rect 30092 9329 30108 9363
rect 30246 9329 30262 9363
rect 30296 9329 30312 9363
rect 30450 9329 30466 9363
rect 30500 9329 30516 9363
rect 30654 9329 30670 9363
rect 30704 9329 30720 9363
rect 30858 9329 30874 9363
rect 30908 9329 30924 9363
rect 31062 9329 31078 9363
rect 31112 9329 31128 9363
rect 31266 9329 31282 9363
rect 31316 9329 31332 9363
rect 31470 9329 31486 9363
rect 31520 9329 31536 9363
rect 31674 9329 31690 9363
rect 31724 9329 31740 9363
rect 31878 9329 31894 9363
rect 31928 9329 31944 9363
rect 32082 9329 32098 9363
rect 32132 9329 32148 9363
rect 32286 9329 32302 9363
rect 32336 9329 32352 9363
rect 32490 9329 32506 9363
rect 32540 9329 32556 9363
rect 32694 9329 32710 9363
rect 32744 9329 32760 9363
rect 32898 9329 32914 9363
rect 32948 9329 32964 9363
rect 33102 9329 33118 9363
rect 33152 9329 33168 9363
rect 33306 9329 33322 9363
rect 33356 9329 33372 9363
rect 33510 9329 33526 9363
rect 33560 9329 33576 9363
rect 33714 9329 33730 9363
rect 33764 9329 33780 9363
rect 33918 9329 33934 9363
rect 33968 9329 33984 9363
rect 34122 9329 34138 9363
rect 34172 9329 34188 9363
rect 34326 9329 34342 9363
rect 34376 9329 34392 9363
rect 34530 9329 34546 9363
rect 34580 9329 34596 9363
rect 34734 9329 34750 9363
rect 34784 9329 34800 9363
rect 34938 9329 34954 9363
rect 34988 9329 35004 9363
rect 35142 9329 35158 9363
rect 35192 9329 35208 9363
rect 35346 9329 35362 9363
rect 35396 9329 35412 9363
rect 35550 9329 35566 9363
rect 35600 9329 35616 9363
rect 35754 9329 35770 9363
rect 35804 9329 35820 9363
rect 35958 9329 35974 9363
rect 36008 9329 36024 9363
rect 36162 9329 36178 9363
rect 36212 9329 36228 9363
rect 36366 9329 36382 9363
rect 36416 9329 36432 9363
rect 36570 9329 36586 9363
rect 36620 9329 36636 9363
rect 36774 9329 36790 9363
rect 36824 9329 36840 9363
rect 36978 9329 36994 9363
rect 37028 9329 37044 9363
rect 37182 9329 37198 9363
rect 37232 9329 37248 9363
rect 37386 9329 37402 9363
rect 37436 9329 37452 9363
rect 37590 9329 37606 9363
rect 37640 9329 37656 9363
rect 37794 9329 37810 9363
rect 37844 9329 37860 9363
rect 37998 9329 38014 9363
rect 38048 9329 38064 9363
rect 38202 9329 38218 9363
rect 38252 9329 38268 9363
rect 38406 9329 38422 9363
rect 38456 9329 38472 9363
rect 38610 9329 38626 9363
rect 38660 9329 38676 9363
rect 38814 9329 38830 9363
rect 38864 9329 38880 9363
rect 39018 9329 39034 9363
rect 39068 9329 39084 9363
rect 39222 9329 39238 9363
rect 39272 9329 39288 9363
rect 39426 9329 39442 9363
rect 39476 9329 39492 9363
rect 39630 9329 39646 9363
rect 39680 9329 39696 9363
rect 39834 9329 39850 9363
rect 39884 9329 39900 9363
rect 40038 9329 40054 9363
rect 40088 9329 40104 9363
rect 40242 9329 40258 9363
rect 40292 9329 40308 9363
rect 40446 9329 40462 9363
rect 40496 9329 40512 9363
rect 40650 9329 40666 9363
rect 40700 9329 40716 9363
rect 40854 9329 40870 9363
rect 40904 9329 40920 9363
rect 41058 9329 41074 9363
rect 41108 9329 41124 9363
rect 41262 9329 41278 9363
rect 41312 9329 41328 9363
rect 41466 9329 41482 9363
rect 41516 9329 41532 9363
rect 41670 9329 41686 9363
rect 41720 9329 41736 9363
rect 41874 9329 41890 9363
rect 41924 9329 41940 9363
rect 42078 9329 42094 9363
rect 42128 9329 42144 9363
rect 42282 9329 42298 9363
rect 42332 9329 42348 9363
rect 42486 9329 42502 9363
rect 42536 9329 42552 9363
rect 42690 9329 42706 9363
rect 42740 9329 42756 9363
rect 42894 9329 42910 9363
rect 42944 9329 42960 9363
rect 43098 9329 43114 9363
rect 43148 9329 43164 9363
rect 43302 9329 43318 9363
rect 43352 9329 43368 9363
rect 43506 9329 43522 9363
rect 43556 9329 43572 9363
rect 43710 9329 43726 9363
rect 43760 9329 43776 9363
rect 43914 9329 43930 9363
rect 43964 9329 43980 9363
rect 44118 9329 44134 9363
rect 44168 9329 44184 9363
rect 44322 9329 44338 9363
rect 44372 9329 44388 9363
rect 44526 9329 44542 9363
rect 44576 9329 44592 9363
rect 44730 9329 44746 9363
rect 44780 9329 44796 9363
rect 44934 9329 44950 9363
rect 44984 9329 45000 9363
rect 45138 9329 45154 9363
rect 45188 9329 45204 9363
rect 45342 9329 45358 9363
rect 45392 9329 45408 9363
rect 45546 9329 45562 9363
rect 45596 9329 45612 9363
rect 45750 9329 45766 9363
rect 45800 9329 45816 9363
rect 45954 9329 45970 9363
rect 46004 9329 46020 9363
rect 46158 9329 46174 9363
rect 46208 9329 46224 9363
rect 46362 9329 46378 9363
rect 46412 9329 46428 9363
rect 46566 9329 46582 9363
rect 46616 9329 46632 9363
rect 46770 9329 46786 9363
rect 46820 9329 46836 9363
rect 46974 9329 46990 9363
rect 47024 9329 47040 9363
rect 47178 9329 47194 9363
rect 47228 9329 47244 9363
rect 47382 9329 47398 9363
rect 47432 9329 47448 9363
rect 47586 9329 47602 9363
rect 47636 9329 47652 9363
rect 47790 9329 47806 9363
rect 47840 9329 47856 9363
rect 47994 9329 48010 9363
rect 48044 9329 48060 9363
rect 48198 9329 48214 9363
rect 48248 9329 48264 9363
rect 48402 9329 48418 9363
rect 48452 9329 48468 9363
rect 48606 9329 48622 9363
rect 48656 9329 48672 9363
rect 48810 9329 48826 9363
rect 48860 9329 48876 9363
rect 49014 9329 49030 9363
rect 49064 9329 49080 9363
rect 49218 9329 49234 9363
rect 49268 9329 49284 9363
rect 49422 9329 49438 9363
rect 49472 9329 49488 9363
rect 49626 9329 49642 9363
rect 49676 9329 49692 9363
rect 49830 9329 49846 9363
rect 49880 9329 49896 9363
rect 50034 9329 50050 9363
rect 50084 9329 50100 9363
rect 50238 9329 50254 9363
rect 50288 9329 50304 9363
rect 50442 9329 50458 9363
rect 50492 9329 50508 9363
rect 50646 9329 50662 9363
rect 50696 9329 50712 9363
rect 50850 9329 50866 9363
rect 50900 9329 50916 9363
rect 51054 9329 51070 9363
rect 51104 9329 51120 9363
rect 51258 9329 51274 9363
rect 51308 9329 51324 9363
rect 51462 9329 51478 9363
rect 51512 9329 51528 9363
rect 51666 9329 51682 9363
rect 51716 9329 51732 9363
rect 51870 9329 51886 9363
rect 51920 9329 51936 9363
rect 52074 9329 52090 9363
rect 52124 9329 52140 9363
rect 52278 9329 52294 9363
rect 52328 9329 52344 9363
rect 52482 9329 52498 9363
rect 52532 9329 52548 9363
rect 52686 9329 52702 9363
rect 52736 9329 52752 9363
rect 52890 9329 52906 9363
rect 52940 9329 52956 9363
rect 53094 9329 53110 9363
rect 53144 9329 53160 9363
rect 53298 9329 53314 9363
rect 53348 9329 53364 9363
rect 53502 9329 53518 9363
rect 53552 9329 53568 9363
rect 53706 9329 53722 9363
rect 53756 9329 53772 9363
rect 53910 9329 53926 9363
rect 53960 9329 53976 9363
rect 54114 9329 54130 9363
rect 54164 9329 54180 9363
rect 54318 9329 54334 9363
rect 54368 9329 54384 9363
rect 54522 9329 54538 9363
rect 54572 9329 54588 9363
rect 54726 9329 54742 9363
rect 54776 9329 54792 9363
rect 54930 9329 54946 9363
rect 54980 9329 54996 9363
rect 55134 9329 55150 9363
rect 55184 9329 55200 9363
rect 55338 9329 55354 9363
rect 55388 9329 55404 9363
rect 55542 9329 55558 9363
rect 55592 9329 55608 9363
rect 55746 9329 55762 9363
rect 55796 9329 55812 9363
rect 55950 9329 55966 9363
rect 56000 9329 56016 9363
rect 56154 9329 56170 9363
rect 56204 9329 56220 9363
rect 56358 9329 56374 9363
rect 56408 9329 56424 9363
rect 56562 9329 56578 9363
rect 56612 9329 56628 9363
rect 56766 9329 56782 9363
rect 56816 9329 56832 9363
rect 56970 9329 56986 9363
rect 57020 9329 57036 9363
rect 57174 9329 57190 9363
rect 57224 9329 57240 9363
rect 57378 9329 57394 9363
rect 57428 9329 57444 9363
rect 57582 9329 57598 9363
rect 57632 9329 57648 9363
rect 57786 9329 57802 9363
rect 57836 9329 57852 9363
rect 57990 9329 58006 9363
rect 58040 9329 58056 9363
rect 58194 9329 58210 9363
rect 58244 9329 58260 9363
rect 58398 9329 58414 9363
rect 58448 9329 58464 9363
rect 58602 9329 58618 9363
rect 58652 9329 58668 9363
rect 58806 9329 58822 9363
rect 58856 9329 58872 9363
rect 59010 9329 59026 9363
rect 59060 9329 59076 9363
rect 59214 9329 59230 9363
rect 59264 9329 59280 9363
rect 59418 9329 59434 9363
rect 59468 9329 59484 9363
rect 59622 9329 59638 9363
rect 59672 9329 59688 9363
rect 59826 9329 59842 9363
rect 59876 9329 59892 9363
rect 60030 9329 60046 9363
rect 60080 9329 60096 9363
rect 60234 9329 60250 9363
rect 60284 9329 60300 9363
rect 8214 7734 8230 7768
rect 8264 7734 8280 7768
rect 8418 7734 8434 7768
rect 8468 7734 8484 7768
rect 8622 7734 8638 7768
rect 8672 7734 8688 7768
rect 8826 7734 8842 7768
rect 8876 7734 8892 7768
rect 9030 7734 9046 7768
rect 9080 7734 9096 7768
rect 9234 7734 9250 7768
rect 9284 7734 9300 7768
rect 9438 7734 9454 7768
rect 9488 7734 9504 7768
rect 9642 7734 9658 7768
rect 9692 7734 9708 7768
rect 9846 7734 9862 7768
rect 9896 7734 9912 7768
rect 10050 7734 10066 7768
rect 10100 7734 10116 7768
rect 10254 7734 10270 7768
rect 10304 7734 10320 7768
rect 10458 7734 10474 7768
rect 10508 7734 10524 7768
rect 10662 7734 10678 7768
rect 10712 7734 10728 7768
rect 10866 7734 10882 7768
rect 10916 7734 10932 7768
rect 11070 7734 11086 7768
rect 11120 7734 11136 7768
rect 11274 7734 11290 7768
rect 11324 7734 11340 7768
rect 11478 7734 11494 7768
rect 11528 7734 11544 7768
rect 11682 7734 11698 7768
rect 11732 7734 11748 7768
rect 11886 7734 11902 7768
rect 11936 7734 11952 7768
rect 12090 7734 12106 7768
rect 12140 7734 12156 7768
rect 12294 7734 12310 7768
rect 12344 7734 12360 7768
rect 12498 7734 12514 7768
rect 12548 7734 12564 7768
rect 12702 7734 12718 7768
rect 12752 7734 12768 7768
rect 12906 7734 12922 7768
rect 12956 7734 12972 7768
rect 13110 7734 13126 7768
rect 13160 7734 13176 7768
rect 13314 7734 13330 7768
rect 13364 7734 13380 7768
rect 13518 7734 13534 7768
rect 13568 7734 13584 7768
rect 13722 7734 13738 7768
rect 13772 7734 13788 7768
rect 13926 7734 13942 7768
rect 13976 7734 13992 7768
rect 14130 7734 14146 7768
rect 14180 7734 14196 7768
rect 14334 7734 14350 7768
rect 14384 7734 14400 7768
rect 14538 7734 14554 7768
rect 14588 7734 14604 7768
rect 14742 7734 14758 7768
rect 14792 7734 14808 7768
rect 14946 7734 14962 7768
rect 14996 7734 15012 7768
rect 15150 7734 15166 7768
rect 15200 7734 15216 7768
rect 15354 7734 15370 7768
rect 15404 7734 15420 7768
rect 15558 7734 15574 7768
rect 15608 7734 15624 7768
rect 15762 7734 15778 7768
rect 15812 7734 15828 7768
rect 15966 7734 15982 7768
rect 16016 7734 16032 7768
rect 16170 7734 16186 7768
rect 16220 7734 16236 7768
rect 16374 7734 16390 7768
rect 16424 7734 16440 7768
rect 16578 7734 16594 7768
rect 16628 7734 16644 7768
rect 16782 7734 16798 7768
rect 16832 7734 16848 7768
rect 16986 7734 17002 7768
rect 17036 7734 17052 7768
rect 17190 7734 17206 7768
rect 17240 7734 17256 7768
rect 17394 7734 17410 7768
rect 17444 7734 17460 7768
rect 17598 7734 17614 7768
rect 17648 7734 17664 7768
rect 17802 7734 17818 7768
rect 17852 7734 17868 7768
rect 18006 7734 18022 7768
rect 18056 7734 18072 7768
rect 18210 7734 18226 7768
rect 18260 7734 18276 7768
rect 18414 7734 18430 7768
rect 18464 7734 18480 7768
rect 18618 7734 18634 7768
rect 18668 7734 18684 7768
rect 18822 7734 18838 7768
rect 18872 7734 18888 7768
rect 19026 7734 19042 7768
rect 19076 7734 19092 7768
rect 19230 7734 19246 7768
rect 19280 7734 19296 7768
rect 19434 7734 19450 7768
rect 19484 7734 19500 7768
rect 19638 7734 19654 7768
rect 19688 7734 19704 7768
rect 19842 7734 19858 7768
rect 19892 7734 19908 7768
rect 20046 7734 20062 7768
rect 20096 7734 20112 7768
rect 20250 7734 20266 7768
rect 20300 7734 20316 7768
rect 20454 7734 20470 7768
rect 20504 7734 20520 7768
rect 20658 7734 20674 7768
rect 20708 7734 20724 7768
rect 20862 7734 20878 7768
rect 20912 7734 20928 7768
rect 21066 7734 21082 7768
rect 21116 7734 21132 7768
rect 21270 7734 21286 7768
rect 21320 7734 21336 7768
rect 21474 7734 21490 7768
rect 21524 7734 21540 7768
rect 21678 7734 21694 7768
rect 21728 7734 21744 7768
rect 21882 7734 21898 7768
rect 21932 7734 21948 7768
rect 22086 7734 22102 7768
rect 22136 7734 22152 7768
rect 22290 7734 22306 7768
rect 22340 7734 22356 7768
rect 22494 7734 22510 7768
rect 22544 7734 22560 7768
rect 22698 7734 22714 7768
rect 22748 7734 22764 7768
rect 22902 7734 22918 7768
rect 22952 7734 22968 7768
rect 23106 7734 23122 7768
rect 23156 7734 23172 7768
rect 23310 7734 23326 7768
rect 23360 7734 23376 7768
rect 23514 7734 23530 7768
rect 23564 7734 23580 7768
rect 23718 7734 23734 7768
rect 23768 7734 23784 7768
rect 23922 7734 23938 7768
rect 23972 7734 23988 7768
rect 24126 7734 24142 7768
rect 24176 7734 24192 7768
rect 24330 7734 24346 7768
rect 24380 7734 24396 7768
rect 24534 7734 24550 7768
rect 24584 7734 24600 7768
rect 24738 7734 24754 7768
rect 24788 7734 24804 7768
rect 24942 7734 24958 7768
rect 24992 7734 25008 7768
rect 25146 7734 25162 7768
rect 25196 7734 25212 7768
rect 25350 7734 25366 7768
rect 25400 7734 25416 7768
rect 25554 7734 25570 7768
rect 25604 7734 25620 7768
rect 25758 7734 25774 7768
rect 25808 7734 25824 7768
rect 25962 7734 25978 7768
rect 26012 7734 26028 7768
rect 26166 7734 26182 7768
rect 26216 7734 26232 7768
rect 26370 7734 26386 7768
rect 26420 7734 26436 7768
rect 26574 7734 26590 7768
rect 26624 7734 26640 7768
rect 26778 7734 26794 7768
rect 26828 7734 26844 7768
rect 26982 7734 26998 7768
rect 27032 7734 27048 7768
rect 27186 7734 27202 7768
rect 27236 7734 27252 7768
rect 27390 7734 27406 7768
rect 27440 7734 27456 7768
rect 27594 7734 27610 7768
rect 27644 7734 27660 7768
rect 27798 7734 27814 7768
rect 27848 7734 27864 7768
rect 28002 7734 28018 7768
rect 28052 7734 28068 7768
rect 28206 7734 28222 7768
rect 28256 7734 28272 7768
rect 28410 7734 28426 7768
rect 28460 7734 28476 7768
rect 28614 7734 28630 7768
rect 28664 7734 28680 7768
rect 28818 7734 28834 7768
rect 28868 7734 28884 7768
rect 29022 7734 29038 7768
rect 29072 7734 29088 7768
rect 29226 7734 29242 7768
rect 29276 7734 29292 7768
rect 29430 7734 29446 7768
rect 29480 7734 29496 7768
rect 29634 7734 29650 7768
rect 29684 7734 29700 7768
rect 29838 7734 29854 7768
rect 29888 7734 29904 7768
rect 30042 7734 30058 7768
rect 30092 7734 30108 7768
rect 30246 7734 30262 7768
rect 30296 7734 30312 7768
rect 30450 7734 30466 7768
rect 30500 7734 30516 7768
rect 30654 7734 30670 7768
rect 30704 7734 30720 7768
rect 30858 7734 30874 7768
rect 30908 7734 30924 7768
rect 31062 7734 31078 7768
rect 31112 7734 31128 7768
rect 31266 7734 31282 7768
rect 31316 7734 31332 7768
rect 31470 7734 31486 7768
rect 31520 7734 31536 7768
rect 31674 7734 31690 7768
rect 31724 7734 31740 7768
rect 31878 7734 31894 7768
rect 31928 7734 31944 7768
rect 32082 7734 32098 7768
rect 32132 7734 32148 7768
rect 32286 7734 32302 7768
rect 32336 7734 32352 7768
rect 32490 7734 32506 7768
rect 32540 7734 32556 7768
rect 32694 7734 32710 7768
rect 32744 7734 32760 7768
rect 32898 7734 32914 7768
rect 32948 7734 32964 7768
rect 33102 7734 33118 7768
rect 33152 7734 33168 7768
rect 33306 7734 33322 7768
rect 33356 7734 33372 7768
rect 33510 7734 33526 7768
rect 33560 7734 33576 7768
rect 33714 7734 33730 7768
rect 33764 7734 33780 7768
rect 33918 7734 33934 7768
rect 33968 7734 33984 7768
rect 34122 7734 34138 7768
rect 34172 7734 34188 7768
rect 34326 7734 34342 7768
rect 34376 7734 34392 7768
rect 34530 7734 34546 7768
rect 34580 7734 34596 7768
rect 34734 7734 34750 7768
rect 34784 7734 34800 7768
rect 34938 7734 34954 7768
rect 34988 7734 35004 7768
rect 35142 7734 35158 7768
rect 35192 7734 35208 7768
rect 35346 7734 35362 7768
rect 35396 7734 35412 7768
rect 35550 7734 35566 7768
rect 35600 7734 35616 7768
rect 35754 7734 35770 7768
rect 35804 7734 35820 7768
rect 35958 7734 35974 7768
rect 36008 7734 36024 7768
rect 36162 7734 36178 7768
rect 36212 7734 36228 7768
rect 36366 7734 36382 7768
rect 36416 7734 36432 7768
rect 36570 7734 36586 7768
rect 36620 7734 36636 7768
rect 36774 7734 36790 7768
rect 36824 7734 36840 7768
rect 36978 7734 36994 7768
rect 37028 7734 37044 7768
rect 37182 7734 37198 7768
rect 37232 7734 37248 7768
rect 37386 7734 37402 7768
rect 37436 7734 37452 7768
rect 37590 7734 37606 7768
rect 37640 7734 37656 7768
rect 37794 7734 37810 7768
rect 37844 7734 37860 7768
rect 37998 7734 38014 7768
rect 38048 7734 38064 7768
rect 38202 7734 38218 7768
rect 38252 7734 38268 7768
rect 38406 7734 38422 7768
rect 38456 7734 38472 7768
rect 38610 7734 38626 7768
rect 38660 7734 38676 7768
rect 38814 7734 38830 7768
rect 38864 7734 38880 7768
rect 39018 7734 39034 7768
rect 39068 7734 39084 7768
rect 39222 7734 39238 7768
rect 39272 7734 39288 7768
rect 39426 7734 39442 7768
rect 39476 7734 39492 7768
rect 39630 7734 39646 7768
rect 39680 7734 39696 7768
rect 39834 7734 39850 7768
rect 39884 7734 39900 7768
rect 40038 7734 40054 7768
rect 40088 7734 40104 7768
rect 40242 7734 40258 7768
rect 40292 7734 40308 7768
rect 40446 7734 40462 7768
rect 40496 7734 40512 7768
rect 40650 7734 40666 7768
rect 40700 7734 40716 7768
rect 40854 7734 40870 7768
rect 40904 7734 40920 7768
rect 41058 7734 41074 7768
rect 41108 7734 41124 7768
rect 41262 7734 41278 7768
rect 41312 7734 41328 7768
rect 41466 7734 41482 7768
rect 41516 7734 41532 7768
rect 41670 7734 41686 7768
rect 41720 7734 41736 7768
rect 41874 7734 41890 7768
rect 41924 7734 41940 7768
rect 42078 7734 42094 7768
rect 42128 7734 42144 7768
rect 42282 7734 42298 7768
rect 42332 7734 42348 7768
rect 42486 7734 42502 7768
rect 42536 7734 42552 7768
rect 42690 7734 42706 7768
rect 42740 7734 42756 7768
rect 42894 7734 42910 7768
rect 42944 7734 42960 7768
rect 43098 7734 43114 7768
rect 43148 7734 43164 7768
rect 43302 7734 43318 7768
rect 43352 7734 43368 7768
rect 43506 7734 43522 7768
rect 43556 7734 43572 7768
rect 43710 7734 43726 7768
rect 43760 7734 43776 7768
rect 43914 7734 43930 7768
rect 43964 7734 43980 7768
rect 44118 7734 44134 7768
rect 44168 7734 44184 7768
rect 44322 7734 44338 7768
rect 44372 7734 44388 7768
rect 44526 7734 44542 7768
rect 44576 7734 44592 7768
rect 44730 7734 44746 7768
rect 44780 7734 44796 7768
rect 44934 7734 44950 7768
rect 44984 7734 45000 7768
rect 45138 7734 45154 7768
rect 45188 7734 45204 7768
rect 45342 7734 45358 7768
rect 45392 7734 45408 7768
rect 45546 7734 45562 7768
rect 45596 7734 45612 7768
rect 45750 7734 45766 7768
rect 45800 7734 45816 7768
rect 45954 7734 45970 7768
rect 46004 7734 46020 7768
rect 46158 7734 46174 7768
rect 46208 7734 46224 7768
rect 46362 7734 46378 7768
rect 46412 7734 46428 7768
rect 46566 7734 46582 7768
rect 46616 7734 46632 7768
rect 46770 7734 46786 7768
rect 46820 7734 46836 7768
rect 46974 7734 46990 7768
rect 47024 7734 47040 7768
rect 47178 7734 47194 7768
rect 47228 7734 47244 7768
rect 47382 7734 47398 7768
rect 47432 7734 47448 7768
rect 47586 7734 47602 7768
rect 47636 7734 47652 7768
rect 47790 7734 47806 7768
rect 47840 7734 47856 7768
rect 47994 7734 48010 7768
rect 48044 7734 48060 7768
rect 48198 7734 48214 7768
rect 48248 7734 48264 7768
rect 48402 7734 48418 7768
rect 48452 7734 48468 7768
rect 48606 7734 48622 7768
rect 48656 7734 48672 7768
rect 48810 7734 48826 7768
rect 48860 7734 48876 7768
rect 49014 7734 49030 7768
rect 49064 7734 49080 7768
rect 49218 7734 49234 7768
rect 49268 7734 49284 7768
rect 49422 7734 49438 7768
rect 49472 7734 49488 7768
rect 49626 7734 49642 7768
rect 49676 7734 49692 7768
rect 49830 7734 49846 7768
rect 49880 7734 49896 7768
rect 50034 7734 50050 7768
rect 50084 7734 50100 7768
rect 50238 7734 50254 7768
rect 50288 7734 50304 7768
rect 50442 7734 50458 7768
rect 50492 7734 50508 7768
rect 50646 7734 50662 7768
rect 50696 7734 50712 7768
rect 50850 7734 50866 7768
rect 50900 7734 50916 7768
rect 51054 7734 51070 7768
rect 51104 7734 51120 7768
rect 51258 7734 51274 7768
rect 51308 7734 51324 7768
rect 51462 7734 51478 7768
rect 51512 7734 51528 7768
rect 51666 7734 51682 7768
rect 51716 7734 51732 7768
rect 51870 7734 51886 7768
rect 51920 7734 51936 7768
rect 52074 7734 52090 7768
rect 52124 7734 52140 7768
rect 52278 7734 52294 7768
rect 52328 7734 52344 7768
rect 52482 7734 52498 7768
rect 52532 7734 52548 7768
rect 52686 7734 52702 7768
rect 52736 7734 52752 7768
rect 52890 7734 52906 7768
rect 52940 7734 52956 7768
rect 53094 7734 53110 7768
rect 53144 7734 53160 7768
rect 53298 7734 53314 7768
rect 53348 7734 53364 7768
rect 53502 7734 53518 7768
rect 53552 7734 53568 7768
rect 53706 7734 53722 7768
rect 53756 7734 53772 7768
rect 53910 7734 53926 7768
rect 53960 7734 53976 7768
rect 54114 7734 54130 7768
rect 54164 7734 54180 7768
rect 54318 7734 54334 7768
rect 54368 7734 54384 7768
rect 54522 7734 54538 7768
rect 54572 7734 54588 7768
rect 54726 7734 54742 7768
rect 54776 7734 54792 7768
rect 54930 7734 54946 7768
rect 54980 7734 54996 7768
rect 55134 7734 55150 7768
rect 55184 7734 55200 7768
rect 55338 7734 55354 7768
rect 55388 7734 55404 7768
rect 55542 7734 55558 7768
rect 55592 7734 55608 7768
rect 55746 7734 55762 7768
rect 55796 7734 55812 7768
rect 55950 7734 55966 7768
rect 56000 7734 56016 7768
rect 56154 7734 56170 7768
rect 56204 7734 56220 7768
rect 56358 7734 56374 7768
rect 56408 7734 56424 7768
rect 56562 7734 56578 7768
rect 56612 7734 56628 7768
rect 56766 7734 56782 7768
rect 56816 7734 56832 7768
rect 56970 7734 56986 7768
rect 57020 7734 57036 7768
rect 57174 7734 57190 7768
rect 57224 7734 57240 7768
rect 57378 7734 57394 7768
rect 57428 7734 57444 7768
rect 57582 7734 57598 7768
rect 57632 7734 57648 7768
rect 57786 7734 57802 7768
rect 57836 7734 57852 7768
rect 57990 7734 58006 7768
rect 58040 7734 58056 7768
rect 58194 7734 58210 7768
rect 58244 7734 58260 7768
rect 58398 7734 58414 7768
rect 58448 7734 58464 7768
rect 58602 7734 58618 7768
rect 58652 7734 58668 7768
rect 58806 7734 58822 7768
rect 58856 7734 58872 7768
rect 59010 7734 59026 7768
rect 59060 7734 59076 7768
rect 59214 7734 59230 7768
rect 59264 7734 59280 7768
rect 59418 7734 59434 7768
rect 59468 7734 59484 7768
rect 59622 7734 59638 7768
rect 59672 7734 59688 7768
rect 59826 7734 59842 7768
rect 59876 7734 59892 7768
rect 60030 7734 60046 7768
rect 60080 7734 60096 7768
rect 60234 7734 60250 7768
rect 60284 7734 60300 7768
rect 337 7093 371 7109
rect 337 7043 371 7059
rect 745 7093 779 7109
rect 745 7043 779 7059
rect 1153 7093 1187 7109
rect 1153 7043 1187 7059
rect 7959 6413 7993 6429
rect 7959 6363 7993 6379
rect 7959 6209 7993 6225
rect 7959 6159 7993 6175
rect 7959 6005 7993 6021
rect 7959 5955 7993 5971
rect 7959 5801 7993 5817
rect 7959 5751 7993 5767
rect 2993 5622 3027 5638
rect 2993 5572 3027 5588
rect 7959 5597 7993 5613
rect 7959 5547 7993 5563
rect 7959 5393 7993 5409
rect 7959 5343 7993 5359
rect 7959 5189 7993 5205
rect 7959 5139 7993 5155
rect 7959 4985 7993 5001
rect 7959 4935 7993 4951
rect 51 2995 85 3011
rect -1386 2957 -1352 2973
rect 51 2945 85 2961
rect -1386 2907 -1352 2923
rect 458 1950 492 1966
rect 458 1900 492 1916
rect 14692 1739 14726 1755
rect 14692 1689 14726 1705
rect 15000 1739 15034 1755
rect 15000 1689 15034 1705
rect 15308 1739 15342 1755
rect 15308 1689 15342 1705
rect 15616 1739 15650 1755
rect 15616 1689 15650 1705
rect 15924 1739 15958 1755
rect 15924 1689 15958 1705
rect 16232 1739 16266 1755
rect 16232 1689 16266 1705
rect 16540 1739 16574 1755
rect 16540 1689 16574 1705
rect 16848 1739 16882 1755
rect 16848 1689 16882 1705
rect 17156 1739 17190 1755
rect 17156 1689 17190 1705
rect 17464 1739 17498 1755
rect 17464 1689 17498 1705
rect 17772 1739 17806 1755
rect 17772 1689 17806 1705
rect 18080 1739 18114 1755
rect 18080 1689 18114 1705
rect 18388 1739 18422 1755
rect 18388 1689 18422 1705
rect 18696 1739 18730 1755
rect 18696 1689 18730 1705
rect 19004 1739 19038 1755
rect 19004 1689 19038 1705
rect 19312 1739 19346 1755
rect 19312 1689 19346 1705
rect 19620 1739 19654 1755
rect 19620 1689 19654 1705
rect 19928 1739 19962 1755
rect 19928 1689 19962 1705
rect 20236 1739 20270 1755
rect 20236 1689 20270 1705
rect 20544 1739 20578 1755
rect 20544 1689 20578 1705
rect 20852 1739 20886 1755
rect 20852 1689 20886 1705
rect 21160 1739 21194 1755
rect 21160 1689 21194 1705
rect 21468 1739 21502 1755
rect 21468 1689 21502 1705
rect 21776 1739 21810 1755
rect 21776 1689 21810 1705
rect 22084 1739 22118 1755
rect 22084 1689 22118 1705
rect 22392 1739 22426 1755
rect 22392 1689 22426 1705
rect 22700 1739 22734 1755
rect 22700 1689 22734 1705
rect 23008 1739 23042 1755
rect 23008 1689 23042 1705
rect 23316 1739 23350 1755
rect 23316 1689 23350 1705
rect 23624 1739 23658 1755
rect 23624 1689 23658 1705
rect 23932 1739 23966 1755
rect 23932 1689 23966 1705
rect 24240 1739 24274 1755
rect 24240 1689 24274 1705
rect 4835 1624 4869 1640
rect 4835 1574 4869 1590
rect 5243 1624 5277 1640
rect 5243 1574 5277 1590
rect 5651 1624 5685 1640
rect 5651 1574 5685 1590
rect 14676 0 14692 34
rect 14726 0 14742 34
rect 14984 0 15000 34
rect 15034 0 15050 34
rect 15292 0 15308 34
rect 15342 0 15358 34
rect 15600 0 15616 34
rect 15650 0 15666 34
rect 15908 0 15924 34
rect 15958 0 15974 34
rect 16216 0 16232 34
rect 16266 0 16282 34
rect 16524 0 16540 34
rect 16574 0 16590 34
rect 16832 0 16848 34
rect 16882 0 16898 34
rect 17140 0 17156 34
rect 17190 0 17206 34
rect 17448 0 17464 34
rect 17498 0 17514 34
rect 17756 0 17772 34
rect 17806 0 17822 34
rect 18064 0 18080 34
rect 18114 0 18130 34
rect 18372 0 18388 34
rect 18422 0 18438 34
rect 18680 0 18696 34
rect 18730 0 18746 34
rect 18988 0 19004 34
rect 19038 0 19054 34
rect 19296 0 19312 34
rect 19346 0 19362 34
rect 19604 0 19620 34
rect 19654 0 19670 34
rect 19912 0 19928 34
rect 19962 0 19978 34
rect 20220 0 20236 34
rect 20270 0 20286 34
rect 20528 0 20544 34
rect 20578 0 20594 34
rect 20836 0 20852 34
rect 20886 0 20902 34
rect 21144 0 21160 34
rect 21194 0 21210 34
rect 21452 0 21468 34
rect 21502 0 21518 34
rect 21760 0 21776 34
rect 21810 0 21826 34
rect 22068 0 22084 34
rect 22118 0 22134 34
rect 22376 0 22392 34
rect 22426 0 22442 34
rect 22684 0 22700 34
rect 22734 0 22750 34
rect 22992 0 23008 34
rect 23042 0 23058 34
rect 23300 0 23316 34
rect 23350 0 23366 34
rect 23608 0 23624 34
rect 23658 0 23674 34
rect 23916 0 23932 34
rect 23966 0 23982 34
rect 24224 0 24240 34
rect 24274 0 24290 34
<< viali >>
rect 7959 11848 7993 11882
rect 7959 11644 7993 11678
rect 7959 11440 7993 11474
rect 7959 11236 7993 11270
rect 7959 11032 7993 11066
rect 7959 10828 7993 10862
rect 7959 10624 7993 10658
rect 7959 10420 7993 10454
rect 8230 9329 8264 9363
rect 8434 9329 8468 9363
rect 8638 9329 8672 9363
rect 8842 9329 8876 9363
rect 9046 9329 9080 9363
rect 9250 9329 9284 9363
rect 9454 9329 9488 9363
rect 9658 9329 9692 9363
rect 9862 9329 9896 9363
rect 10066 9329 10100 9363
rect 10270 9329 10304 9363
rect 10474 9329 10508 9363
rect 10678 9329 10712 9363
rect 10882 9329 10916 9363
rect 11086 9329 11120 9363
rect 11290 9329 11324 9363
rect 11494 9329 11528 9363
rect 11698 9329 11732 9363
rect 11902 9329 11936 9363
rect 12106 9329 12140 9363
rect 12310 9329 12344 9363
rect 12514 9329 12548 9363
rect 12718 9329 12752 9363
rect 12922 9329 12956 9363
rect 13126 9329 13160 9363
rect 13330 9329 13364 9363
rect 13534 9329 13568 9363
rect 13738 9329 13772 9363
rect 13942 9329 13976 9363
rect 14146 9329 14180 9363
rect 14350 9329 14384 9363
rect 14554 9329 14588 9363
rect 14758 9329 14792 9363
rect 14962 9329 14996 9363
rect 15166 9329 15200 9363
rect 15370 9329 15404 9363
rect 15574 9329 15608 9363
rect 15778 9329 15812 9363
rect 15982 9329 16016 9363
rect 16186 9329 16220 9363
rect 16390 9329 16424 9363
rect 16594 9329 16628 9363
rect 16798 9329 16832 9363
rect 17002 9329 17036 9363
rect 17206 9329 17240 9363
rect 17410 9329 17444 9363
rect 17614 9329 17648 9363
rect 17818 9329 17852 9363
rect 18022 9329 18056 9363
rect 18226 9329 18260 9363
rect 18430 9329 18464 9363
rect 18634 9329 18668 9363
rect 18838 9329 18872 9363
rect 19042 9329 19076 9363
rect 19246 9329 19280 9363
rect 19450 9329 19484 9363
rect 19654 9329 19688 9363
rect 19858 9329 19892 9363
rect 20062 9329 20096 9363
rect 20266 9329 20300 9363
rect 20470 9329 20504 9363
rect 20674 9329 20708 9363
rect 20878 9329 20912 9363
rect 21082 9329 21116 9363
rect 21286 9329 21320 9363
rect 21490 9329 21524 9363
rect 21694 9329 21728 9363
rect 21898 9329 21932 9363
rect 22102 9329 22136 9363
rect 22306 9329 22340 9363
rect 22510 9329 22544 9363
rect 22714 9329 22748 9363
rect 22918 9329 22952 9363
rect 23122 9329 23156 9363
rect 23326 9329 23360 9363
rect 23530 9329 23564 9363
rect 23734 9329 23768 9363
rect 23938 9329 23972 9363
rect 24142 9329 24176 9363
rect 24346 9329 24380 9363
rect 24550 9329 24584 9363
rect 24754 9329 24788 9363
rect 24958 9329 24992 9363
rect 25162 9329 25196 9363
rect 25366 9329 25400 9363
rect 25570 9329 25604 9363
rect 25774 9329 25808 9363
rect 25978 9329 26012 9363
rect 26182 9329 26216 9363
rect 26386 9329 26420 9363
rect 26590 9329 26624 9363
rect 26794 9329 26828 9363
rect 26998 9329 27032 9363
rect 27202 9329 27236 9363
rect 27406 9329 27440 9363
rect 27610 9329 27644 9363
rect 27814 9329 27848 9363
rect 28018 9329 28052 9363
rect 28222 9329 28256 9363
rect 28426 9329 28460 9363
rect 28630 9329 28664 9363
rect 28834 9329 28868 9363
rect 29038 9329 29072 9363
rect 29242 9329 29276 9363
rect 29446 9329 29480 9363
rect 29650 9329 29684 9363
rect 29854 9329 29888 9363
rect 30058 9329 30092 9363
rect 30262 9329 30296 9363
rect 30466 9329 30500 9363
rect 30670 9329 30704 9363
rect 30874 9329 30908 9363
rect 31078 9329 31112 9363
rect 31282 9329 31316 9363
rect 31486 9329 31520 9363
rect 31690 9329 31724 9363
rect 31894 9329 31928 9363
rect 32098 9329 32132 9363
rect 32302 9329 32336 9363
rect 32506 9329 32540 9363
rect 32710 9329 32744 9363
rect 32914 9329 32948 9363
rect 33118 9329 33152 9363
rect 33322 9329 33356 9363
rect 33526 9329 33560 9363
rect 33730 9329 33764 9363
rect 33934 9329 33968 9363
rect 34138 9329 34172 9363
rect 34342 9329 34376 9363
rect 34546 9329 34580 9363
rect 34750 9329 34784 9363
rect 34954 9329 34988 9363
rect 35158 9329 35192 9363
rect 35362 9329 35396 9363
rect 35566 9329 35600 9363
rect 35770 9329 35804 9363
rect 35974 9329 36008 9363
rect 36178 9329 36212 9363
rect 36382 9329 36416 9363
rect 36586 9329 36620 9363
rect 36790 9329 36824 9363
rect 36994 9329 37028 9363
rect 37198 9329 37232 9363
rect 37402 9329 37436 9363
rect 37606 9329 37640 9363
rect 37810 9329 37844 9363
rect 38014 9329 38048 9363
rect 38218 9329 38252 9363
rect 38422 9329 38456 9363
rect 38626 9329 38660 9363
rect 38830 9329 38864 9363
rect 39034 9329 39068 9363
rect 39238 9329 39272 9363
rect 39442 9329 39476 9363
rect 39646 9329 39680 9363
rect 39850 9329 39884 9363
rect 40054 9329 40088 9363
rect 40258 9329 40292 9363
rect 40462 9329 40496 9363
rect 40666 9329 40700 9363
rect 40870 9329 40904 9363
rect 41074 9329 41108 9363
rect 41278 9329 41312 9363
rect 41482 9329 41516 9363
rect 41686 9329 41720 9363
rect 41890 9329 41924 9363
rect 42094 9329 42128 9363
rect 42298 9329 42332 9363
rect 42502 9329 42536 9363
rect 42706 9329 42740 9363
rect 42910 9329 42944 9363
rect 43114 9329 43148 9363
rect 43318 9329 43352 9363
rect 43522 9329 43556 9363
rect 43726 9329 43760 9363
rect 43930 9329 43964 9363
rect 44134 9329 44168 9363
rect 44338 9329 44372 9363
rect 44542 9329 44576 9363
rect 44746 9329 44780 9363
rect 44950 9329 44984 9363
rect 45154 9329 45188 9363
rect 45358 9329 45392 9363
rect 45562 9329 45596 9363
rect 45766 9329 45800 9363
rect 45970 9329 46004 9363
rect 46174 9329 46208 9363
rect 46378 9329 46412 9363
rect 46582 9329 46616 9363
rect 46786 9329 46820 9363
rect 46990 9329 47024 9363
rect 47194 9329 47228 9363
rect 47398 9329 47432 9363
rect 47602 9329 47636 9363
rect 47806 9329 47840 9363
rect 48010 9329 48044 9363
rect 48214 9329 48248 9363
rect 48418 9329 48452 9363
rect 48622 9329 48656 9363
rect 48826 9329 48860 9363
rect 49030 9329 49064 9363
rect 49234 9329 49268 9363
rect 49438 9329 49472 9363
rect 49642 9329 49676 9363
rect 49846 9329 49880 9363
rect 50050 9329 50084 9363
rect 50254 9329 50288 9363
rect 50458 9329 50492 9363
rect 50662 9329 50696 9363
rect 50866 9329 50900 9363
rect 51070 9329 51104 9363
rect 51274 9329 51308 9363
rect 51478 9329 51512 9363
rect 51682 9329 51716 9363
rect 51886 9329 51920 9363
rect 52090 9329 52124 9363
rect 52294 9329 52328 9363
rect 52498 9329 52532 9363
rect 52702 9329 52736 9363
rect 52906 9329 52940 9363
rect 53110 9329 53144 9363
rect 53314 9329 53348 9363
rect 53518 9329 53552 9363
rect 53722 9329 53756 9363
rect 53926 9329 53960 9363
rect 54130 9329 54164 9363
rect 54334 9329 54368 9363
rect 54538 9329 54572 9363
rect 54742 9329 54776 9363
rect 54946 9329 54980 9363
rect 55150 9329 55184 9363
rect 55354 9329 55388 9363
rect 55558 9329 55592 9363
rect 55762 9329 55796 9363
rect 55966 9329 56000 9363
rect 56170 9329 56204 9363
rect 56374 9329 56408 9363
rect 56578 9329 56612 9363
rect 56782 9329 56816 9363
rect 56986 9329 57020 9363
rect 57190 9329 57224 9363
rect 57394 9329 57428 9363
rect 57598 9329 57632 9363
rect 57802 9329 57836 9363
rect 58006 9329 58040 9363
rect 58210 9329 58244 9363
rect 58414 9329 58448 9363
rect 58618 9329 58652 9363
rect 58822 9329 58856 9363
rect 59026 9329 59060 9363
rect 59230 9329 59264 9363
rect 59434 9329 59468 9363
rect 59638 9329 59672 9363
rect 59842 9329 59876 9363
rect 60046 9329 60080 9363
rect 60250 9329 60284 9363
rect 8230 7734 8264 7768
rect 8434 7734 8468 7768
rect 8638 7734 8672 7768
rect 8842 7734 8876 7768
rect 9046 7734 9080 7768
rect 9250 7734 9284 7768
rect 9454 7734 9488 7768
rect 9658 7734 9692 7768
rect 9862 7734 9896 7768
rect 10066 7734 10100 7768
rect 10270 7734 10304 7768
rect 10474 7734 10508 7768
rect 10678 7734 10712 7768
rect 10882 7734 10916 7768
rect 11086 7734 11120 7768
rect 11290 7734 11324 7768
rect 11494 7734 11528 7768
rect 11698 7734 11732 7768
rect 11902 7734 11936 7768
rect 12106 7734 12140 7768
rect 12310 7734 12344 7768
rect 12514 7734 12548 7768
rect 12718 7734 12752 7768
rect 12922 7734 12956 7768
rect 13126 7734 13160 7768
rect 13330 7734 13364 7768
rect 13534 7734 13568 7768
rect 13738 7734 13772 7768
rect 13942 7734 13976 7768
rect 14146 7734 14180 7768
rect 14350 7734 14384 7768
rect 14554 7734 14588 7768
rect 14758 7734 14792 7768
rect 14962 7734 14996 7768
rect 15166 7734 15200 7768
rect 15370 7734 15404 7768
rect 15574 7734 15608 7768
rect 15778 7734 15812 7768
rect 15982 7734 16016 7768
rect 16186 7734 16220 7768
rect 16390 7734 16424 7768
rect 16594 7734 16628 7768
rect 16798 7734 16832 7768
rect 17002 7734 17036 7768
rect 17206 7734 17240 7768
rect 17410 7734 17444 7768
rect 17614 7734 17648 7768
rect 17818 7734 17852 7768
rect 18022 7734 18056 7768
rect 18226 7734 18260 7768
rect 18430 7734 18464 7768
rect 18634 7734 18668 7768
rect 18838 7734 18872 7768
rect 19042 7734 19076 7768
rect 19246 7734 19280 7768
rect 19450 7734 19484 7768
rect 19654 7734 19688 7768
rect 19858 7734 19892 7768
rect 20062 7734 20096 7768
rect 20266 7734 20300 7768
rect 20470 7734 20504 7768
rect 20674 7734 20708 7768
rect 20878 7734 20912 7768
rect 21082 7734 21116 7768
rect 21286 7734 21320 7768
rect 21490 7734 21524 7768
rect 21694 7734 21728 7768
rect 21898 7734 21932 7768
rect 22102 7734 22136 7768
rect 22306 7734 22340 7768
rect 22510 7734 22544 7768
rect 22714 7734 22748 7768
rect 22918 7734 22952 7768
rect 23122 7734 23156 7768
rect 23326 7734 23360 7768
rect 23530 7734 23564 7768
rect 23734 7734 23768 7768
rect 23938 7734 23972 7768
rect 24142 7734 24176 7768
rect 24346 7734 24380 7768
rect 24550 7734 24584 7768
rect 24754 7734 24788 7768
rect 24958 7734 24992 7768
rect 25162 7734 25196 7768
rect 25366 7734 25400 7768
rect 25570 7734 25604 7768
rect 25774 7734 25808 7768
rect 25978 7734 26012 7768
rect 26182 7734 26216 7768
rect 26386 7734 26420 7768
rect 26590 7734 26624 7768
rect 26794 7734 26828 7768
rect 26998 7734 27032 7768
rect 27202 7734 27236 7768
rect 27406 7734 27440 7768
rect 27610 7734 27644 7768
rect 27814 7734 27848 7768
rect 28018 7734 28052 7768
rect 28222 7734 28256 7768
rect 28426 7734 28460 7768
rect 28630 7734 28664 7768
rect 28834 7734 28868 7768
rect 29038 7734 29072 7768
rect 29242 7734 29276 7768
rect 29446 7734 29480 7768
rect 29650 7734 29684 7768
rect 29854 7734 29888 7768
rect 30058 7734 30092 7768
rect 30262 7734 30296 7768
rect 30466 7734 30500 7768
rect 30670 7734 30704 7768
rect 30874 7734 30908 7768
rect 31078 7734 31112 7768
rect 31282 7734 31316 7768
rect 31486 7734 31520 7768
rect 31690 7734 31724 7768
rect 31894 7734 31928 7768
rect 32098 7734 32132 7768
rect 32302 7734 32336 7768
rect 32506 7734 32540 7768
rect 32710 7734 32744 7768
rect 32914 7734 32948 7768
rect 33118 7734 33152 7768
rect 33322 7734 33356 7768
rect 33526 7734 33560 7768
rect 33730 7734 33764 7768
rect 33934 7734 33968 7768
rect 34138 7734 34172 7768
rect 34342 7734 34376 7768
rect 34546 7734 34580 7768
rect 34750 7734 34784 7768
rect 34954 7734 34988 7768
rect 35158 7734 35192 7768
rect 35362 7734 35396 7768
rect 35566 7734 35600 7768
rect 35770 7734 35804 7768
rect 35974 7734 36008 7768
rect 36178 7734 36212 7768
rect 36382 7734 36416 7768
rect 36586 7734 36620 7768
rect 36790 7734 36824 7768
rect 36994 7734 37028 7768
rect 37198 7734 37232 7768
rect 37402 7734 37436 7768
rect 37606 7734 37640 7768
rect 37810 7734 37844 7768
rect 38014 7734 38048 7768
rect 38218 7734 38252 7768
rect 38422 7734 38456 7768
rect 38626 7734 38660 7768
rect 38830 7734 38864 7768
rect 39034 7734 39068 7768
rect 39238 7734 39272 7768
rect 39442 7734 39476 7768
rect 39646 7734 39680 7768
rect 39850 7734 39884 7768
rect 40054 7734 40088 7768
rect 40258 7734 40292 7768
rect 40462 7734 40496 7768
rect 40666 7734 40700 7768
rect 40870 7734 40904 7768
rect 41074 7734 41108 7768
rect 41278 7734 41312 7768
rect 41482 7734 41516 7768
rect 41686 7734 41720 7768
rect 41890 7734 41924 7768
rect 42094 7734 42128 7768
rect 42298 7734 42332 7768
rect 42502 7734 42536 7768
rect 42706 7734 42740 7768
rect 42910 7734 42944 7768
rect 43114 7734 43148 7768
rect 43318 7734 43352 7768
rect 43522 7734 43556 7768
rect 43726 7734 43760 7768
rect 43930 7734 43964 7768
rect 44134 7734 44168 7768
rect 44338 7734 44372 7768
rect 44542 7734 44576 7768
rect 44746 7734 44780 7768
rect 44950 7734 44984 7768
rect 45154 7734 45188 7768
rect 45358 7734 45392 7768
rect 45562 7734 45596 7768
rect 45766 7734 45800 7768
rect 45970 7734 46004 7768
rect 46174 7734 46208 7768
rect 46378 7734 46412 7768
rect 46582 7734 46616 7768
rect 46786 7734 46820 7768
rect 46990 7734 47024 7768
rect 47194 7734 47228 7768
rect 47398 7734 47432 7768
rect 47602 7734 47636 7768
rect 47806 7734 47840 7768
rect 48010 7734 48044 7768
rect 48214 7734 48248 7768
rect 48418 7734 48452 7768
rect 48622 7734 48656 7768
rect 48826 7734 48860 7768
rect 49030 7734 49064 7768
rect 49234 7734 49268 7768
rect 49438 7734 49472 7768
rect 49642 7734 49676 7768
rect 49846 7734 49880 7768
rect 50050 7734 50084 7768
rect 50254 7734 50288 7768
rect 50458 7734 50492 7768
rect 50662 7734 50696 7768
rect 50866 7734 50900 7768
rect 51070 7734 51104 7768
rect 51274 7734 51308 7768
rect 51478 7734 51512 7768
rect 51682 7734 51716 7768
rect 51886 7734 51920 7768
rect 52090 7734 52124 7768
rect 52294 7734 52328 7768
rect 52498 7734 52532 7768
rect 52702 7734 52736 7768
rect 52906 7734 52940 7768
rect 53110 7734 53144 7768
rect 53314 7734 53348 7768
rect 53518 7734 53552 7768
rect 53722 7734 53756 7768
rect 53926 7734 53960 7768
rect 54130 7734 54164 7768
rect 54334 7734 54368 7768
rect 54538 7734 54572 7768
rect 54742 7734 54776 7768
rect 54946 7734 54980 7768
rect 55150 7734 55184 7768
rect 55354 7734 55388 7768
rect 55558 7734 55592 7768
rect 55762 7734 55796 7768
rect 55966 7734 56000 7768
rect 56170 7734 56204 7768
rect 56374 7734 56408 7768
rect 56578 7734 56612 7768
rect 56782 7734 56816 7768
rect 56986 7734 57020 7768
rect 57190 7734 57224 7768
rect 57394 7734 57428 7768
rect 57598 7734 57632 7768
rect 57802 7734 57836 7768
rect 58006 7734 58040 7768
rect 58210 7734 58244 7768
rect 58414 7734 58448 7768
rect 58618 7734 58652 7768
rect 58822 7734 58856 7768
rect 59026 7734 59060 7768
rect 59230 7734 59264 7768
rect 59434 7734 59468 7768
rect 59638 7734 59672 7768
rect 59842 7734 59876 7768
rect 60046 7734 60080 7768
rect 60250 7734 60284 7768
rect 337 7059 371 7093
rect 745 7059 779 7093
rect 1153 7059 1187 7093
rect 7959 6379 7993 6413
rect 7959 6175 7993 6209
rect 7959 5971 7993 6005
rect 7959 5767 7993 5801
rect 2993 5588 3027 5622
rect 7959 5563 7993 5597
rect 7959 5359 7993 5393
rect 7959 5155 7993 5189
rect 7959 4951 7993 4985
rect -1386 2923 -1352 2957
rect 51 2961 85 2995
rect 458 1916 492 1950
rect 14692 1705 14726 1739
rect 15000 1705 15034 1739
rect 15308 1705 15342 1739
rect 15616 1705 15650 1739
rect 15924 1705 15958 1739
rect 16232 1705 16266 1739
rect 16540 1705 16574 1739
rect 16848 1705 16882 1739
rect 17156 1705 17190 1739
rect 17464 1705 17498 1739
rect 17772 1705 17806 1739
rect 18080 1705 18114 1739
rect 18388 1705 18422 1739
rect 18696 1705 18730 1739
rect 19004 1705 19038 1739
rect 19312 1705 19346 1739
rect 19620 1705 19654 1739
rect 19928 1705 19962 1739
rect 20236 1705 20270 1739
rect 20544 1705 20578 1739
rect 20852 1705 20886 1739
rect 21160 1705 21194 1739
rect 21468 1705 21502 1739
rect 21776 1705 21810 1739
rect 22084 1705 22118 1739
rect 22392 1705 22426 1739
rect 22700 1705 22734 1739
rect 23008 1705 23042 1739
rect 23316 1705 23350 1739
rect 23624 1705 23658 1739
rect 23932 1705 23966 1739
rect 24240 1705 24274 1739
rect 4835 1590 4869 1624
rect 5243 1590 5277 1624
rect 5651 1590 5685 1624
rect 14692 0 14726 34
rect 15000 0 15034 34
rect 15308 0 15342 34
rect 15616 0 15650 34
rect 15924 0 15958 34
rect 16232 0 16266 34
rect 16540 0 16574 34
rect 16848 0 16882 34
rect 17156 0 17190 34
rect 17464 0 17498 34
rect 17772 0 17806 34
rect 18080 0 18114 34
rect 18388 0 18422 34
rect 18696 0 18730 34
rect 19004 0 19038 34
rect 19312 0 19346 34
rect 19620 0 19654 34
rect 19928 0 19962 34
rect 20236 0 20270 34
rect 20544 0 20578 34
rect 20852 0 20886 34
rect 21160 0 21194 34
rect 21468 0 21502 34
rect 21776 0 21810 34
rect 22084 0 22118 34
rect 22392 0 22426 34
rect 22700 0 22734 34
rect 23008 0 23042 34
rect 23316 0 23350 34
rect 23624 0 23658 34
rect 23932 0 23966 34
rect 24240 0 24274 34
<< metal1 >>
rect 8201 12170 8207 12222
rect 8259 12170 8265 12222
rect 60249 12170 60255 12222
rect 60307 12170 60313 12222
rect 2731 11959 2737 12011
rect 2789 11959 2795 12011
rect 3979 11959 3985 12011
rect 4037 11959 4043 12011
rect 5577 11959 5583 12011
rect 5635 11959 5641 12011
rect 7225 11959 7231 12011
rect 7283 11959 7289 12011
rect 7947 11882 8005 11888
rect 7947 11848 7959 11882
rect 7993 11879 8005 11882
rect 8106 11879 8112 11891
rect 7993 11851 8112 11879
rect 7993 11848 8005 11851
rect 7947 11842 8005 11848
rect 8106 11839 8112 11851
rect 8164 11839 8170 11891
rect 7947 11678 8005 11684
rect 7947 11644 7959 11678
rect 7993 11675 8005 11678
rect 8106 11675 8112 11687
rect 7993 11647 8112 11675
rect 7993 11644 8005 11647
rect 7947 11638 8005 11644
rect 8106 11635 8112 11647
rect 8164 11635 8170 11687
rect 7947 11474 8005 11480
rect 7947 11440 7959 11474
rect 7993 11471 8005 11474
rect 8106 11471 8112 11483
rect 7993 11443 8112 11471
rect 7993 11440 8005 11443
rect 7947 11434 8005 11440
rect 8106 11431 8112 11443
rect 8164 11431 8170 11483
rect 7947 11270 8005 11276
rect 7947 11236 7959 11270
rect 7993 11267 8005 11270
rect 8106 11267 8112 11279
rect 7993 11239 8112 11267
rect 7993 11236 8005 11239
rect 7947 11230 8005 11236
rect 8106 11227 8112 11239
rect 8164 11227 8170 11279
rect 7947 11066 8005 11072
rect 7947 11032 7959 11066
rect 7993 11063 8005 11066
rect 8106 11063 8112 11075
rect 7993 11035 8112 11063
rect 7993 11032 8005 11035
rect 7947 11026 8005 11032
rect 8106 11023 8112 11035
rect 8164 11023 8170 11075
rect 7947 10862 8005 10868
rect 7947 10828 7959 10862
rect 7993 10859 8005 10862
rect 8106 10859 8112 10871
rect 7993 10831 8112 10859
rect 7993 10828 8005 10831
rect 7947 10822 8005 10828
rect 8106 10819 8112 10831
rect 8164 10819 8170 10871
rect 7947 10658 8005 10664
rect 7947 10624 7959 10658
rect 7993 10655 8005 10658
rect 8106 10655 8112 10667
rect 7993 10627 8112 10655
rect 7993 10624 8005 10627
rect 7947 10618 8005 10624
rect 8106 10615 8112 10627
rect 8164 10615 8170 10667
rect 7947 10454 8005 10460
rect 7947 10420 7959 10454
rect 7993 10451 8005 10454
rect 8106 10451 8112 10463
rect 7993 10423 8112 10451
rect 7993 10420 8005 10423
rect 7947 10414 8005 10420
rect 8106 10411 8112 10423
rect 8164 10411 8170 10463
rect 2731 10243 2737 10295
rect 2789 10243 2795 10295
rect 3979 10243 3985 10295
rect 4037 10243 4043 10295
rect 5577 10243 5583 10295
rect 5635 10243 5641 10295
rect 7225 10243 7231 10295
rect 7283 10243 7289 10295
rect 109 9820 115 9872
rect 167 9820 173 9872
rect 8148 9806 8154 9818
rect 6375 9778 8154 9806
rect 1333 9395 1339 9447
rect 1391 9395 1397 9447
rect 1403 9187 1409 9199
rect 1351 9159 1409 9187
rect 1403 9147 1409 9159
rect 1461 9147 1467 9199
rect 109 8868 115 8920
rect 167 8868 173 8920
rect 1333 8443 1339 8495
rect 1391 8443 1397 8495
rect 109 7831 115 7883
rect 167 7831 173 7883
rect 1333 7209 1339 7261
rect 1391 7209 1397 7261
rect 322 7050 328 7102
rect 380 7050 386 7102
rect 730 7050 736 7102
rect 788 7050 794 7102
rect 1138 7050 1144 7102
rect 1196 7050 1202 7102
rect 6375 6787 6403 9778
rect 8148 9766 8154 9778
rect 8206 9766 8212 9818
rect 8233 9375 8261 9424
rect 8437 9375 8465 9424
rect 8641 9375 8669 9424
rect 8845 9375 8873 9424
rect 9049 9375 9077 9424
rect 9253 9375 9281 9424
rect 9457 9375 9485 9424
rect 9661 9375 9689 9424
rect 9865 9375 9893 9424
rect 10069 9375 10097 9424
rect 10273 9375 10301 9424
rect 10477 9375 10505 9424
rect 10681 9375 10709 9424
rect 10885 9375 10913 9424
rect 11089 9375 11117 9424
rect 11293 9375 11321 9424
rect 11497 9375 11525 9424
rect 11701 9375 11729 9424
rect 11905 9375 11933 9424
rect 12109 9375 12137 9424
rect 12313 9375 12341 9424
rect 12517 9375 12545 9424
rect 12721 9375 12749 9424
rect 12925 9375 12953 9424
rect 13129 9375 13157 9424
rect 13333 9375 13361 9424
rect 13537 9375 13565 9424
rect 13741 9375 13769 9424
rect 13945 9375 13973 9424
rect 14149 9375 14177 9424
rect 14353 9375 14381 9424
rect 14557 9375 14585 9424
rect 14761 9375 14789 9424
rect 14965 9375 14993 9424
rect 15169 9375 15197 9424
rect 15373 9375 15401 9424
rect 15577 9375 15605 9424
rect 15781 9375 15809 9424
rect 15985 9375 16013 9424
rect 16189 9375 16217 9424
rect 16393 9375 16421 9424
rect 16597 9375 16625 9424
rect 16801 9375 16829 9424
rect 17005 9375 17033 9424
rect 17209 9375 17237 9424
rect 17413 9375 17441 9424
rect 17617 9375 17645 9424
rect 17821 9375 17849 9424
rect 18025 9375 18053 9424
rect 18229 9375 18257 9424
rect 18433 9375 18461 9424
rect 18637 9375 18665 9424
rect 18841 9375 18869 9424
rect 19045 9375 19073 9424
rect 19249 9375 19277 9424
rect 19453 9375 19481 9424
rect 19657 9375 19685 9424
rect 19861 9375 19889 9424
rect 20065 9375 20093 9424
rect 20269 9375 20297 9424
rect 20473 9375 20501 9424
rect 20677 9375 20705 9424
rect 20881 9375 20909 9424
rect 21085 9375 21113 9424
rect 21289 9375 21317 9424
rect 21493 9375 21521 9424
rect 21697 9375 21725 9424
rect 21901 9375 21929 9424
rect 22105 9375 22133 9424
rect 22309 9375 22337 9424
rect 22513 9375 22541 9424
rect 22717 9375 22745 9424
rect 22921 9375 22949 9424
rect 23125 9375 23153 9424
rect 23329 9375 23357 9424
rect 23533 9375 23561 9424
rect 23737 9375 23765 9424
rect 23941 9375 23969 9424
rect 24145 9375 24173 9424
rect 24349 9375 24377 9424
rect 24553 9375 24581 9424
rect 24757 9375 24785 9424
rect 24961 9375 24989 9424
rect 25165 9375 25193 9424
rect 25369 9375 25397 9424
rect 25573 9375 25601 9424
rect 25777 9375 25805 9424
rect 25981 9375 26009 9424
rect 26185 9375 26213 9424
rect 26389 9375 26417 9424
rect 26593 9375 26621 9424
rect 26797 9375 26825 9424
rect 27001 9375 27029 9424
rect 27205 9375 27233 9424
rect 27409 9375 27437 9424
rect 27613 9375 27641 9424
rect 27817 9375 27845 9424
rect 28021 9375 28049 9424
rect 28225 9375 28253 9424
rect 28429 9375 28457 9424
rect 28633 9375 28661 9424
rect 28837 9375 28865 9424
rect 29041 9375 29069 9424
rect 29245 9375 29273 9424
rect 29449 9375 29477 9424
rect 29653 9375 29681 9424
rect 29857 9375 29885 9424
rect 30061 9375 30089 9424
rect 30265 9375 30293 9424
rect 30469 9375 30497 9424
rect 30673 9375 30701 9424
rect 30877 9375 30905 9424
rect 31081 9375 31109 9424
rect 31285 9375 31313 9424
rect 31489 9375 31517 9424
rect 31693 9375 31721 9424
rect 31897 9375 31925 9424
rect 32101 9375 32129 9424
rect 32305 9375 32333 9424
rect 32509 9375 32537 9424
rect 32713 9375 32741 9424
rect 32917 9375 32945 9424
rect 33121 9375 33149 9424
rect 33325 9375 33353 9424
rect 33529 9375 33557 9424
rect 33733 9375 33761 9424
rect 33937 9375 33965 9424
rect 34141 9375 34169 9424
rect 34345 9375 34373 9424
rect 34549 9375 34577 9424
rect 34753 9375 34781 9424
rect 34957 9375 34985 9424
rect 35161 9375 35189 9424
rect 35365 9375 35393 9424
rect 35569 9375 35597 9424
rect 35773 9375 35801 9424
rect 35977 9375 36005 9424
rect 36181 9375 36209 9424
rect 36385 9375 36413 9424
rect 36589 9375 36617 9424
rect 36793 9375 36821 9424
rect 36997 9375 37025 9424
rect 37201 9375 37229 9424
rect 37405 9375 37433 9424
rect 37609 9375 37637 9424
rect 37813 9375 37841 9424
rect 38017 9375 38045 9424
rect 38221 9375 38249 9424
rect 38425 9375 38453 9424
rect 38629 9375 38657 9424
rect 38833 9375 38861 9424
rect 39037 9375 39065 9424
rect 39241 9375 39269 9424
rect 39445 9375 39473 9424
rect 39649 9375 39677 9424
rect 39853 9375 39881 9424
rect 40057 9375 40085 9424
rect 40261 9375 40289 9424
rect 40465 9375 40493 9424
rect 40669 9375 40697 9424
rect 40873 9375 40901 9424
rect 41077 9375 41105 9424
rect 41281 9375 41309 9424
rect 41485 9375 41513 9424
rect 41689 9375 41717 9424
rect 41893 9375 41921 9424
rect 42097 9375 42125 9424
rect 42301 9375 42329 9424
rect 42505 9375 42533 9424
rect 42709 9375 42737 9424
rect 42913 9375 42941 9424
rect 43117 9375 43145 9424
rect 43321 9375 43349 9424
rect 43525 9375 43553 9424
rect 43729 9375 43757 9424
rect 43933 9375 43961 9424
rect 44137 9375 44165 9424
rect 44341 9375 44369 9424
rect 44545 9375 44573 9424
rect 44749 9375 44777 9424
rect 44953 9375 44981 9424
rect 45157 9375 45185 9424
rect 45361 9375 45389 9424
rect 45565 9375 45593 9424
rect 45769 9375 45797 9424
rect 45973 9375 46001 9424
rect 46177 9375 46205 9424
rect 46381 9375 46409 9424
rect 46585 9375 46613 9424
rect 46789 9375 46817 9424
rect 46993 9375 47021 9424
rect 47197 9375 47225 9424
rect 47401 9375 47429 9424
rect 47605 9375 47633 9424
rect 47809 9375 47837 9424
rect 48013 9375 48041 9424
rect 48217 9375 48245 9424
rect 48421 9375 48449 9424
rect 48625 9375 48653 9424
rect 48829 9375 48857 9424
rect 49033 9375 49061 9424
rect 49237 9375 49265 9424
rect 49441 9375 49469 9424
rect 49645 9375 49673 9424
rect 49849 9375 49877 9424
rect 50053 9375 50081 9424
rect 50257 9375 50285 9424
rect 50461 9375 50489 9424
rect 50665 9375 50693 9424
rect 50869 9375 50897 9424
rect 51073 9375 51101 9424
rect 51277 9375 51305 9424
rect 51481 9375 51509 9424
rect 51685 9375 51713 9424
rect 51889 9375 51917 9424
rect 52093 9375 52121 9424
rect 52297 9375 52325 9424
rect 52501 9375 52529 9424
rect 52705 9375 52733 9424
rect 52909 9375 52937 9424
rect 53113 9375 53141 9424
rect 53317 9375 53345 9424
rect 53521 9375 53549 9424
rect 53725 9375 53753 9424
rect 53929 9375 53957 9424
rect 54133 9375 54161 9424
rect 54337 9375 54365 9424
rect 54541 9375 54569 9424
rect 54745 9375 54773 9424
rect 54949 9375 54977 9424
rect 55153 9375 55181 9424
rect 55357 9375 55385 9424
rect 55561 9375 55589 9424
rect 55765 9375 55793 9424
rect 55969 9375 55997 9424
rect 56173 9375 56201 9424
rect 56377 9375 56405 9424
rect 56581 9375 56609 9424
rect 56785 9375 56813 9424
rect 56989 9375 57017 9424
rect 57193 9375 57221 9424
rect 57397 9375 57425 9424
rect 57601 9375 57629 9424
rect 57805 9375 57833 9424
rect 58009 9375 58037 9424
rect 58213 9375 58241 9424
rect 58417 9375 58445 9424
rect 58621 9375 58649 9424
rect 58825 9375 58853 9424
rect 59029 9375 59057 9424
rect 59233 9375 59261 9424
rect 59437 9375 59465 9424
rect 59641 9375 59669 9424
rect 59845 9375 59873 9424
rect 60049 9375 60077 9424
rect 60253 9375 60281 9424
rect 8224 9363 8270 9375
rect 8224 9329 8230 9363
rect 8264 9329 8270 9363
rect 8224 9317 8270 9329
rect 8428 9363 8474 9375
rect 8428 9329 8434 9363
rect 8468 9329 8474 9363
rect 8428 9317 8474 9329
rect 8632 9363 8678 9375
rect 8632 9329 8638 9363
rect 8672 9329 8678 9363
rect 8632 9317 8678 9329
rect 8836 9363 8882 9375
rect 8836 9329 8842 9363
rect 8876 9329 8882 9363
rect 8836 9317 8882 9329
rect 9040 9363 9086 9375
rect 9040 9329 9046 9363
rect 9080 9329 9086 9363
rect 9040 9317 9086 9329
rect 9244 9363 9290 9375
rect 9244 9329 9250 9363
rect 9284 9329 9290 9363
rect 9244 9317 9290 9329
rect 9448 9363 9494 9375
rect 9448 9329 9454 9363
rect 9488 9329 9494 9363
rect 9448 9317 9494 9329
rect 9652 9363 9698 9375
rect 9652 9329 9658 9363
rect 9692 9329 9698 9363
rect 9652 9317 9698 9329
rect 9856 9363 9902 9375
rect 9856 9329 9862 9363
rect 9896 9329 9902 9363
rect 9856 9317 9902 9329
rect 10060 9363 10106 9375
rect 10060 9329 10066 9363
rect 10100 9329 10106 9363
rect 10060 9317 10106 9329
rect 10264 9363 10310 9375
rect 10264 9329 10270 9363
rect 10304 9329 10310 9363
rect 10264 9317 10310 9329
rect 10468 9363 10514 9375
rect 10468 9329 10474 9363
rect 10508 9329 10514 9363
rect 10468 9317 10514 9329
rect 10672 9363 10718 9375
rect 10672 9329 10678 9363
rect 10712 9329 10718 9363
rect 10672 9317 10718 9329
rect 10876 9363 10922 9375
rect 10876 9329 10882 9363
rect 10916 9329 10922 9363
rect 10876 9317 10922 9329
rect 11080 9363 11126 9375
rect 11080 9329 11086 9363
rect 11120 9329 11126 9363
rect 11080 9317 11126 9329
rect 11284 9363 11330 9375
rect 11284 9329 11290 9363
rect 11324 9329 11330 9363
rect 11284 9317 11330 9329
rect 11488 9363 11534 9375
rect 11488 9329 11494 9363
rect 11528 9329 11534 9363
rect 11488 9317 11534 9329
rect 11692 9363 11738 9375
rect 11692 9329 11698 9363
rect 11732 9329 11738 9363
rect 11692 9317 11738 9329
rect 11896 9363 11942 9375
rect 11896 9329 11902 9363
rect 11936 9329 11942 9363
rect 11896 9317 11942 9329
rect 12100 9363 12146 9375
rect 12100 9329 12106 9363
rect 12140 9329 12146 9363
rect 12100 9317 12146 9329
rect 12304 9363 12350 9375
rect 12304 9329 12310 9363
rect 12344 9329 12350 9363
rect 12304 9317 12350 9329
rect 12508 9363 12554 9375
rect 12508 9329 12514 9363
rect 12548 9329 12554 9363
rect 12508 9317 12554 9329
rect 12712 9363 12758 9375
rect 12712 9329 12718 9363
rect 12752 9329 12758 9363
rect 12712 9317 12758 9329
rect 12916 9363 12962 9375
rect 12916 9329 12922 9363
rect 12956 9329 12962 9363
rect 12916 9317 12962 9329
rect 13120 9363 13166 9375
rect 13120 9329 13126 9363
rect 13160 9329 13166 9363
rect 13120 9317 13166 9329
rect 13324 9363 13370 9375
rect 13324 9329 13330 9363
rect 13364 9329 13370 9363
rect 13324 9317 13370 9329
rect 13528 9363 13574 9375
rect 13528 9329 13534 9363
rect 13568 9329 13574 9363
rect 13528 9317 13574 9329
rect 13732 9363 13778 9375
rect 13732 9329 13738 9363
rect 13772 9329 13778 9363
rect 13732 9317 13778 9329
rect 13936 9363 13982 9375
rect 13936 9329 13942 9363
rect 13976 9329 13982 9363
rect 13936 9317 13982 9329
rect 14140 9363 14186 9375
rect 14140 9329 14146 9363
rect 14180 9329 14186 9363
rect 14140 9317 14186 9329
rect 14344 9363 14390 9375
rect 14344 9329 14350 9363
rect 14384 9329 14390 9363
rect 14344 9317 14390 9329
rect 14548 9363 14594 9375
rect 14548 9329 14554 9363
rect 14588 9329 14594 9363
rect 14548 9317 14594 9329
rect 14752 9363 14798 9375
rect 14752 9329 14758 9363
rect 14792 9329 14798 9363
rect 14752 9317 14798 9329
rect 14956 9363 15002 9375
rect 14956 9329 14962 9363
rect 14996 9329 15002 9363
rect 14956 9317 15002 9329
rect 15160 9363 15206 9375
rect 15160 9329 15166 9363
rect 15200 9329 15206 9363
rect 15160 9317 15206 9329
rect 15364 9363 15410 9375
rect 15364 9329 15370 9363
rect 15404 9329 15410 9363
rect 15364 9317 15410 9329
rect 15568 9363 15614 9375
rect 15568 9329 15574 9363
rect 15608 9329 15614 9363
rect 15568 9317 15614 9329
rect 15772 9363 15818 9375
rect 15772 9329 15778 9363
rect 15812 9329 15818 9363
rect 15772 9317 15818 9329
rect 15976 9363 16022 9375
rect 15976 9329 15982 9363
rect 16016 9329 16022 9363
rect 15976 9317 16022 9329
rect 16180 9363 16226 9375
rect 16180 9329 16186 9363
rect 16220 9329 16226 9363
rect 16180 9317 16226 9329
rect 16384 9363 16430 9375
rect 16384 9329 16390 9363
rect 16424 9329 16430 9363
rect 16384 9317 16430 9329
rect 16588 9363 16634 9375
rect 16588 9329 16594 9363
rect 16628 9329 16634 9363
rect 16588 9317 16634 9329
rect 16792 9363 16838 9375
rect 16792 9329 16798 9363
rect 16832 9329 16838 9363
rect 16792 9317 16838 9329
rect 16996 9363 17042 9375
rect 16996 9329 17002 9363
rect 17036 9329 17042 9363
rect 16996 9317 17042 9329
rect 17200 9363 17246 9375
rect 17200 9329 17206 9363
rect 17240 9329 17246 9363
rect 17200 9317 17246 9329
rect 17404 9363 17450 9375
rect 17404 9329 17410 9363
rect 17444 9329 17450 9363
rect 17404 9317 17450 9329
rect 17608 9363 17654 9375
rect 17608 9329 17614 9363
rect 17648 9329 17654 9363
rect 17608 9317 17654 9329
rect 17812 9363 17858 9375
rect 17812 9329 17818 9363
rect 17852 9329 17858 9363
rect 17812 9317 17858 9329
rect 18016 9363 18062 9375
rect 18016 9329 18022 9363
rect 18056 9329 18062 9363
rect 18016 9317 18062 9329
rect 18220 9363 18266 9375
rect 18220 9329 18226 9363
rect 18260 9329 18266 9363
rect 18220 9317 18266 9329
rect 18424 9363 18470 9375
rect 18424 9329 18430 9363
rect 18464 9329 18470 9363
rect 18424 9317 18470 9329
rect 18628 9363 18674 9375
rect 18628 9329 18634 9363
rect 18668 9329 18674 9363
rect 18628 9317 18674 9329
rect 18832 9363 18878 9375
rect 18832 9329 18838 9363
rect 18872 9329 18878 9363
rect 18832 9317 18878 9329
rect 19036 9363 19082 9375
rect 19036 9329 19042 9363
rect 19076 9329 19082 9363
rect 19036 9317 19082 9329
rect 19240 9363 19286 9375
rect 19240 9329 19246 9363
rect 19280 9329 19286 9363
rect 19240 9317 19286 9329
rect 19444 9363 19490 9375
rect 19444 9329 19450 9363
rect 19484 9329 19490 9363
rect 19444 9317 19490 9329
rect 19648 9363 19694 9375
rect 19648 9329 19654 9363
rect 19688 9329 19694 9363
rect 19648 9317 19694 9329
rect 19852 9363 19898 9375
rect 19852 9329 19858 9363
rect 19892 9329 19898 9363
rect 19852 9317 19898 9329
rect 20056 9363 20102 9375
rect 20056 9329 20062 9363
rect 20096 9329 20102 9363
rect 20056 9317 20102 9329
rect 20260 9363 20306 9375
rect 20260 9329 20266 9363
rect 20300 9329 20306 9363
rect 20260 9317 20306 9329
rect 20464 9363 20510 9375
rect 20464 9329 20470 9363
rect 20504 9329 20510 9363
rect 20464 9317 20510 9329
rect 20668 9363 20714 9375
rect 20668 9329 20674 9363
rect 20708 9329 20714 9363
rect 20668 9317 20714 9329
rect 20872 9363 20918 9375
rect 20872 9329 20878 9363
rect 20912 9329 20918 9363
rect 20872 9317 20918 9329
rect 21076 9363 21122 9375
rect 21076 9329 21082 9363
rect 21116 9329 21122 9363
rect 21076 9317 21122 9329
rect 21280 9363 21326 9375
rect 21280 9329 21286 9363
rect 21320 9329 21326 9363
rect 21280 9317 21326 9329
rect 21484 9363 21530 9375
rect 21484 9329 21490 9363
rect 21524 9329 21530 9363
rect 21484 9317 21530 9329
rect 21688 9363 21734 9375
rect 21688 9329 21694 9363
rect 21728 9329 21734 9363
rect 21688 9317 21734 9329
rect 21892 9363 21938 9375
rect 21892 9329 21898 9363
rect 21932 9329 21938 9363
rect 21892 9317 21938 9329
rect 22096 9363 22142 9375
rect 22096 9329 22102 9363
rect 22136 9329 22142 9363
rect 22096 9317 22142 9329
rect 22300 9363 22346 9375
rect 22300 9329 22306 9363
rect 22340 9329 22346 9363
rect 22300 9317 22346 9329
rect 22504 9363 22550 9375
rect 22504 9329 22510 9363
rect 22544 9329 22550 9363
rect 22504 9317 22550 9329
rect 22708 9363 22754 9375
rect 22708 9329 22714 9363
rect 22748 9329 22754 9363
rect 22708 9317 22754 9329
rect 22912 9363 22958 9375
rect 22912 9329 22918 9363
rect 22952 9329 22958 9363
rect 22912 9317 22958 9329
rect 23116 9363 23162 9375
rect 23116 9329 23122 9363
rect 23156 9329 23162 9363
rect 23116 9317 23162 9329
rect 23320 9363 23366 9375
rect 23320 9329 23326 9363
rect 23360 9329 23366 9363
rect 23320 9317 23366 9329
rect 23524 9363 23570 9375
rect 23524 9329 23530 9363
rect 23564 9329 23570 9363
rect 23524 9317 23570 9329
rect 23728 9363 23774 9375
rect 23728 9329 23734 9363
rect 23768 9329 23774 9363
rect 23728 9317 23774 9329
rect 23932 9363 23978 9375
rect 23932 9329 23938 9363
rect 23972 9329 23978 9363
rect 23932 9317 23978 9329
rect 24136 9363 24182 9375
rect 24136 9329 24142 9363
rect 24176 9329 24182 9363
rect 24136 9317 24182 9329
rect 24340 9363 24386 9375
rect 24340 9329 24346 9363
rect 24380 9329 24386 9363
rect 24340 9317 24386 9329
rect 24544 9363 24590 9375
rect 24544 9329 24550 9363
rect 24584 9329 24590 9363
rect 24544 9317 24590 9329
rect 24748 9363 24794 9375
rect 24748 9329 24754 9363
rect 24788 9329 24794 9363
rect 24748 9317 24794 9329
rect 24952 9363 24998 9375
rect 24952 9329 24958 9363
rect 24992 9329 24998 9363
rect 24952 9317 24998 9329
rect 25156 9363 25202 9375
rect 25156 9329 25162 9363
rect 25196 9329 25202 9363
rect 25156 9317 25202 9329
rect 25360 9363 25406 9375
rect 25360 9329 25366 9363
rect 25400 9329 25406 9363
rect 25360 9317 25406 9329
rect 25564 9363 25610 9375
rect 25564 9329 25570 9363
rect 25604 9329 25610 9363
rect 25564 9317 25610 9329
rect 25768 9363 25814 9375
rect 25768 9329 25774 9363
rect 25808 9329 25814 9363
rect 25768 9317 25814 9329
rect 25972 9363 26018 9375
rect 25972 9329 25978 9363
rect 26012 9329 26018 9363
rect 25972 9317 26018 9329
rect 26176 9363 26222 9375
rect 26176 9329 26182 9363
rect 26216 9329 26222 9363
rect 26176 9317 26222 9329
rect 26380 9363 26426 9375
rect 26380 9329 26386 9363
rect 26420 9329 26426 9363
rect 26380 9317 26426 9329
rect 26584 9363 26630 9375
rect 26584 9329 26590 9363
rect 26624 9329 26630 9363
rect 26584 9317 26630 9329
rect 26788 9363 26834 9375
rect 26788 9329 26794 9363
rect 26828 9329 26834 9363
rect 26788 9317 26834 9329
rect 26992 9363 27038 9375
rect 26992 9329 26998 9363
rect 27032 9329 27038 9363
rect 26992 9317 27038 9329
rect 27196 9363 27242 9375
rect 27196 9329 27202 9363
rect 27236 9329 27242 9363
rect 27196 9317 27242 9329
rect 27400 9363 27446 9375
rect 27400 9329 27406 9363
rect 27440 9329 27446 9363
rect 27400 9317 27446 9329
rect 27604 9363 27650 9375
rect 27604 9329 27610 9363
rect 27644 9329 27650 9363
rect 27604 9317 27650 9329
rect 27808 9363 27854 9375
rect 27808 9329 27814 9363
rect 27848 9329 27854 9363
rect 27808 9317 27854 9329
rect 28012 9363 28058 9375
rect 28012 9329 28018 9363
rect 28052 9329 28058 9363
rect 28012 9317 28058 9329
rect 28216 9363 28262 9375
rect 28216 9329 28222 9363
rect 28256 9329 28262 9363
rect 28216 9317 28262 9329
rect 28420 9363 28466 9375
rect 28420 9329 28426 9363
rect 28460 9329 28466 9363
rect 28420 9317 28466 9329
rect 28624 9363 28670 9375
rect 28624 9329 28630 9363
rect 28664 9329 28670 9363
rect 28624 9317 28670 9329
rect 28828 9363 28874 9375
rect 28828 9329 28834 9363
rect 28868 9329 28874 9363
rect 28828 9317 28874 9329
rect 29032 9363 29078 9375
rect 29032 9329 29038 9363
rect 29072 9329 29078 9363
rect 29032 9317 29078 9329
rect 29236 9363 29282 9375
rect 29236 9329 29242 9363
rect 29276 9329 29282 9363
rect 29236 9317 29282 9329
rect 29440 9363 29486 9375
rect 29440 9329 29446 9363
rect 29480 9329 29486 9363
rect 29440 9317 29486 9329
rect 29644 9363 29690 9375
rect 29644 9329 29650 9363
rect 29684 9329 29690 9363
rect 29644 9317 29690 9329
rect 29848 9363 29894 9375
rect 29848 9329 29854 9363
rect 29888 9329 29894 9363
rect 29848 9317 29894 9329
rect 30052 9363 30098 9375
rect 30052 9329 30058 9363
rect 30092 9329 30098 9363
rect 30052 9317 30098 9329
rect 30256 9363 30302 9375
rect 30256 9329 30262 9363
rect 30296 9329 30302 9363
rect 30256 9317 30302 9329
rect 30460 9363 30506 9375
rect 30460 9329 30466 9363
rect 30500 9329 30506 9363
rect 30460 9317 30506 9329
rect 30664 9363 30710 9375
rect 30664 9329 30670 9363
rect 30704 9329 30710 9363
rect 30664 9317 30710 9329
rect 30868 9363 30914 9375
rect 30868 9329 30874 9363
rect 30908 9329 30914 9363
rect 30868 9317 30914 9329
rect 31072 9363 31118 9375
rect 31072 9329 31078 9363
rect 31112 9329 31118 9363
rect 31072 9317 31118 9329
rect 31276 9363 31322 9375
rect 31276 9329 31282 9363
rect 31316 9329 31322 9363
rect 31276 9317 31322 9329
rect 31480 9363 31526 9375
rect 31480 9329 31486 9363
rect 31520 9329 31526 9363
rect 31480 9317 31526 9329
rect 31684 9363 31730 9375
rect 31684 9329 31690 9363
rect 31724 9329 31730 9363
rect 31684 9317 31730 9329
rect 31888 9363 31934 9375
rect 31888 9329 31894 9363
rect 31928 9329 31934 9363
rect 31888 9317 31934 9329
rect 32092 9363 32138 9375
rect 32092 9329 32098 9363
rect 32132 9329 32138 9363
rect 32092 9317 32138 9329
rect 32296 9363 32342 9375
rect 32296 9329 32302 9363
rect 32336 9329 32342 9363
rect 32296 9317 32342 9329
rect 32500 9363 32546 9375
rect 32500 9329 32506 9363
rect 32540 9329 32546 9363
rect 32500 9317 32546 9329
rect 32704 9363 32750 9375
rect 32704 9329 32710 9363
rect 32744 9329 32750 9363
rect 32704 9317 32750 9329
rect 32908 9363 32954 9375
rect 32908 9329 32914 9363
rect 32948 9329 32954 9363
rect 32908 9317 32954 9329
rect 33112 9363 33158 9375
rect 33112 9329 33118 9363
rect 33152 9329 33158 9363
rect 33112 9317 33158 9329
rect 33316 9363 33362 9375
rect 33316 9329 33322 9363
rect 33356 9329 33362 9363
rect 33316 9317 33362 9329
rect 33520 9363 33566 9375
rect 33520 9329 33526 9363
rect 33560 9329 33566 9363
rect 33520 9317 33566 9329
rect 33724 9363 33770 9375
rect 33724 9329 33730 9363
rect 33764 9329 33770 9363
rect 33724 9317 33770 9329
rect 33928 9363 33974 9375
rect 33928 9329 33934 9363
rect 33968 9329 33974 9363
rect 33928 9317 33974 9329
rect 34132 9363 34178 9375
rect 34132 9329 34138 9363
rect 34172 9329 34178 9363
rect 34132 9317 34178 9329
rect 34336 9363 34382 9375
rect 34336 9329 34342 9363
rect 34376 9329 34382 9363
rect 34336 9317 34382 9329
rect 34540 9363 34586 9375
rect 34540 9329 34546 9363
rect 34580 9329 34586 9363
rect 34540 9317 34586 9329
rect 34744 9363 34790 9375
rect 34744 9329 34750 9363
rect 34784 9329 34790 9363
rect 34744 9317 34790 9329
rect 34948 9363 34994 9375
rect 34948 9329 34954 9363
rect 34988 9329 34994 9363
rect 34948 9317 34994 9329
rect 35152 9363 35198 9375
rect 35152 9329 35158 9363
rect 35192 9329 35198 9363
rect 35152 9317 35198 9329
rect 35356 9363 35402 9375
rect 35356 9329 35362 9363
rect 35396 9329 35402 9363
rect 35356 9317 35402 9329
rect 35560 9363 35606 9375
rect 35560 9329 35566 9363
rect 35600 9329 35606 9363
rect 35560 9317 35606 9329
rect 35764 9363 35810 9375
rect 35764 9329 35770 9363
rect 35804 9329 35810 9363
rect 35764 9317 35810 9329
rect 35968 9363 36014 9375
rect 35968 9329 35974 9363
rect 36008 9329 36014 9363
rect 35968 9317 36014 9329
rect 36172 9363 36218 9375
rect 36172 9329 36178 9363
rect 36212 9329 36218 9363
rect 36172 9317 36218 9329
rect 36376 9363 36422 9375
rect 36376 9329 36382 9363
rect 36416 9329 36422 9363
rect 36376 9317 36422 9329
rect 36580 9363 36626 9375
rect 36580 9329 36586 9363
rect 36620 9329 36626 9363
rect 36580 9317 36626 9329
rect 36784 9363 36830 9375
rect 36784 9329 36790 9363
rect 36824 9329 36830 9363
rect 36784 9317 36830 9329
rect 36988 9363 37034 9375
rect 36988 9329 36994 9363
rect 37028 9329 37034 9363
rect 36988 9317 37034 9329
rect 37192 9363 37238 9375
rect 37192 9329 37198 9363
rect 37232 9329 37238 9363
rect 37192 9317 37238 9329
rect 37396 9363 37442 9375
rect 37396 9329 37402 9363
rect 37436 9329 37442 9363
rect 37396 9317 37442 9329
rect 37600 9363 37646 9375
rect 37600 9329 37606 9363
rect 37640 9329 37646 9363
rect 37600 9317 37646 9329
rect 37804 9363 37850 9375
rect 37804 9329 37810 9363
rect 37844 9329 37850 9363
rect 37804 9317 37850 9329
rect 38008 9363 38054 9375
rect 38008 9329 38014 9363
rect 38048 9329 38054 9363
rect 38008 9317 38054 9329
rect 38212 9363 38258 9375
rect 38212 9329 38218 9363
rect 38252 9329 38258 9363
rect 38212 9317 38258 9329
rect 38416 9363 38462 9375
rect 38416 9329 38422 9363
rect 38456 9329 38462 9363
rect 38416 9317 38462 9329
rect 38620 9363 38666 9375
rect 38620 9329 38626 9363
rect 38660 9329 38666 9363
rect 38620 9317 38666 9329
rect 38824 9363 38870 9375
rect 38824 9329 38830 9363
rect 38864 9329 38870 9363
rect 38824 9317 38870 9329
rect 39028 9363 39074 9375
rect 39028 9329 39034 9363
rect 39068 9329 39074 9363
rect 39028 9317 39074 9329
rect 39232 9363 39278 9375
rect 39232 9329 39238 9363
rect 39272 9329 39278 9363
rect 39232 9317 39278 9329
rect 39436 9363 39482 9375
rect 39436 9329 39442 9363
rect 39476 9329 39482 9363
rect 39436 9317 39482 9329
rect 39640 9363 39686 9375
rect 39640 9329 39646 9363
rect 39680 9329 39686 9363
rect 39640 9317 39686 9329
rect 39844 9363 39890 9375
rect 39844 9329 39850 9363
rect 39884 9329 39890 9363
rect 39844 9317 39890 9329
rect 40048 9363 40094 9375
rect 40048 9329 40054 9363
rect 40088 9329 40094 9363
rect 40048 9317 40094 9329
rect 40252 9363 40298 9375
rect 40252 9329 40258 9363
rect 40292 9329 40298 9363
rect 40252 9317 40298 9329
rect 40456 9363 40502 9375
rect 40456 9329 40462 9363
rect 40496 9329 40502 9363
rect 40456 9317 40502 9329
rect 40660 9363 40706 9375
rect 40660 9329 40666 9363
rect 40700 9329 40706 9363
rect 40660 9317 40706 9329
rect 40864 9363 40910 9375
rect 40864 9329 40870 9363
rect 40904 9329 40910 9363
rect 40864 9317 40910 9329
rect 41068 9363 41114 9375
rect 41068 9329 41074 9363
rect 41108 9329 41114 9363
rect 41068 9317 41114 9329
rect 41272 9363 41318 9375
rect 41272 9329 41278 9363
rect 41312 9329 41318 9363
rect 41272 9317 41318 9329
rect 41476 9363 41522 9375
rect 41476 9329 41482 9363
rect 41516 9329 41522 9363
rect 41476 9317 41522 9329
rect 41680 9363 41726 9375
rect 41680 9329 41686 9363
rect 41720 9329 41726 9363
rect 41680 9317 41726 9329
rect 41884 9363 41930 9375
rect 41884 9329 41890 9363
rect 41924 9329 41930 9363
rect 41884 9317 41930 9329
rect 42088 9363 42134 9375
rect 42088 9329 42094 9363
rect 42128 9329 42134 9363
rect 42088 9317 42134 9329
rect 42292 9363 42338 9375
rect 42292 9329 42298 9363
rect 42332 9329 42338 9363
rect 42292 9317 42338 9329
rect 42496 9363 42542 9375
rect 42496 9329 42502 9363
rect 42536 9329 42542 9363
rect 42496 9317 42542 9329
rect 42700 9363 42746 9375
rect 42700 9329 42706 9363
rect 42740 9329 42746 9363
rect 42700 9317 42746 9329
rect 42904 9363 42950 9375
rect 42904 9329 42910 9363
rect 42944 9329 42950 9363
rect 42904 9317 42950 9329
rect 43108 9363 43154 9375
rect 43108 9329 43114 9363
rect 43148 9329 43154 9363
rect 43108 9317 43154 9329
rect 43312 9363 43358 9375
rect 43312 9329 43318 9363
rect 43352 9329 43358 9363
rect 43312 9317 43358 9329
rect 43516 9363 43562 9375
rect 43516 9329 43522 9363
rect 43556 9329 43562 9363
rect 43516 9317 43562 9329
rect 43720 9363 43766 9375
rect 43720 9329 43726 9363
rect 43760 9329 43766 9363
rect 43720 9317 43766 9329
rect 43924 9363 43970 9375
rect 43924 9329 43930 9363
rect 43964 9329 43970 9363
rect 43924 9317 43970 9329
rect 44128 9363 44174 9375
rect 44128 9329 44134 9363
rect 44168 9329 44174 9363
rect 44128 9317 44174 9329
rect 44332 9363 44378 9375
rect 44332 9329 44338 9363
rect 44372 9329 44378 9363
rect 44332 9317 44378 9329
rect 44536 9363 44582 9375
rect 44536 9329 44542 9363
rect 44576 9329 44582 9363
rect 44536 9317 44582 9329
rect 44740 9363 44786 9375
rect 44740 9329 44746 9363
rect 44780 9329 44786 9363
rect 44740 9317 44786 9329
rect 44944 9363 44990 9375
rect 44944 9329 44950 9363
rect 44984 9329 44990 9363
rect 44944 9317 44990 9329
rect 45148 9363 45194 9375
rect 45148 9329 45154 9363
rect 45188 9329 45194 9363
rect 45148 9317 45194 9329
rect 45352 9363 45398 9375
rect 45352 9329 45358 9363
rect 45392 9329 45398 9363
rect 45352 9317 45398 9329
rect 45556 9363 45602 9375
rect 45556 9329 45562 9363
rect 45596 9329 45602 9363
rect 45556 9317 45602 9329
rect 45760 9363 45806 9375
rect 45760 9329 45766 9363
rect 45800 9329 45806 9363
rect 45760 9317 45806 9329
rect 45964 9363 46010 9375
rect 45964 9329 45970 9363
rect 46004 9329 46010 9363
rect 45964 9317 46010 9329
rect 46168 9363 46214 9375
rect 46168 9329 46174 9363
rect 46208 9329 46214 9363
rect 46168 9317 46214 9329
rect 46372 9363 46418 9375
rect 46372 9329 46378 9363
rect 46412 9329 46418 9363
rect 46372 9317 46418 9329
rect 46576 9363 46622 9375
rect 46576 9329 46582 9363
rect 46616 9329 46622 9363
rect 46576 9317 46622 9329
rect 46780 9363 46826 9375
rect 46780 9329 46786 9363
rect 46820 9329 46826 9363
rect 46780 9317 46826 9329
rect 46984 9363 47030 9375
rect 46984 9329 46990 9363
rect 47024 9329 47030 9363
rect 46984 9317 47030 9329
rect 47188 9363 47234 9375
rect 47188 9329 47194 9363
rect 47228 9329 47234 9363
rect 47188 9317 47234 9329
rect 47392 9363 47438 9375
rect 47392 9329 47398 9363
rect 47432 9329 47438 9363
rect 47392 9317 47438 9329
rect 47596 9363 47642 9375
rect 47596 9329 47602 9363
rect 47636 9329 47642 9363
rect 47596 9317 47642 9329
rect 47800 9363 47846 9375
rect 47800 9329 47806 9363
rect 47840 9329 47846 9363
rect 47800 9317 47846 9329
rect 48004 9363 48050 9375
rect 48004 9329 48010 9363
rect 48044 9329 48050 9363
rect 48004 9317 48050 9329
rect 48208 9363 48254 9375
rect 48208 9329 48214 9363
rect 48248 9329 48254 9363
rect 48208 9317 48254 9329
rect 48412 9363 48458 9375
rect 48412 9329 48418 9363
rect 48452 9329 48458 9363
rect 48412 9317 48458 9329
rect 48616 9363 48662 9375
rect 48616 9329 48622 9363
rect 48656 9329 48662 9363
rect 48616 9317 48662 9329
rect 48820 9363 48866 9375
rect 48820 9329 48826 9363
rect 48860 9329 48866 9363
rect 48820 9317 48866 9329
rect 49024 9363 49070 9375
rect 49024 9329 49030 9363
rect 49064 9329 49070 9363
rect 49024 9317 49070 9329
rect 49228 9363 49274 9375
rect 49228 9329 49234 9363
rect 49268 9329 49274 9363
rect 49228 9317 49274 9329
rect 49432 9363 49478 9375
rect 49432 9329 49438 9363
rect 49472 9329 49478 9363
rect 49432 9317 49478 9329
rect 49636 9363 49682 9375
rect 49636 9329 49642 9363
rect 49676 9329 49682 9363
rect 49636 9317 49682 9329
rect 49840 9363 49886 9375
rect 49840 9329 49846 9363
rect 49880 9329 49886 9363
rect 49840 9317 49886 9329
rect 50044 9363 50090 9375
rect 50044 9329 50050 9363
rect 50084 9329 50090 9363
rect 50044 9317 50090 9329
rect 50248 9363 50294 9375
rect 50248 9329 50254 9363
rect 50288 9329 50294 9363
rect 50248 9317 50294 9329
rect 50452 9363 50498 9375
rect 50452 9329 50458 9363
rect 50492 9329 50498 9363
rect 50452 9317 50498 9329
rect 50656 9363 50702 9375
rect 50656 9329 50662 9363
rect 50696 9329 50702 9363
rect 50656 9317 50702 9329
rect 50860 9363 50906 9375
rect 50860 9329 50866 9363
rect 50900 9329 50906 9363
rect 50860 9317 50906 9329
rect 51064 9363 51110 9375
rect 51064 9329 51070 9363
rect 51104 9329 51110 9363
rect 51064 9317 51110 9329
rect 51268 9363 51314 9375
rect 51268 9329 51274 9363
rect 51308 9329 51314 9363
rect 51268 9317 51314 9329
rect 51472 9363 51518 9375
rect 51472 9329 51478 9363
rect 51512 9329 51518 9363
rect 51472 9317 51518 9329
rect 51676 9363 51722 9375
rect 51676 9329 51682 9363
rect 51716 9329 51722 9363
rect 51676 9317 51722 9329
rect 51880 9363 51926 9375
rect 51880 9329 51886 9363
rect 51920 9329 51926 9363
rect 51880 9317 51926 9329
rect 52084 9363 52130 9375
rect 52084 9329 52090 9363
rect 52124 9329 52130 9363
rect 52084 9317 52130 9329
rect 52288 9363 52334 9375
rect 52288 9329 52294 9363
rect 52328 9329 52334 9363
rect 52288 9317 52334 9329
rect 52492 9363 52538 9375
rect 52492 9329 52498 9363
rect 52532 9329 52538 9363
rect 52492 9317 52538 9329
rect 52696 9363 52742 9375
rect 52696 9329 52702 9363
rect 52736 9329 52742 9363
rect 52696 9317 52742 9329
rect 52900 9363 52946 9375
rect 52900 9329 52906 9363
rect 52940 9329 52946 9363
rect 52900 9317 52946 9329
rect 53104 9363 53150 9375
rect 53104 9329 53110 9363
rect 53144 9329 53150 9363
rect 53104 9317 53150 9329
rect 53308 9363 53354 9375
rect 53308 9329 53314 9363
rect 53348 9329 53354 9363
rect 53308 9317 53354 9329
rect 53512 9363 53558 9375
rect 53512 9329 53518 9363
rect 53552 9329 53558 9363
rect 53512 9317 53558 9329
rect 53716 9363 53762 9375
rect 53716 9329 53722 9363
rect 53756 9329 53762 9363
rect 53716 9317 53762 9329
rect 53920 9363 53966 9375
rect 53920 9329 53926 9363
rect 53960 9329 53966 9363
rect 53920 9317 53966 9329
rect 54124 9363 54170 9375
rect 54124 9329 54130 9363
rect 54164 9329 54170 9363
rect 54124 9317 54170 9329
rect 54328 9363 54374 9375
rect 54328 9329 54334 9363
rect 54368 9329 54374 9363
rect 54328 9317 54374 9329
rect 54532 9363 54578 9375
rect 54532 9329 54538 9363
rect 54572 9329 54578 9363
rect 54532 9317 54578 9329
rect 54736 9363 54782 9375
rect 54736 9329 54742 9363
rect 54776 9329 54782 9363
rect 54736 9317 54782 9329
rect 54940 9363 54986 9375
rect 54940 9329 54946 9363
rect 54980 9329 54986 9363
rect 54940 9317 54986 9329
rect 55144 9363 55190 9375
rect 55144 9329 55150 9363
rect 55184 9329 55190 9363
rect 55144 9317 55190 9329
rect 55348 9363 55394 9375
rect 55348 9329 55354 9363
rect 55388 9329 55394 9363
rect 55348 9317 55394 9329
rect 55552 9363 55598 9375
rect 55552 9329 55558 9363
rect 55592 9329 55598 9363
rect 55552 9317 55598 9329
rect 55756 9363 55802 9375
rect 55756 9329 55762 9363
rect 55796 9329 55802 9363
rect 55756 9317 55802 9329
rect 55960 9363 56006 9375
rect 55960 9329 55966 9363
rect 56000 9329 56006 9363
rect 55960 9317 56006 9329
rect 56164 9363 56210 9375
rect 56164 9329 56170 9363
rect 56204 9329 56210 9363
rect 56164 9317 56210 9329
rect 56368 9363 56414 9375
rect 56368 9329 56374 9363
rect 56408 9329 56414 9363
rect 56368 9317 56414 9329
rect 56572 9363 56618 9375
rect 56572 9329 56578 9363
rect 56612 9329 56618 9363
rect 56572 9317 56618 9329
rect 56776 9363 56822 9375
rect 56776 9329 56782 9363
rect 56816 9329 56822 9363
rect 56776 9317 56822 9329
rect 56980 9363 57026 9375
rect 56980 9329 56986 9363
rect 57020 9329 57026 9363
rect 56980 9317 57026 9329
rect 57184 9363 57230 9375
rect 57184 9329 57190 9363
rect 57224 9329 57230 9363
rect 57184 9317 57230 9329
rect 57388 9363 57434 9375
rect 57388 9329 57394 9363
rect 57428 9329 57434 9363
rect 57388 9317 57434 9329
rect 57592 9363 57638 9375
rect 57592 9329 57598 9363
rect 57632 9329 57638 9363
rect 57592 9317 57638 9329
rect 57796 9363 57842 9375
rect 57796 9329 57802 9363
rect 57836 9329 57842 9363
rect 57796 9317 57842 9329
rect 58000 9363 58046 9375
rect 58000 9329 58006 9363
rect 58040 9329 58046 9363
rect 58000 9317 58046 9329
rect 58204 9363 58250 9375
rect 58204 9329 58210 9363
rect 58244 9329 58250 9363
rect 58204 9317 58250 9329
rect 58408 9363 58454 9375
rect 58408 9329 58414 9363
rect 58448 9329 58454 9363
rect 58408 9317 58454 9329
rect 58612 9363 58658 9375
rect 58612 9329 58618 9363
rect 58652 9329 58658 9363
rect 58612 9317 58658 9329
rect 58816 9363 58862 9375
rect 58816 9329 58822 9363
rect 58856 9329 58862 9363
rect 58816 9317 58862 9329
rect 59020 9363 59066 9375
rect 59020 9329 59026 9363
rect 59060 9329 59066 9363
rect 59020 9317 59066 9329
rect 59224 9363 59270 9375
rect 59224 9329 59230 9363
rect 59264 9329 59270 9363
rect 59224 9317 59270 9329
rect 59428 9363 59474 9375
rect 59428 9329 59434 9363
rect 59468 9329 59474 9363
rect 59428 9317 59474 9329
rect 59632 9363 59678 9375
rect 59632 9329 59638 9363
rect 59672 9329 59678 9363
rect 59632 9317 59678 9329
rect 59836 9363 59882 9375
rect 59836 9329 59842 9363
rect 59876 9329 59882 9363
rect 59836 9317 59882 9329
rect 60040 9363 60086 9375
rect 60040 9329 60046 9363
rect 60080 9329 60086 9363
rect 60040 9317 60086 9329
rect 60244 9363 60290 9375
rect 60244 9329 60250 9363
rect 60284 9329 60290 9363
rect 60244 9317 60290 9329
rect 8095 8728 8101 8780
rect 8153 8728 8159 8780
rect 60319 8728 60325 8780
rect 60377 8728 60383 8780
rect 8095 7812 8101 7864
rect 8153 7812 8159 7864
rect 60319 7812 60325 7864
rect 60377 7812 60383 7864
rect 8224 7768 8270 7780
rect 8224 7734 8230 7768
rect 8264 7734 8270 7768
rect 8224 7722 8270 7734
rect 8428 7768 8474 7780
rect 8428 7734 8434 7768
rect 8468 7734 8474 7768
rect 8428 7722 8474 7734
rect 8632 7768 8678 7780
rect 8632 7734 8638 7768
rect 8672 7734 8678 7768
rect 8632 7722 8678 7734
rect 8836 7768 8882 7780
rect 8836 7734 8842 7768
rect 8876 7734 8882 7768
rect 8836 7722 8882 7734
rect 9040 7768 9086 7780
rect 9040 7734 9046 7768
rect 9080 7734 9086 7768
rect 9040 7722 9086 7734
rect 9244 7768 9290 7780
rect 9244 7734 9250 7768
rect 9284 7734 9290 7768
rect 9244 7722 9290 7734
rect 9448 7768 9494 7780
rect 9448 7734 9454 7768
rect 9488 7734 9494 7768
rect 9448 7722 9494 7734
rect 9652 7768 9698 7780
rect 9652 7734 9658 7768
rect 9692 7734 9698 7768
rect 9652 7722 9698 7734
rect 9856 7768 9902 7780
rect 9856 7734 9862 7768
rect 9896 7734 9902 7768
rect 9856 7722 9902 7734
rect 10060 7768 10106 7780
rect 10060 7734 10066 7768
rect 10100 7734 10106 7768
rect 10060 7722 10106 7734
rect 10264 7768 10310 7780
rect 10264 7734 10270 7768
rect 10304 7734 10310 7768
rect 10264 7722 10310 7734
rect 10468 7768 10514 7780
rect 10468 7734 10474 7768
rect 10508 7734 10514 7768
rect 10468 7722 10514 7734
rect 10672 7768 10718 7780
rect 10672 7734 10678 7768
rect 10712 7734 10718 7768
rect 10672 7722 10718 7734
rect 10876 7768 10922 7780
rect 10876 7734 10882 7768
rect 10916 7734 10922 7768
rect 10876 7722 10922 7734
rect 11080 7768 11126 7780
rect 11080 7734 11086 7768
rect 11120 7734 11126 7768
rect 11080 7722 11126 7734
rect 11284 7768 11330 7780
rect 11284 7734 11290 7768
rect 11324 7734 11330 7768
rect 11284 7722 11330 7734
rect 11488 7768 11534 7780
rect 11488 7734 11494 7768
rect 11528 7734 11534 7768
rect 11488 7722 11534 7734
rect 11692 7768 11738 7780
rect 11692 7734 11698 7768
rect 11732 7734 11738 7768
rect 11692 7722 11738 7734
rect 11896 7768 11942 7780
rect 11896 7734 11902 7768
rect 11936 7734 11942 7768
rect 11896 7722 11942 7734
rect 12100 7768 12146 7780
rect 12100 7734 12106 7768
rect 12140 7734 12146 7768
rect 12100 7722 12146 7734
rect 12304 7768 12350 7780
rect 12304 7734 12310 7768
rect 12344 7734 12350 7768
rect 12304 7722 12350 7734
rect 12508 7768 12554 7780
rect 12508 7734 12514 7768
rect 12548 7734 12554 7768
rect 12508 7722 12554 7734
rect 12712 7768 12758 7780
rect 12712 7734 12718 7768
rect 12752 7734 12758 7768
rect 12712 7722 12758 7734
rect 12916 7768 12962 7780
rect 12916 7734 12922 7768
rect 12956 7734 12962 7768
rect 12916 7722 12962 7734
rect 13120 7768 13166 7780
rect 13120 7734 13126 7768
rect 13160 7734 13166 7768
rect 13120 7722 13166 7734
rect 13324 7768 13370 7780
rect 13324 7734 13330 7768
rect 13364 7734 13370 7768
rect 13324 7722 13370 7734
rect 13528 7768 13574 7780
rect 13528 7734 13534 7768
rect 13568 7734 13574 7768
rect 13528 7722 13574 7734
rect 13732 7768 13778 7780
rect 13732 7734 13738 7768
rect 13772 7734 13778 7768
rect 13732 7722 13778 7734
rect 13936 7768 13982 7780
rect 13936 7734 13942 7768
rect 13976 7734 13982 7768
rect 13936 7722 13982 7734
rect 14140 7768 14186 7780
rect 14140 7734 14146 7768
rect 14180 7734 14186 7768
rect 14140 7722 14186 7734
rect 14344 7768 14390 7780
rect 14344 7734 14350 7768
rect 14384 7734 14390 7768
rect 14344 7722 14390 7734
rect 14548 7768 14594 7780
rect 14548 7734 14554 7768
rect 14588 7734 14594 7768
rect 14548 7722 14594 7734
rect 14752 7768 14798 7780
rect 14752 7734 14758 7768
rect 14792 7734 14798 7768
rect 14752 7722 14798 7734
rect 14956 7768 15002 7780
rect 14956 7734 14962 7768
rect 14996 7734 15002 7768
rect 14956 7722 15002 7734
rect 15160 7768 15206 7780
rect 15160 7734 15166 7768
rect 15200 7734 15206 7768
rect 15160 7722 15206 7734
rect 15364 7768 15410 7780
rect 15364 7734 15370 7768
rect 15404 7734 15410 7768
rect 15364 7722 15410 7734
rect 15568 7768 15614 7780
rect 15568 7734 15574 7768
rect 15608 7734 15614 7768
rect 15568 7722 15614 7734
rect 15772 7768 15818 7780
rect 15772 7734 15778 7768
rect 15812 7734 15818 7768
rect 15772 7722 15818 7734
rect 15976 7768 16022 7780
rect 15976 7734 15982 7768
rect 16016 7734 16022 7768
rect 15976 7722 16022 7734
rect 16180 7768 16226 7780
rect 16180 7734 16186 7768
rect 16220 7734 16226 7768
rect 16180 7722 16226 7734
rect 16384 7768 16430 7780
rect 16384 7734 16390 7768
rect 16424 7734 16430 7768
rect 16384 7722 16430 7734
rect 16588 7768 16634 7780
rect 16588 7734 16594 7768
rect 16628 7734 16634 7768
rect 16588 7722 16634 7734
rect 16792 7768 16838 7780
rect 16792 7734 16798 7768
rect 16832 7734 16838 7768
rect 16792 7722 16838 7734
rect 16996 7768 17042 7780
rect 16996 7734 17002 7768
rect 17036 7734 17042 7768
rect 16996 7722 17042 7734
rect 17200 7768 17246 7780
rect 17200 7734 17206 7768
rect 17240 7734 17246 7768
rect 17200 7722 17246 7734
rect 17404 7768 17450 7780
rect 17404 7734 17410 7768
rect 17444 7734 17450 7768
rect 17404 7722 17450 7734
rect 17608 7768 17654 7780
rect 17608 7734 17614 7768
rect 17648 7734 17654 7768
rect 17608 7722 17654 7734
rect 17812 7768 17858 7780
rect 17812 7734 17818 7768
rect 17852 7734 17858 7768
rect 17812 7722 17858 7734
rect 18016 7768 18062 7780
rect 18016 7734 18022 7768
rect 18056 7734 18062 7768
rect 18016 7722 18062 7734
rect 18220 7768 18266 7780
rect 18220 7734 18226 7768
rect 18260 7734 18266 7768
rect 18220 7722 18266 7734
rect 18424 7768 18470 7780
rect 18424 7734 18430 7768
rect 18464 7734 18470 7768
rect 18424 7722 18470 7734
rect 18628 7768 18674 7780
rect 18628 7734 18634 7768
rect 18668 7734 18674 7768
rect 18628 7722 18674 7734
rect 18832 7768 18878 7780
rect 18832 7734 18838 7768
rect 18872 7734 18878 7768
rect 18832 7722 18878 7734
rect 19036 7768 19082 7780
rect 19036 7734 19042 7768
rect 19076 7734 19082 7768
rect 19036 7722 19082 7734
rect 19240 7768 19286 7780
rect 19240 7734 19246 7768
rect 19280 7734 19286 7768
rect 19240 7722 19286 7734
rect 19444 7768 19490 7780
rect 19444 7734 19450 7768
rect 19484 7734 19490 7768
rect 19444 7722 19490 7734
rect 19648 7768 19694 7780
rect 19648 7734 19654 7768
rect 19688 7734 19694 7768
rect 19648 7722 19694 7734
rect 19852 7768 19898 7780
rect 19852 7734 19858 7768
rect 19892 7734 19898 7768
rect 19852 7722 19898 7734
rect 20056 7768 20102 7780
rect 20056 7734 20062 7768
rect 20096 7734 20102 7768
rect 20056 7722 20102 7734
rect 20260 7768 20306 7780
rect 20260 7734 20266 7768
rect 20300 7734 20306 7768
rect 20260 7722 20306 7734
rect 20464 7768 20510 7780
rect 20464 7734 20470 7768
rect 20504 7734 20510 7768
rect 20464 7722 20510 7734
rect 20668 7768 20714 7780
rect 20668 7734 20674 7768
rect 20708 7734 20714 7768
rect 20668 7722 20714 7734
rect 20872 7768 20918 7780
rect 20872 7734 20878 7768
rect 20912 7734 20918 7768
rect 20872 7722 20918 7734
rect 21076 7768 21122 7780
rect 21076 7734 21082 7768
rect 21116 7734 21122 7768
rect 21076 7722 21122 7734
rect 21280 7768 21326 7780
rect 21280 7734 21286 7768
rect 21320 7734 21326 7768
rect 21280 7722 21326 7734
rect 21484 7768 21530 7780
rect 21484 7734 21490 7768
rect 21524 7734 21530 7768
rect 21484 7722 21530 7734
rect 21688 7768 21734 7780
rect 21688 7734 21694 7768
rect 21728 7734 21734 7768
rect 21688 7722 21734 7734
rect 21892 7768 21938 7780
rect 21892 7734 21898 7768
rect 21932 7734 21938 7768
rect 21892 7722 21938 7734
rect 22096 7768 22142 7780
rect 22096 7734 22102 7768
rect 22136 7734 22142 7768
rect 22096 7722 22142 7734
rect 22300 7768 22346 7780
rect 22300 7734 22306 7768
rect 22340 7734 22346 7768
rect 22300 7722 22346 7734
rect 22504 7768 22550 7780
rect 22504 7734 22510 7768
rect 22544 7734 22550 7768
rect 22504 7722 22550 7734
rect 22708 7768 22754 7780
rect 22708 7734 22714 7768
rect 22748 7734 22754 7768
rect 22708 7722 22754 7734
rect 22912 7768 22958 7780
rect 22912 7734 22918 7768
rect 22952 7734 22958 7768
rect 22912 7722 22958 7734
rect 23116 7768 23162 7780
rect 23116 7734 23122 7768
rect 23156 7734 23162 7768
rect 23116 7722 23162 7734
rect 23320 7768 23366 7780
rect 23320 7734 23326 7768
rect 23360 7734 23366 7768
rect 23320 7722 23366 7734
rect 23524 7768 23570 7780
rect 23524 7734 23530 7768
rect 23564 7734 23570 7768
rect 23524 7722 23570 7734
rect 23728 7768 23774 7780
rect 23728 7734 23734 7768
rect 23768 7734 23774 7768
rect 23728 7722 23774 7734
rect 23932 7768 23978 7780
rect 23932 7734 23938 7768
rect 23972 7734 23978 7768
rect 23932 7722 23978 7734
rect 24136 7768 24182 7780
rect 24136 7734 24142 7768
rect 24176 7734 24182 7768
rect 24136 7722 24182 7734
rect 24340 7768 24386 7780
rect 24340 7734 24346 7768
rect 24380 7734 24386 7768
rect 24340 7722 24386 7734
rect 24544 7768 24590 7780
rect 24544 7734 24550 7768
rect 24584 7734 24590 7768
rect 24544 7722 24590 7734
rect 24748 7768 24794 7780
rect 24748 7734 24754 7768
rect 24788 7734 24794 7768
rect 24748 7722 24794 7734
rect 24952 7768 24998 7780
rect 24952 7734 24958 7768
rect 24992 7734 24998 7768
rect 24952 7722 24998 7734
rect 25156 7768 25202 7780
rect 25156 7734 25162 7768
rect 25196 7734 25202 7768
rect 25156 7722 25202 7734
rect 25360 7768 25406 7780
rect 25360 7734 25366 7768
rect 25400 7734 25406 7768
rect 25360 7722 25406 7734
rect 25564 7768 25610 7780
rect 25564 7734 25570 7768
rect 25604 7734 25610 7768
rect 25564 7722 25610 7734
rect 25768 7768 25814 7780
rect 25768 7734 25774 7768
rect 25808 7734 25814 7768
rect 25768 7722 25814 7734
rect 25972 7768 26018 7780
rect 25972 7734 25978 7768
rect 26012 7734 26018 7768
rect 25972 7722 26018 7734
rect 26176 7768 26222 7780
rect 26176 7734 26182 7768
rect 26216 7734 26222 7768
rect 26176 7722 26222 7734
rect 26380 7768 26426 7780
rect 26380 7734 26386 7768
rect 26420 7734 26426 7768
rect 26380 7722 26426 7734
rect 26584 7768 26630 7780
rect 26584 7734 26590 7768
rect 26624 7734 26630 7768
rect 26584 7722 26630 7734
rect 26788 7768 26834 7780
rect 26788 7734 26794 7768
rect 26828 7734 26834 7768
rect 26788 7722 26834 7734
rect 26992 7768 27038 7780
rect 26992 7734 26998 7768
rect 27032 7734 27038 7768
rect 26992 7722 27038 7734
rect 27196 7768 27242 7780
rect 27196 7734 27202 7768
rect 27236 7734 27242 7768
rect 27196 7722 27242 7734
rect 27400 7768 27446 7780
rect 27400 7734 27406 7768
rect 27440 7734 27446 7768
rect 27400 7722 27446 7734
rect 27604 7768 27650 7780
rect 27604 7734 27610 7768
rect 27644 7734 27650 7768
rect 27604 7722 27650 7734
rect 27808 7768 27854 7780
rect 27808 7734 27814 7768
rect 27848 7734 27854 7768
rect 27808 7722 27854 7734
rect 28012 7768 28058 7780
rect 28012 7734 28018 7768
rect 28052 7734 28058 7768
rect 28012 7722 28058 7734
rect 28216 7768 28262 7780
rect 28216 7734 28222 7768
rect 28256 7734 28262 7768
rect 28216 7722 28262 7734
rect 28420 7768 28466 7780
rect 28420 7734 28426 7768
rect 28460 7734 28466 7768
rect 28420 7722 28466 7734
rect 28624 7768 28670 7780
rect 28624 7734 28630 7768
rect 28664 7734 28670 7768
rect 28624 7722 28670 7734
rect 28828 7768 28874 7780
rect 28828 7734 28834 7768
rect 28868 7734 28874 7768
rect 28828 7722 28874 7734
rect 29032 7768 29078 7780
rect 29032 7734 29038 7768
rect 29072 7734 29078 7768
rect 29032 7722 29078 7734
rect 29236 7768 29282 7780
rect 29236 7734 29242 7768
rect 29276 7734 29282 7768
rect 29236 7722 29282 7734
rect 29440 7768 29486 7780
rect 29440 7734 29446 7768
rect 29480 7734 29486 7768
rect 29440 7722 29486 7734
rect 29644 7768 29690 7780
rect 29644 7734 29650 7768
rect 29684 7734 29690 7768
rect 29644 7722 29690 7734
rect 29848 7768 29894 7780
rect 29848 7734 29854 7768
rect 29888 7734 29894 7768
rect 29848 7722 29894 7734
rect 30052 7768 30098 7780
rect 30052 7734 30058 7768
rect 30092 7734 30098 7768
rect 30052 7722 30098 7734
rect 30256 7768 30302 7780
rect 30256 7734 30262 7768
rect 30296 7734 30302 7768
rect 30256 7722 30302 7734
rect 30460 7768 30506 7780
rect 30460 7734 30466 7768
rect 30500 7734 30506 7768
rect 30460 7722 30506 7734
rect 30664 7768 30710 7780
rect 30664 7734 30670 7768
rect 30704 7734 30710 7768
rect 30664 7722 30710 7734
rect 30868 7768 30914 7780
rect 30868 7734 30874 7768
rect 30908 7734 30914 7768
rect 30868 7722 30914 7734
rect 31072 7768 31118 7780
rect 31072 7734 31078 7768
rect 31112 7734 31118 7768
rect 31072 7722 31118 7734
rect 31276 7768 31322 7780
rect 31276 7734 31282 7768
rect 31316 7734 31322 7768
rect 31276 7722 31322 7734
rect 31480 7768 31526 7780
rect 31480 7734 31486 7768
rect 31520 7734 31526 7768
rect 31480 7722 31526 7734
rect 31684 7768 31730 7780
rect 31684 7734 31690 7768
rect 31724 7734 31730 7768
rect 31684 7722 31730 7734
rect 31888 7768 31934 7780
rect 31888 7734 31894 7768
rect 31928 7734 31934 7768
rect 31888 7722 31934 7734
rect 32092 7768 32138 7780
rect 32092 7734 32098 7768
rect 32132 7734 32138 7768
rect 32092 7722 32138 7734
rect 32296 7768 32342 7780
rect 32296 7734 32302 7768
rect 32336 7734 32342 7768
rect 32296 7722 32342 7734
rect 32500 7768 32546 7780
rect 32500 7734 32506 7768
rect 32540 7734 32546 7768
rect 32500 7722 32546 7734
rect 32704 7768 32750 7780
rect 32704 7734 32710 7768
rect 32744 7734 32750 7768
rect 32704 7722 32750 7734
rect 32908 7768 32954 7780
rect 32908 7734 32914 7768
rect 32948 7734 32954 7768
rect 32908 7722 32954 7734
rect 33112 7768 33158 7780
rect 33112 7734 33118 7768
rect 33152 7734 33158 7768
rect 33112 7722 33158 7734
rect 33316 7768 33362 7780
rect 33316 7734 33322 7768
rect 33356 7734 33362 7768
rect 33316 7722 33362 7734
rect 33520 7768 33566 7780
rect 33520 7734 33526 7768
rect 33560 7734 33566 7768
rect 33520 7722 33566 7734
rect 33724 7768 33770 7780
rect 33724 7734 33730 7768
rect 33764 7734 33770 7768
rect 33724 7722 33770 7734
rect 33928 7768 33974 7780
rect 33928 7734 33934 7768
rect 33968 7734 33974 7768
rect 33928 7722 33974 7734
rect 34132 7768 34178 7780
rect 34132 7734 34138 7768
rect 34172 7734 34178 7768
rect 34132 7722 34178 7734
rect 34336 7768 34382 7780
rect 34336 7734 34342 7768
rect 34376 7734 34382 7768
rect 34336 7722 34382 7734
rect 34540 7768 34586 7780
rect 34540 7734 34546 7768
rect 34580 7734 34586 7768
rect 34540 7722 34586 7734
rect 34744 7768 34790 7780
rect 34744 7734 34750 7768
rect 34784 7734 34790 7768
rect 34744 7722 34790 7734
rect 34948 7768 34994 7780
rect 34948 7734 34954 7768
rect 34988 7734 34994 7768
rect 34948 7722 34994 7734
rect 35152 7768 35198 7780
rect 35152 7734 35158 7768
rect 35192 7734 35198 7768
rect 35152 7722 35198 7734
rect 35356 7768 35402 7780
rect 35356 7734 35362 7768
rect 35396 7734 35402 7768
rect 35356 7722 35402 7734
rect 35560 7768 35606 7780
rect 35560 7734 35566 7768
rect 35600 7734 35606 7768
rect 35560 7722 35606 7734
rect 35764 7768 35810 7780
rect 35764 7734 35770 7768
rect 35804 7734 35810 7768
rect 35764 7722 35810 7734
rect 35968 7768 36014 7780
rect 35968 7734 35974 7768
rect 36008 7734 36014 7768
rect 35968 7722 36014 7734
rect 36172 7768 36218 7780
rect 36172 7734 36178 7768
rect 36212 7734 36218 7768
rect 36172 7722 36218 7734
rect 36376 7768 36422 7780
rect 36376 7734 36382 7768
rect 36416 7734 36422 7768
rect 36376 7722 36422 7734
rect 36580 7768 36626 7780
rect 36580 7734 36586 7768
rect 36620 7734 36626 7768
rect 36580 7722 36626 7734
rect 36784 7768 36830 7780
rect 36784 7734 36790 7768
rect 36824 7734 36830 7768
rect 36784 7722 36830 7734
rect 36988 7768 37034 7780
rect 36988 7734 36994 7768
rect 37028 7734 37034 7768
rect 36988 7722 37034 7734
rect 37192 7768 37238 7780
rect 37192 7734 37198 7768
rect 37232 7734 37238 7768
rect 37192 7722 37238 7734
rect 37396 7768 37442 7780
rect 37396 7734 37402 7768
rect 37436 7734 37442 7768
rect 37396 7722 37442 7734
rect 37600 7768 37646 7780
rect 37600 7734 37606 7768
rect 37640 7734 37646 7768
rect 37600 7722 37646 7734
rect 37804 7768 37850 7780
rect 37804 7734 37810 7768
rect 37844 7734 37850 7768
rect 37804 7722 37850 7734
rect 38008 7768 38054 7780
rect 38008 7734 38014 7768
rect 38048 7734 38054 7768
rect 38008 7722 38054 7734
rect 38212 7768 38258 7780
rect 38212 7734 38218 7768
rect 38252 7734 38258 7768
rect 38212 7722 38258 7734
rect 38416 7768 38462 7780
rect 38416 7734 38422 7768
rect 38456 7734 38462 7768
rect 38416 7722 38462 7734
rect 38620 7768 38666 7780
rect 38620 7734 38626 7768
rect 38660 7734 38666 7768
rect 38620 7722 38666 7734
rect 38824 7768 38870 7780
rect 38824 7734 38830 7768
rect 38864 7734 38870 7768
rect 38824 7722 38870 7734
rect 39028 7768 39074 7780
rect 39028 7734 39034 7768
rect 39068 7734 39074 7768
rect 39028 7722 39074 7734
rect 39232 7768 39278 7780
rect 39232 7734 39238 7768
rect 39272 7734 39278 7768
rect 39232 7722 39278 7734
rect 39436 7768 39482 7780
rect 39436 7734 39442 7768
rect 39476 7734 39482 7768
rect 39436 7722 39482 7734
rect 39640 7768 39686 7780
rect 39640 7734 39646 7768
rect 39680 7734 39686 7768
rect 39640 7722 39686 7734
rect 39844 7768 39890 7780
rect 39844 7734 39850 7768
rect 39884 7734 39890 7768
rect 39844 7722 39890 7734
rect 40048 7768 40094 7780
rect 40048 7734 40054 7768
rect 40088 7734 40094 7768
rect 40048 7722 40094 7734
rect 40252 7768 40298 7780
rect 40252 7734 40258 7768
rect 40292 7734 40298 7768
rect 40252 7722 40298 7734
rect 40456 7768 40502 7780
rect 40456 7734 40462 7768
rect 40496 7734 40502 7768
rect 40456 7722 40502 7734
rect 40660 7768 40706 7780
rect 40660 7734 40666 7768
rect 40700 7734 40706 7768
rect 40660 7722 40706 7734
rect 40864 7768 40910 7780
rect 40864 7734 40870 7768
rect 40904 7734 40910 7768
rect 40864 7722 40910 7734
rect 41068 7768 41114 7780
rect 41068 7734 41074 7768
rect 41108 7734 41114 7768
rect 41068 7722 41114 7734
rect 41272 7768 41318 7780
rect 41272 7734 41278 7768
rect 41312 7734 41318 7768
rect 41272 7722 41318 7734
rect 41476 7768 41522 7780
rect 41476 7734 41482 7768
rect 41516 7734 41522 7768
rect 41476 7722 41522 7734
rect 41680 7768 41726 7780
rect 41680 7734 41686 7768
rect 41720 7734 41726 7768
rect 41680 7722 41726 7734
rect 41884 7768 41930 7780
rect 41884 7734 41890 7768
rect 41924 7734 41930 7768
rect 41884 7722 41930 7734
rect 42088 7768 42134 7780
rect 42088 7734 42094 7768
rect 42128 7734 42134 7768
rect 42088 7722 42134 7734
rect 42292 7768 42338 7780
rect 42292 7734 42298 7768
rect 42332 7734 42338 7768
rect 42292 7722 42338 7734
rect 42496 7768 42542 7780
rect 42496 7734 42502 7768
rect 42536 7734 42542 7768
rect 42496 7722 42542 7734
rect 42700 7768 42746 7780
rect 42700 7734 42706 7768
rect 42740 7734 42746 7768
rect 42700 7722 42746 7734
rect 42904 7768 42950 7780
rect 42904 7734 42910 7768
rect 42944 7734 42950 7768
rect 42904 7722 42950 7734
rect 43108 7768 43154 7780
rect 43108 7734 43114 7768
rect 43148 7734 43154 7768
rect 43108 7722 43154 7734
rect 43312 7768 43358 7780
rect 43312 7734 43318 7768
rect 43352 7734 43358 7768
rect 43312 7722 43358 7734
rect 43516 7768 43562 7780
rect 43516 7734 43522 7768
rect 43556 7734 43562 7768
rect 43516 7722 43562 7734
rect 43720 7768 43766 7780
rect 43720 7734 43726 7768
rect 43760 7734 43766 7768
rect 43720 7722 43766 7734
rect 43924 7768 43970 7780
rect 43924 7734 43930 7768
rect 43964 7734 43970 7768
rect 43924 7722 43970 7734
rect 44128 7768 44174 7780
rect 44128 7734 44134 7768
rect 44168 7734 44174 7768
rect 44128 7722 44174 7734
rect 44332 7768 44378 7780
rect 44332 7734 44338 7768
rect 44372 7734 44378 7768
rect 44332 7722 44378 7734
rect 44536 7768 44582 7780
rect 44536 7734 44542 7768
rect 44576 7734 44582 7768
rect 44536 7722 44582 7734
rect 44740 7768 44786 7780
rect 44740 7734 44746 7768
rect 44780 7734 44786 7768
rect 44740 7722 44786 7734
rect 44944 7768 44990 7780
rect 44944 7734 44950 7768
rect 44984 7734 44990 7768
rect 44944 7722 44990 7734
rect 45148 7768 45194 7780
rect 45148 7734 45154 7768
rect 45188 7734 45194 7768
rect 45148 7722 45194 7734
rect 45352 7768 45398 7780
rect 45352 7734 45358 7768
rect 45392 7734 45398 7768
rect 45352 7722 45398 7734
rect 45556 7768 45602 7780
rect 45556 7734 45562 7768
rect 45596 7734 45602 7768
rect 45556 7722 45602 7734
rect 45760 7768 45806 7780
rect 45760 7734 45766 7768
rect 45800 7734 45806 7768
rect 45760 7722 45806 7734
rect 45964 7768 46010 7780
rect 45964 7734 45970 7768
rect 46004 7734 46010 7768
rect 45964 7722 46010 7734
rect 46168 7768 46214 7780
rect 46168 7734 46174 7768
rect 46208 7734 46214 7768
rect 46168 7722 46214 7734
rect 46372 7768 46418 7780
rect 46372 7734 46378 7768
rect 46412 7734 46418 7768
rect 46372 7722 46418 7734
rect 46576 7768 46622 7780
rect 46576 7734 46582 7768
rect 46616 7734 46622 7768
rect 46576 7722 46622 7734
rect 46780 7768 46826 7780
rect 46780 7734 46786 7768
rect 46820 7734 46826 7768
rect 46780 7722 46826 7734
rect 46984 7768 47030 7780
rect 46984 7734 46990 7768
rect 47024 7734 47030 7768
rect 46984 7722 47030 7734
rect 47188 7768 47234 7780
rect 47188 7734 47194 7768
rect 47228 7734 47234 7768
rect 47188 7722 47234 7734
rect 47392 7768 47438 7780
rect 47392 7734 47398 7768
rect 47432 7734 47438 7768
rect 47392 7722 47438 7734
rect 47596 7768 47642 7780
rect 47596 7734 47602 7768
rect 47636 7734 47642 7768
rect 47596 7722 47642 7734
rect 47800 7768 47846 7780
rect 47800 7734 47806 7768
rect 47840 7734 47846 7768
rect 47800 7722 47846 7734
rect 48004 7768 48050 7780
rect 48004 7734 48010 7768
rect 48044 7734 48050 7768
rect 48004 7722 48050 7734
rect 48208 7768 48254 7780
rect 48208 7734 48214 7768
rect 48248 7734 48254 7768
rect 48208 7722 48254 7734
rect 48412 7768 48458 7780
rect 48412 7734 48418 7768
rect 48452 7734 48458 7768
rect 48412 7722 48458 7734
rect 48616 7768 48662 7780
rect 48616 7734 48622 7768
rect 48656 7734 48662 7768
rect 48616 7722 48662 7734
rect 48820 7768 48866 7780
rect 48820 7734 48826 7768
rect 48860 7734 48866 7768
rect 48820 7722 48866 7734
rect 49024 7768 49070 7780
rect 49024 7734 49030 7768
rect 49064 7734 49070 7768
rect 49024 7722 49070 7734
rect 49228 7768 49274 7780
rect 49228 7734 49234 7768
rect 49268 7734 49274 7768
rect 49228 7722 49274 7734
rect 49432 7768 49478 7780
rect 49432 7734 49438 7768
rect 49472 7734 49478 7768
rect 49432 7722 49478 7734
rect 49636 7768 49682 7780
rect 49636 7734 49642 7768
rect 49676 7734 49682 7768
rect 49636 7722 49682 7734
rect 49840 7768 49886 7780
rect 49840 7734 49846 7768
rect 49880 7734 49886 7768
rect 49840 7722 49886 7734
rect 50044 7768 50090 7780
rect 50044 7734 50050 7768
rect 50084 7734 50090 7768
rect 50044 7722 50090 7734
rect 50248 7768 50294 7780
rect 50248 7734 50254 7768
rect 50288 7734 50294 7768
rect 50248 7722 50294 7734
rect 50452 7768 50498 7780
rect 50452 7734 50458 7768
rect 50492 7734 50498 7768
rect 50452 7722 50498 7734
rect 50656 7768 50702 7780
rect 50656 7734 50662 7768
rect 50696 7734 50702 7768
rect 50656 7722 50702 7734
rect 50860 7768 50906 7780
rect 50860 7734 50866 7768
rect 50900 7734 50906 7768
rect 50860 7722 50906 7734
rect 51064 7768 51110 7780
rect 51064 7734 51070 7768
rect 51104 7734 51110 7768
rect 51064 7722 51110 7734
rect 51268 7768 51314 7780
rect 51268 7734 51274 7768
rect 51308 7734 51314 7768
rect 51268 7722 51314 7734
rect 51472 7768 51518 7780
rect 51472 7734 51478 7768
rect 51512 7734 51518 7768
rect 51472 7722 51518 7734
rect 51676 7768 51722 7780
rect 51676 7734 51682 7768
rect 51716 7734 51722 7768
rect 51676 7722 51722 7734
rect 51880 7768 51926 7780
rect 51880 7734 51886 7768
rect 51920 7734 51926 7768
rect 51880 7722 51926 7734
rect 52084 7768 52130 7780
rect 52084 7734 52090 7768
rect 52124 7734 52130 7768
rect 52084 7722 52130 7734
rect 52288 7768 52334 7780
rect 52288 7734 52294 7768
rect 52328 7734 52334 7768
rect 52288 7722 52334 7734
rect 52492 7768 52538 7780
rect 52492 7734 52498 7768
rect 52532 7734 52538 7768
rect 52492 7722 52538 7734
rect 52696 7768 52742 7780
rect 52696 7734 52702 7768
rect 52736 7734 52742 7768
rect 52696 7722 52742 7734
rect 52900 7768 52946 7780
rect 52900 7734 52906 7768
rect 52940 7734 52946 7768
rect 52900 7722 52946 7734
rect 53104 7768 53150 7780
rect 53104 7734 53110 7768
rect 53144 7734 53150 7768
rect 53104 7722 53150 7734
rect 53308 7768 53354 7780
rect 53308 7734 53314 7768
rect 53348 7734 53354 7768
rect 53308 7722 53354 7734
rect 53512 7768 53558 7780
rect 53512 7734 53518 7768
rect 53552 7734 53558 7768
rect 53512 7722 53558 7734
rect 53716 7768 53762 7780
rect 53716 7734 53722 7768
rect 53756 7734 53762 7768
rect 53716 7722 53762 7734
rect 53920 7768 53966 7780
rect 53920 7734 53926 7768
rect 53960 7734 53966 7768
rect 53920 7722 53966 7734
rect 54124 7768 54170 7780
rect 54124 7734 54130 7768
rect 54164 7734 54170 7768
rect 54124 7722 54170 7734
rect 54328 7768 54374 7780
rect 54328 7734 54334 7768
rect 54368 7734 54374 7768
rect 54328 7722 54374 7734
rect 54532 7768 54578 7780
rect 54532 7734 54538 7768
rect 54572 7734 54578 7768
rect 54532 7722 54578 7734
rect 54736 7768 54782 7780
rect 54736 7734 54742 7768
rect 54776 7734 54782 7768
rect 54736 7722 54782 7734
rect 54940 7768 54986 7780
rect 54940 7734 54946 7768
rect 54980 7734 54986 7768
rect 54940 7722 54986 7734
rect 55144 7768 55190 7780
rect 55144 7734 55150 7768
rect 55184 7734 55190 7768
rect 55144 7722 55190 7734
rect 55348 7768 55394 7780
rect 55348 7734 55354 7768
rect 55388 7734 55394 7768
rect 55348 7722 55394 7734
rect 55552 7768 55598 7780
rect 55552 7734 55558 7768
rect 55592 7734 55598 7768
rect 55552 7722 55598 7734
rect 55756 7768 55802 7780
rect 55756 7734 55762 7768
rect 55796 7734 55802 7768
rect 55756 7722 55802 7734
rect 55960 7768 56006 7780
rect 55960 7734 55966 7768
rect 56000 7734 56006 7768
rect 55960 7722 56006 7734
rect 56164 7768 56210 7780
rect 56164 7734 56170 7768
rect 56204 7734 56210 7768
rect 56164 7722 56210 7734
rect 56368 7768 56414 7780
rect 56368 7734 56374 7768
rect 56408 7734 56414 7768
rect 56368 7722 56414 7734
rect 56572 7768 56618 7780
rect 56572 7734 56578 7768
rect 56612 7734 56618 7768
rect 56572 7722 56618 7734
rect 56776 7768 56822 7780
rect 56776 7734 56782 7768
rect 56816 7734 56822 7768
rect 56776 7722 56822 7734
rect 56980 7768 57026 7780
rect 56980 7734 56986 7768
rect 57020 7734 57026 7768
rect 56980 7722 57026 7734
rect 57184 7768 57230 7780
rect 57184 7734 57190 7768
rect 57224 7734 57230 7768
rect 57184 7722 57230 7734
rect 57388 7768 57434 7780
rect 57388 7734 57394 7768
rect 57428 7734 57434 7768
rect 57388 7722 57434 7734
rect 57592 7768 57638 7780
rect 57592 7734 57598 7768
rect 57632 7734 57638 7768
rect 57592 7722 57638 7734
rect 57796 7768 57842 7780
rect 57796 7734 57802 7768
rect 57836 7734 57842 7768
rect 57796 7722 57842 7734
rect 58000 7768 58046 7780
rect 58000 7734 58006 7768
rect 58040 7734 58046 7768
rect 58000 7722 58046 7734
rect 58204 7768 58250 7780
rect 58204 7734 58210 7768
rect 58244 7734 58250 7768
rect 58204 7722 58250 7734
rect 58408 7768 58454 7780
rect 58408 7734 58414 7768
rect 58448 7734 58454 7768
rect 58408 7722 58454 7734
rect 58612 7768 58658 7780
rect 58612 7734 58618 7768
rect 58652 7734 58658 7768
rect 58612 7722 58658 7734
rect 58816 7768 58862 7780
rect 58816 7734 58822 7768
rect 58856 7734 58862 7768
rect 58816 7722 58862 7734
rect 59020 7768 59066 7780
rect 59020 7734 59026 7768
rect 59060 7734 59066 7768
rect 59020 7722 59066 7734
rect 59224 7768 59270 7780
rect 59224 7734 59230 7768
rect 59264 7734 59270 7768
rect 59224 7722 59270 7734
rect 59428 7768 59474 7780
rect 59428 7734 59434 7768
rect 59468 7734 59474 7768
rect 59428 7722 59474 7734
rect 59632 7768 59678 7780
rect 59632 7734 59638 7768
rect 59672 7734 59678 7768
rect 59632 7722 59678 7734
rect 59836 7768 59882 7780
rect 59836 7734 59842 7768
rect 59876 7734 59882 7768
rect 59836 7722 59882 7734
rect 60040 7768 60086 7780
rect 60040 7734 60046 7768
rect 60080 7734 60086 7768
rect 60040 7722 60086 7734
rect 60244 7768 60290 7780
rect 60244 7734 60250 7768
rect 60284 7734 60290 7768
rect 60244 7722 60290 7734
rect 8233 7216 8261 7722
rect 8437 7216 8465 7722
rect 8641 7216 8669 7722
rect 8845 7216 8873 7722
rect 9049 7216 9077 7722
rect 9253 7216 9281 7722
rect 9457 7216 9485 7722
rect 9661 7216 9689 7722
rect 9865 7216 9893 7722
rect 10069 7216 10097 7722
rect 10273 7216 10301 7722
rect 10477 7216 10505 7722
rect 10681 7216 10709 7722
rect 10885 7216 10913 7722
rect 11089 7216 11117 7722
rect 11293 7216 11321 7722
rect 11497 7216 11525 7722
rect 11701 7216 11729 7722
rect 11905 7216 11933 7722
rect 12109 7216 12137 7722
rect 12313 7216 12341 7722
rect 12517 7216 12545 7722
rect 12721 7216 12749 7722
rect 12925 7216 12953 7722
rect 13129 7216 13157 7722
rect 13333 7216 13361 7722
rect 13537 7216 13565 7722
rect 13741 7216 13769 7722
rect 13945 7216 13973 7722
rect 14149 7216 14177 7722
rect 14353 7216 14381 7722
rect 14557 7216 14585 7722
rect 14761 7216 14789 7722
rect 14965 7216 14993 7722
rect 15169 7216 15197 7722
rect 15373 7216 15401 7722
rect 15577 7216 15605 7722
rect 15781 7216 15809 7722
rect 15985 7216 16013 7722
rect 16189 7216 16217 7722
rect 16393 7216 16421 7722
rect 16597 7216 16625 7722
rect 16801 7216 16829 7722
rect 17005 7216 17033 7722
rect 17209 7216 17237 7722
rect 17413 7216 17441 7722
rect 17617 7216 17645 7722
rect 17821 7216 17849 7722
rect 18025 7216 18053 7722
rect 18229 7216 18257 7722
rect 18433 7216 18461 7722
rect 18637 7216 18665 7722
rect 18841 7216 18869 7722
rect 19045 7216 19073 7722
rect 19249 7216 19277 7722
rect 19453 7216 19481 7722
rect 19657 7216 19685 7722
rect 19861 7216 19889 7722
rect 20065 7216 20093 7722
rect 20269 7216 20297 7722
rect 20473 7216 20501 7722
rect 20677 7216 20705 7722
rect 20881 7216 20909 7722
rect 21085 7216 21113 7722
rect 21289 7216 21317 7722
rect 21493 7216 21521 7722
rect 21697 7216 21725 7722
rect 21901 7216 21929 7722
rect 22105 7216 22133 7722
rect 22309 7216 22337 7722
rect 22513 7216 22541 7722
rect 22717 7216 22745 7722
rect 22921 7216 22949 7722
rect 23125 7216 23153 7722
rect 23329 7216 23357 7722
rect 23533 7216 23561 7722
rect 23737 7216 23765 7722
rect 23941 7216 23969 7722
rect 24145 7216 24173 7722
rect 24349 7216 24377 7722
rect 24553 7216 24581 7722
rect 24757 7216 24785 7722
rect 24961 7216 24989 7722
rect 25165 7216 25193 7722
rect 25369 7216 25397 7722
rect 25573 7216 25601 7722
rect 25777 7216 25805 7722
rect 25981 7216 26009 7722
rect 26185 7216 26213 7722
rect 26389 7216 26417 7722
rect 26593 7216 26621 7722
rect 26797 7216 26825 7722
rect 27001 7216 27029 7722
rect 27205 7216 27233 7722
rect 27409 7216 27437 7722
rect 27613 7216 27641 7722
rect 27817 7216 27845 7722
rect 28021 7216 28049 7722
rect 28225 7216 28253 7722
rect 28429 7216 28457 7722
rect 28633 7216 28661 7722
rect 28837 7216 28865 7722
rect 29041 7216 29069 7722
rect 29245 7216 29273 7722
rect 29449 7216 29477 7722
rect 29653 7216 29681 7722
rect 29857 7216 29885 7722
rect 30061 7216 30089 7722
rect 30265 7216 30293 7722
rect 30469 7216 30497 7722
rect 30673 7216 30701 7722
rect 30877 7216 30905 7722
rect 31081 7216 31109 7722
rect 31285 7216 31313 7722
rect 31489 7216 31517 7722
rect 31693 7216 31721 7722
rect 31897 7216 31925 7722
rect 32101 7216 32129 7722
rect 32305 7216 32333 7722
rect 32509 7216 32537 7722
rect 32713 7216 32741 7722
rect 32917 7216 32945 7722
rect 33121 7216 33149 7722
rect 33325 7216 33353 7722
rect 33529 7216 33557 7722
rect 33733 7216 33761 7722
rect 33937 7216 33965 7722
rect 34141 7216 34169 7722
rect 34345 7216 34373 7722
rect 34549 7216 34577 7722
rect 34753 7216 34781 7722
rect 34957 7216 34985 7722
rect 35161 7216 35189 7722
rect 35365 7216 35393 7722
rect 35569 7216 35597 7722
rect 35773 7216 35801 7722
rect 35977 7216 36005 7722
rect 36181 7216 36209 7722
rect 36385 7216 36413 7722
rect 36589 7216 36617 7722
rect 36793 7216 36821 7722
rect 36997 7216 37025 7722
rect 37201 7216 37229 7722
rect 37405 7216 37433 7722
rect 37609 7216 37637 7722
rect 37813 7216 37841 7722
rect 38017 7216 38045 7722
rect 38221 7216 38249 7722
rect 38425 7216 38453 7722
rect 38629 7216 38657 7722
rect 38833 7216 38861 7722
rect 39037 7216 39065 7722
rect 39241 7216 39269 7722
rect 39445 7216 39473 7722
rect 39649 7216 39677 7722
rect 39853 7216 39881 7722
rect 40057 7216 40085 7722
rect 40261 7216 40289 7722
rect 40465 7216 40493 7722
rect 40669 7216 40697 7722
rect 40873 7216 40901 7722
rect 41077 7216 41105 7722
rect 41281 7216 41309 7722
rect 41485 7216 41513 7722
rect 41689 7216 41717 7722
rect 41893 7216 41921 7722
rect 42097 7216 42125 7722
rect 42301 7216 42329 7722
rect 42505 7216 42533 7722
rect 42709 7216 42737 7722
rect 42913 7216 42941 7722
rect 43117 7216 43145 7722
rect 43321 7216 43349 7722
rect 43525 7216 43553 7722
rect 43729 7216 43757 7722
rect 43933 7216 43961 7722
rect 44137 7216 44165 7722
rect 44341 7216 44369 7722
rect 44545 7216 44573 7722
rect 44749 7216 44777 7722
rect 44953 7216 44981 7722
rect 45157 7216 45185 7722
rect 45361 7216 45389 7722
rect 45565 7216 45593 7722
rect 45769 7216 45797 7722
rect 45973 7216 46001 7722
rect 46177 7216 46205 7722
rect 46381 7216 46409 7722
rect 46585 7216 46613 7722
rect 46789 7216 46817 7722
rect 46993 7216 47021 7722
rect 47197 7216 47225 7722
rect 47401 7216 47429 7722
rect 47605 7216 47633 7722
rect 47809 7216 47837 7722
rect 48013 7216 48041 7722
rect 48217 7216 48245 7722
rect 48421 7216 48449 7722
rect 48625 7216 48653 7722
rect 48829 7216 48857 7722
rect 49033 7216 49061 7722
rect 49237 7216 49265 7722
rect 49441 7216 49469 7722
rect 49645 7216 49673 7722
rect 49849 7216 49877 7722
rect 50053 7216 50081 7722
rect 50257 7216 50285 7722
rect 50461 7216 50489 7722
rect 50665 7216 50693 7722
rect 50869 7216 50897 7722
rect 51073 7216 51101 7722
rect 51277 7216 51305 7722
rect 51481 7216 51509 7722
rect 51685 7216 51713 7722
rect 51889 7216 51917 7722
rect 52093 7216 52121 7722
rect 52297 7216 52325 7722
rect 52501 7216 52529 7722
rect 52705 7216 52733 7722
rect 52909 7216 52937 7722
rect 53113 7216 53141 7722
rect 53317 7216 53345 7722
rect 53521 7216 53549 7722
rect 53725 7216 53753 7722
rect 53929 7216 53957 7722
rect 54133 7216 54161 7722
rect 54337 7216 54365 7722
rect 54541 7216 54569 7722
rect 54745 7216 54773 7722
rect 54949 7216 54977 7722
rect 55153 7216 55181 7722
rect 55357 7216 55385 7722
rect 55561 7216 55589 7722
rect 55765 7216 55793 7722
rect 55969 7216 55997 7722
rect 56173 7216 56201 7722
rect 56377 7216 56405 7722
rect 56581 7216 56609 7722
rect 56785 7216 56813 7722
rect 56989 7216 57017 7722
rect 57193 7216 57221 7722
rect 57397 7216 57425 7722
rect 57601 7216 57629 7722
rect 57805 7216 57833 7722
rect 58009 7216 58037 7722
rect 58213 7216 58241 7722
rect 58417 7216 58445 7722
rect 58621 7216 58649 7722
rect 58825 7216 58853 7722
rect 59029 7216 59057 7722
rect 59233 7216 59261 7722
rect 59437 7216 59465 7722
rect 59641 7216 59669 7722
rect 59845 7216 59873 7722
rect 60049 7216 60077 7722
rect 60253 7216 60281 7722
rect 4278 6759 6403 6787
rect 2981 5622 3039 5628
rect 2981 5588 2993 5622
rect 3027 5619 3039 5622
rect 4278 5619 4306 6759
rect 7003 6490 7009 6542
rect 7061 6490 7067 6542
rect 7625 6490 7631 6542
rect 7683 6490 7689 6542
rect 7944 6370 7950 6422
rect 8002 6370 8008 6422
rect 7944 6166 7950 6218
rect 8002 6166 8008 6218
rect 7944 5962 7950 6014
rect 8002 5962 8008 6014
rect 7944 5758 7950 5810
rect 8002 5758 8008 5810
rect 3027 5591 4306 5619
rect 3027 5588 3039 5591
rect 2981 5582 3039 5588
rect 4278 3718 4306 5591
rect 7944 5554 7950 5606
rect 8002 5554 8008 5606
rect 7944 5350 7950 5402
rect 8002 5350 8008 5402
rect 7944 5146 7950 5198
rect 8002 5146 8008 5198
rect 7944 4942 7950 4994
rect 8002 4942 8008 4994
rect 7003 4774 7009 4826
rect 7061 4774 7067 4826
rect 7625 4774 7631 4826
rect 7683 4774 7689 4826
rect 8215 4724 8221 4776
rect 8273 4724 8279 4776
rect 9847 4724 9853 4776
rect 9905 4724 9911 4776
rect 11479 4724 11485 4776
rect 11537 4724 11543 4776
rect 13111 4724 13117 4776
rect 13169 4724 13175 4776
rect 14743 4724 14749 4776
rect 14801 4724 14807 4776
rect 16375 4724 16381 4776
rect 16433 4724 16439 4776
rect 18007 4724 18013 4776
rect 18065 4724 18071 4776
rect 19639 4724 19645 4776
rect 19697 4724 19703 4776
rect 21271 4724 21277 4776
rect 21329 4724 21335 4776
rect 22903 4724 22909 4776
rect 22961 4724 22967 4776
rect 24535 4724 24541 4776
rect 24593 4724 24599 4776
rect 26167 4724 26173 4776
rect 26225 4724 26231 4776
rect 27799 4724 27805 4776
rect 27857 4724 27863 4776
rect 29431 4724 29437 4776
rect 29489 4724 29495 4776
rect 31063 4724 31069 4776
rect 31121 4724 31127 4776
rect 32695 4724 32701 4776
rect 32753 4724 32759 4776
rect 34327 4724 34333 4776
rect 34385 4724 34391 4776
rect 35959 4724 35965 4776
rect 36017 4724 36023 4776
rect 37591 4724 37597 4776
rect 37649 4724 37655 4776
rect 39223 4724 39229 4776
rect 39281 4724 39287 4776
rect 40855 4724 40861 4776
rect 40913 4724 40919 4776
rect 42487 4724 42493 4776
rect 42545 4724 42551 4776
rect 44119 4724 44125 4776
rect 44177 4724 44183 4776
rect 45751 4724 45757 4776
rect 45809 4724 45815 4776
rect 47383 4724 47389 4776
rect 47441 4724 47447 4776
rect 49015 4724 49021 4776
rect 49073 4724 49079 4776
rect 50647 4724 50653 4776
rect 50705 4724 50711 4776
rect 52279 4724 52285 4776
rect 52337 4724 52343 4776
rect 53911 4724 53917 4776
rect 53969 4724 53975 4776
rect 55543 4724 55549 4776
rect 55601 4724 55607 4776
rect 57175 4724 57181 4776
rect 57233 4724 57239 4776
rect 58807 4724 58813 4776
rect 58865 4724 58871 4776
rect 4607 4351 4613 4403
rect 4665 4351 4671 4403
rect 24225 4061 24231 4113
rect 24283 4101 24289 4113
rect 58807 4101 58813 4113
rect 24283 4073 58813 4101
rect 24283 4061 24289 4073
rect 58807 4061 58813 4073
rect 58865 4061 58871 4113
rect 5831 3926 5837 3978
rect 5889 3926 5895 3978
rect 23917 3959 23923 4011
rect 23975 3999 23981 4011
rect 57175 3999 57181 4011
rect 23975 3971 57181 3999
rect 23975 3959 23981 3971
rect 57175 3959 57181 3971
rect 57233 3959 57239 4011
rect 23609 3857 23615 3909
rect 23667 3897 23673 3909
rect 55543 3897 55549 3909
rect 23667 3869 55549 3897
rect 23667 3857 23673 3869
rect 55543 3857 55549 3869
rect 55601 3857 55607 3909
rect 17449 3755 17455 3807
rect 17507 3795 17513 3807
rect 22903 3795 22909 3807
rect 17507 3767 22909 3795
rect 17507 3755 17513 3767
rect 22903 3755 22909 3767
rect 22961 3755 22967 3807
rect 23301 3755 23307 3807
rect 23359 3795 23365 3807
rect 53911 3795 53917 3807
rect 23359 3767 53917 3795
rect 23359 3755 23365 3767
rect 53911 3755 53917 3767
rect 53969 3755 53975 3807
rect 4278 3690 5237 3718
rect 22993 3653 22999 3705
rect 23051 3693 23057 3705
rect 52279 3693 52285 3705
rect 23051 3665 52285 3693
rect 23051 3653 23057 3665
rect 52279 3653 52285 3665
rect 52337 3653 52343 3705
rect 22685 3551 22691 3603
rect 22743 3591 22749 3603
rect 50647 3591 50653 3603
rect 22743 3563 50653 3591
rect 22743 3551 22749 3563
rect 50647 3551 50653 3563
rect 50705 3551 50711 3603
rect 4607 3399 4613 3451
rect 4665 3399 4671 3451
rect 22377 3449 22383 3501
rect 22435 3489 22441 3501
rect 49015 3489 49021 3501
rect 22435 3461 49021 3489
rect 22435 3449 22441 3461
rect 49015 3449 49021 3461
rect 49073 3449 49079 3501
rect 22069 3347 22075 3399
rect 22127 3387 22133 3399
rect 47383 3387 47389 3399
rect 22127 3359 47389 3387
rect 22127 3347 22133 3359
rect 47383 3347 47389 3359
rect 47441 3347 47447 3399
rect 21761 3245 21767 3297
rect 21819 3285 21825 3297
rect 45751 3285 45757 3297
rect 21819 3257 45757 3285
rect 21819 3245 21825 3257
rect 45751 3245 45757 3257
rect 45809 3245 45815 3297
rect 21145 3143 21151 3195
rect 21203 3183 21209 3195
rect 42487 3183 42493 3195
rect 21203 3155 42493 3183
rect 21203 3143 21209 3155
rect 42487 3143 42493 3155
rect 42545 3143 42551 3195
rect 20837 3041 20843 3093
rect 20895 3081 20901 3093
rect 40855 3081 40861 3093
rect 20895 3053 40861 3081
rect 20895 3041 20901 3053
rect 40855 3041 40861 3053
rect 40913 3041 40919 3093
rect -1401 2914 -1395 2966
rect -1343 2914 -1337 2966
rect 36 2952 42 3004
rect 94 2952 100 3004
rect 5831 2974 5837 3026
rect 5889 2974 5895 3026
rect 20529 2939 20535 2991
rect 20587 2979 20593 2991
rect 39223 2979 39229 2991
rect 20587 2951 39229 2979
rect 20587 2939 20593 2951
rect 39223 2939 39229 2951
rect 39281 2939 39287 2991
rect 20221 2837 20227 2889
rect 20279 2877 20285 2889
rect 37591 2877 37597 2889
rect 20279 2849 37597 2877
rect 20279 2837 20285 2849
rect 37591 2837 37597 2849
rect 37649 2837 37655 2889
rect 16833 2735 16839 2787
rect 16891 2775 16897 2787
rect 19639 2775 19645 2787
rect 16891 2747 19645 2775
rect 16891 2735 16897 2747
rect 19639 2735 19645 2747
rect 19697 2735 19703 2787
rect 19913 2735 19919 2787
rect 19971 2775 19977 2787
rect 35959 2775 35965 2787
rect 19971 2747 35965 2775
rect 19971 2735 19977 2747
rect 35959 2735 35965 2747
rect 36017 2735 36023 2787
rect 19605 2633 19611 2685
rect 19663 2673 19669 2685
rect 34327 2673 34333 2685
rect 19663 2645 34333 2673
rect 19663 2633 19669 2645
rect 34327 2633 34333 2645
rect 34385 2633 34391 2685
rect 19297 2531 19303 2583
rect 19355 2571 19361 2583
rect 32695 2571 32701 2583
rect 19355 2543 32701 2571
rect 19355 2531 19361 2543
rect 32695 2531 32701 2543
rect 32753 2531 32759 2583
rect 18989 2429 18995 2481
rect 19047 2469 19053 2481
rect 31063 2469 31069 2481
rect 19047 2441 31069 2469
rect 19047 2429 19053 2441
rect 31063 2429 31069 2441
rect 31121 2429 31127 2481
rect 4607 2362 4613 2414
rect 4665 2362 4671 2414
rect 14743 2327 14749 2379
rect 14801 2367 14807 2379
rect 15909 2367 15915 2379
rect 14801 2339 15915 2367
rect 14801 2327 14807 2339
rect 15909 2327 15915 2339
rect 15967 2327 15973 2379
rect 18681 2327 18687 2379
rect 18739 2367 18745 2379
rect 29431 2367 29437 2379
rect 18739 2339 29437 2367
rect 18739 2327 18745 2339
rect 29431 2327 29437 2339
rect 29489 2327 29495 2379
rect 13111 2225 13117 2277
rect 13169 2265 13175 2277
rect 15601 2265 15607 2277
rect 13169 2237 15607 2265
rect 13169 2225 13175 2237
rect 15601 2225 15607 2237
rect 15659 2225 15665 2277
rect 16525 2225 16531 2277
rect 16583 2265 16589 2277
rect 18007 2265 18013 2277
rect 16583 2237 18013 2265
rect 16583 2225 16589 2237
rect 18007 2225 18013 2237
rect 18065 2225 18071 2277
rect 18373 2225 18379 2277
rect 18431 2265 18437 2277
rect 27799 2265 27805 2277
rect 18431 2237 27805 2265
rect 18431 2225 18437 2237
rect 27799 2225 27805 2237
rect 27857 2225 27863 2277
rect 11479 2123 11485 2175
rect 11537 2163 11543 2175
rect 15293 2163 15299 2175
rect 11537 2135 15299 2163
rect 11537 2123 11543 2135
rect 15293 2123 15299 2135
rect 15351 2123 15357 2175
rect 18065 2123 18071 2175
rect 18123 2163 18129 2175
rect 26167 2163 26173 2175
rect 18123 2135 26173 2163
rect 18123 2123 18129 2135
rect 26167 2123 26173 2135
rect 26225 2123 26231 2175
rect 9847 2021 9853 2073
rect 9905 2061 9911 2073
rect 14985 2061 14991 2073
rect 9905 2033 14991 2061
rect 9905 2021 9911 2033
rect 14985 2021 14991 2033
rect 15043 2021 15049 2073
rect 17757 2021 17763 2073
rect 17815 2061 17821 2073
rect 24535 2061 24541 2073
rect 17815 2033 24541 2061
rect 17815 2021 17821 2033
rect 24535 2021 24541 2033
rect 24593 2021 24599 2073
rect 443 1907 449 1959
rect 501 1907 507 1959
rect 8215 1919 8221 1971
rect 8273 1959 8279 1971
rect 14677 1959 14683 1971
rect 8273 1931 14683 1959
rect 8273 1919 8279 1931
rect 14677 1919 14683 1931
rect 14735 1919 14741 1971
rect 16217 1919 16223 1971
rect 16275 1959 16281 1971
rect 16375 1959 16381 1971
rect 16275 1931 16381 1959
rect 16275 1919 16281 1931
rect 16375 1919 16381 1931
rect 16433 1919 16439 1971
rect 17141 1919 17147 1971
rect 17199 1959 17205 1971
rect 21271 1959 21277 1971
rect 17199 1931 21277 1959
rect 17199 1919 17205 1931
rect 21271 1919 21277 1931
rect 21329 1919 21335 1971
rect 21453 1919 21459 1971
rect 21511 1959 21517 1971
rect 44119 1959 44125 1971
rect 21511 1931 44125 1959
rect 21511 1919 21517 1931
rect 44119 1919 44125 1931
rect 44177 1919 44183 1971
rect 5831 1740 5837 1792
rect 5889 1740 5895 1792
rect 14677 1696 14683 1748
rect 14735 1696 14741 1748
rect 14985 1696 14991 1748
rect 15043 1696 15049 1748
rect 15293 1696 15299 1748
rect 15351 1696 15357 1748
rect 15601 1696 15607 1748
rect 15659 1696 15665 1748
rect 15909 1696 15915 1748
rect 15967 1696 15973 1748
rect 16217 1696 16223 1748
rect 16275 1696 16281 1748
rect 16525 1696 16531 1748
rect 16583 1696 16589 1748
rect 16833 1696 16839 1748
rect 16891 1696 16897 1748
rect 17141 1696 17147 1748
rect 17199 1696 17205 1748
rect 17449 1696 17455 1748
rect 17507 1696 17513 1748
rect 17757 1696 17763 1748
rect 17815 1696 17821 1748
rect 18065 1696 18071 1748
rect 18123 1696 18129 1748
rect 18373 1696 18379 1748
rect 18431 1696 18437 1748
rect 18681 1696 18687 1748
rect 18739 1696 18745 1748
rect 18989 1696 18995 1748
rect 19047 1696 19053 1748
rect 19297 1696 19303 1748
rect 19355 1696 19361 1748
rect 19605 1696 19611 1748
rect 19663 1696 19669 1748
rect 19913 1696 19919 1748
rect 19971 1696 19977 1748
rect 20221 1696 20227 1748
rect 20279 1696 20285 1748
rect 20529 1696 20535 1748
rect 20587 1696 20593 1748
rect 20837 1696 20843 1748
rect 20895 1696 20901 1748
rect 21145 1696 21151 1748
rect 21203 1696 21209 1748
rect 21453 1696 21459 1748
rect 21511 1696 21517 1748
rect 21761 1696 21767 1748
rect 21819 1696 21825 1748
rect 22069 1696 22075 1748
rect 22127 1696 22133 1748
rect 22377 1696 22383 1748
rect 22435 1696 22441 1748
rect 22685 1696 22691 1748
rect 22743 1696 22749 1748
rect 22993 1696 22999 1748
rect 23051 1696 23057 1748
rect 23301 1696 23307 1748
rect 23359 1696 23365 1748
rect 23609 1696 23615 1748
rect 23667 1696 23673 1748
rect 23917 1696 23923 1748
rect 23975 1696 23981 1748
rect 24225 1696 24231 1748
rect 24283 1696 24289 1748
rect 4820 1581 4826 1633
rect 4878 1581 4884 1633
rect 5228 1581 5234 1633
rect 5286 1581 5292 1633
rect 5636 1581 5642 1633
rect 5694 1581 5700 1633
rect 14509 1426 14515 1478
rect 14567 1426 14573 1478
rect 24345 1426 24351 1478
rect 24403 1426 24409 1478
rect 14509 510 14515 562
rect 14567 510 14573 562
rect 24345 510 24351 562
rect 24403 510 24409 562
rect 14683 43 14735 49
rect 14683 -15 14735 -9
rect 14991 43 15043 49
rect 14991 -15 15043 -9
rect 15299 43 15351 49
rect 15299 -15 15351 -9
rect 15607 43 15659 49
rect 15607 -15 15659 -9
rect 15915 43 15967 49
rect 15915 -15 15967 -9
rect 16223 43 16275 49
rect 16223 -15 16275 -9
rect 16531 43 16583 49
rect 16531 -15 16583 -9
rect 16839 43 16891 49
rect 16839 -15 16891 -9
rect 17147 43 17199 49
rect 17147 -15 17199 -9
rect 17455 43 17507 49
rect 17455 -15 17507 -9
rect 17763 43 17815 49
rect 17763 -15 17815 -9
rect 18071 43 18123 49
rect 18071 -15 18123 -9
rect 18379 43 18431 49
rect 18379 -15 18431 -9
rect 18687 43 18739 49
rect 18687 -15 18739 -9
rect 18995 43 19047 49
rect 18995 -15 19047 -9
rect 19303 43 19355 49
rect 19303 -15 19355 -9
rect 19611 43 19663 49
rect 19611 -15 19663 -9
rect 19919 43 19971 49
rect 19919 -15 19971 -9
rect 20227 43 20279 49
rect 20227 -15 20279 -9
rect 20535 43 20587 49
rect 20535 -15 20587 -9
rect 20843 43 20895 49
rect 20843 -15 20895 -9
rect 21151 43 21203 49
rect 21151 -15 21203 -9
rect 21459 43 21511 49
rect 21459 -15 21511 -9
rect 21767 43 21819 49
rect 21767 -15 21819 -9
rect 22075 43 22127 49
rect 22075 -15 22127 -9
rect 22383 43 22435 49
rect 22383 -15 22435 -9
rect 22691 43 22743 49
rect 22691 -15 22743 -9
rect 22999 43 23051 49
rect 22999 -15 23051 -9
rect 23307 43 23359 49
rect 23307 -15 23359 -9
rect 23615 43 23667 49
rect 23615 -15 23667 -9
rect 23923 43 23975 49
rect 23923 -15 23975 -9
rect 24231 43 24283 49
rect 24231 -15 24283 -9
<< via1 >>
rect 8207 12170 8259 12222
rect 60255 12170 60307 12222
rect 2737 11959 2789 12011
rect 3985 11959 4037 12011
rect 5583 11959 5635 12011
rect 7231 11959 7283 12011
rect 8112 11839 8164 11891
rect 8112 11635 8164 11687
rect 8112 11431 8164 11483
rect 8112 11227 8164 11279
rect 8112 11023 8164 11075
rect 8112 10819 8164 10871
rect 8112 10615 8164 10667
rect 8112 10411 8164 10463
rect 2737 10243 2789 10295
rect 3985 10243 4037 10295
rect 5583 10243 5635 10295
rect 7231 10243 7283 10295
rect 115 9820 167 9872
rect 1339 9395 1391 9447
rect 1409 9147 1461 9199
rect 115 8868 167 8920
rect 1339 8443 1391 8495
rect 115 7831 167 7883
rect 1339 7209 1391 7261
rect 328 7093 380 7102
rect 328 7059 337 7093
rect 337 7059 371 7093
rect 371 7059 380 7093
rect 328 7050 380 7059
rect 736 7093 788 7102
rect 736 7059 745 7093
rect 745 7059 779 7093
rect 779 7059 788 7093
rect 736 7050 788 7059
rect 1144 7093 1196 7102
rect 1144 7059 1153 7093
rect 1153 7059 1187 7093
rect 1187 7059 1196 7093
rect 1144 7050 1196 7059
rect 8154 9766 8206 9818
rect 8101 8728 8153 8780
rect 60325 8728 60377 8780
rect 8101 7812 8153 7864
rect 60325 7812 60377 7864
rect 7009 6490 7061 6542
rect 7631 6490 7683 6542
rect 7950 6413 8002 6422
rect 7950 6379 7959 6413
rect 7959 6379 7993 6413
rect 7993 6379 8002 6413
rect 7950 6370 8002 6379
rect 7950 6209 8002 6218
rect 7950 6175 7959 6209
rect 7959 6175 7993 6209
rect 7993 6175 8002 6209
rect 7950 6166 8002 6175
rect 7950 6005 8002 6014
rect 7950 5971 7959 6005
rect 7959 5971 7993 6005
rect 7993 5971 8002 6005
rect 7950 5962 8002 5971
rect 7950 5801 8002 5810
rect 7950 5767 7959 5801
rect 7959 5767 7993 5801
rect 7993 5767 8002 5801
rect 7950 5758 8002 5767
rect 7950 5597 8002 5606
rect 7950 5563 7959 5597
rect 7959 5563 7993 5597
rect 7993 5563 8002 5597
rect 7950 5554 8002 5563
rect 7950 5393 8002 5402
rect 7950 5359 7959 5393
rect 7959 5359 7993 5393
rect 7993 5359 8002 5393
rect 7950 5350 8002 5359
rect 7950 5189 8002 5198
rect 7950 5155 7959 5189
rect 7959 5155 7993 5189
rect 7993 5155 8002 5189
rect 7950 5146 8002 5155
rect 7950 4985 8002 4994
rect 7950 4951 7959 4985
rect 7959 4951 7993 4985
rect 7993 4951 8002 4985
rect 7950 4942 8002 4951
rect 7009 4774 7061 4826
rect 7631 4774 7683 4826
rect 8221 4724 8273 4776
rect 9853 4724 9905 4776
rect 11485 4724 11537 4776
rect 13117 4724 13169 4776
rect 14749 4724 14801 4776
rect 16381 4724 16433 4776
rect 18013 4724 18065 4776
rect 19645 4724 19697 4776
rect 21277 4724 21329 4776
rect 22909 4724 22961 4776
rect 24541 4724 24593 4776
rect 26173 4724 26225 4776
rect 27805 4724 27857 4776
rect 29437 4724 29489 4776
rect 31069 4724 31121 4776
rect 32701 4724 32753 4776
rect 34333 4724 34385 4776
rect 35965 4724 36017 4776
rect 37597 4724 37649 4776
rect 39229 4724 39281 4776
rect 40861 4724 40913 4776
rect 42493 4724 42545 4776
rect 44125 4724 44177 4776
rect 45757 4724 45809 4776
rect 47389 4724 47441 4776
rect 49021 4724 49073 4776
rect 50653 4724 50705 4776
rect 52285 4724 52337 4776
rect 53917 4724 53969 4776
rect 55549 4724 55601 4776
rect 57181 4724 57233 4776
rect 58813 4724 58865 4776
rect 4613 4351 4665 4403
rect 24231 4061 24283 4113
rect 58813 4061 58865 4113
rect 5837 3926 5889 3978
rect 23923 3959 23975 4011
rect 57181 3959 57233 4011
rect 23615 3857 23667 3909
rect 55549 3857 55601 3909
rect 17455 3755 17507 3807
rect 22909 3755 22961 3807
rect 23307 3755 23359 3807
rect 53917 3755 53969 3807
rect 22999 3653 23051 3705
rect 52285 3653 52337 3705
rect 22691 3551 22743 3603
rect 50653 3551 50705 3603
rect 4613 3399 4665 3451
rect 22383 3449 22435 3501
rect 49021 3449 49073 3501
rect 22075 3347 22127 3399
rect 47389 3347 47441 3399
rect 21767 3245 21819 3297
rect 45757 3245 45809 3297
rect 21151 3143 21203 3195
rect 42493 3143 42545 3195
rect 20843 3041 20895 3093
rect 40861 3041 40913 3093
rect -1395 2957 -1343 2966
rect -1395 2923 -1386 2957
rect -1386 2923 -1352 2957
rect -1352 2923 -1343 2957
rect -1395 2914 -1343 2923
rect 42 2995 94 3004
rect 42 2961 51 2995
rect 51 2961 85 2995
rect 85 2961 94 2995
rect 42 2952 94 2961
rect 5837 2974 5889 3026
rect 20535 2939 20587 2991
rect 39229 2939 39281 2991
rect 20227 2837 20279 2889
rect 37597 2837 37649 2889
rect 16839 2735 16891 2787
rect 19645 2735 19697 2787
rect 19919 2735 19971 2787
rect 35965 2735 36017 2787
rect 19611 2633 19663 2685
rect 34333 2633 34385 2685
rect 19303 2531 19355 2583
rect 32701 2531 32753 2583
rect 18995 2429 19047 2481
rect 31069 2429 31121 2481
rect 4613 2362 4665 2414
rect 14749 2327 14801 2379
rect 15915 2327 15967 2379
rect 18687 2327 18739 2379
rect 29437 2327 29489 2379
rect 13117 2225 13169 2277
rect 15607 2225 15659 2277
rect 16531 2225 16583 2277
rect 18013 2225 18065 2277
rect 18379 2225 18431 2277
rect 27805 2225 27857 2277
rect 11485 2123 11537 2175
rect 15299 2123 15351 2175
rect 18071 2123 18123 2175
rect 26173 2123 26225 2175
rect 9853 2021 9905 2073
rect 14991 2021 15043 2073
rect 17763 2021 17815 2073
rect 24541 2021 24593 2073
rect 449 1950 501 1959
rect 449 1916 458 1950
rect 458 1916 492 1950
rect 492 1916 501 1950
rect 449 1907 501 1916
rect 8221 1919 8273 1971
rect 14683 1919 14735 1971
rect 16223 1919 16275 1971
rect 16381 1919 16433 1971
rect 17147 1919 17199 1971
rect 21277 1919 21329 1971
rect 21459 1919 21511 1971
rect 44125 1919 44177 1971
rect 5837 1740 5889 1792
rect 14683 1739 14735 1748
rect 14683 1705 14692 1739
rect 14692 1705 14726 1739
rect 14726 1705 14735 1739
rect 14683 1696 14735 1705
rect 14991 1739 15043 1748
rect 14991 1705 15000 1739
rect 15000 1705 15034 1739
rect 15034 1705 15043 1739
rect 14991 1696 15043 1705
rect 15299 1739 15351 1748
rect 15299 1705 15308 1739
rect 15308 1705 15342 1739
rect 15342 1705 15351 1739
rect 15299 1696 15351 1705
rect 15607 1739 15659 1748
rect 15607 1705 15616 1739
rect 15616 1705 15650 1739
rect 15650 1705 15659 1739
rect 15607 1696 15659 1705
rect 15915 1739 15967 1748
rect 15915 1705 15924 1739
rect 15924 1705 15958 1739
rect 15958 1705 15967 1739
rect 15915 1696 15967 1705
rect 16223 1739 16275 1748
rect 16223 1705 16232 1739
rect 16232 1705 16266 1739
rect 16266 1705 16275 1739
rect 16223 1696 16275 1705
rect 16531 1739 16583 1748
rect 16531 1705 16540 1739
rect 16540 1705 16574 1739
rect 16574 1705 16583 1739
rect 16531 1696 16583 1705
rect 16839 1739 16891 1748
rect 16839 1705 16848 1739
rect 16848 1705 16882 1739
rect 16882 1705 16891 1739
rect 16839 1696 16891 1705
rect 17147 1739 17199 1748
rect 17147 1705 17156 1739
rect 17156 1705 17190 1739
rect 17190 1705 17199 1739
rect 17147 1696 17199 1705
rect 17455 1739 17507 1748
rect 17455 1705 17464 1739
rect 17464 1705 17498 1739
rect 17498 1705 17507 1739
rect 17455 1696 17507 1705
rect 17763 1739 17815 1748
rect 17763 1705 17772 1739
rect 17772 1705 17806 1739
rect 17806 1705 17815 1739
rect 17763 1696 17815 1705
rect 18071 1739 18123 1748
rect 18071 1705 18080 1739
rect 18080 1705 18114 1739
rect 18114 1705 18123 1739
rect 18071 1696 18123 1705
rect 18379 1739 18431 1748
rect 18379 1705 18388 1739
rect 18388 1705 18422 1739
rect 18422 1705 18431 1739
rect 18379 1696 18431 1705
rect 18687 1739 18739 1748
rect 18687 1705 18696 1739
rect 18696 1705 18730 1739
rect 18730 1705 18739 1739
rect 18687 1696 18739 1705
rect 18995 1739 19047 1748
rect 18995 1705 19004 1739
rect 19004 1705 19038 1739
rect 19038 1705 19047 1739
rect 18995 1696 19047 1705
rect 19303 1739 19355 1748
rect 19303 1705 19312 1739
rect 19312 1705 19346 1739
rect 19346 1705 19355 1739
rect 19303 1696 19355 1705
rect 19611 1739 19663 1748
rect 19611 1705 19620 1739
rect 19620 1705 19654 1739
rect 19654 1705 19663 1739
rect 19611 1696 19663 1705
rect 19919 1739 19971 1748
rect 19919 1705 19928 1739
rect 19928 1705 19962 1739
rect 19962 1705 19971 1739
rect 19919 1696 19971 1705
rect 20227 1739 20279 1748
rect 20227 1705 20236 1739
rect 20236 1705 20270 1739
rect 20270 1705 20279 1739
rect 20227 1696 20279 1705
rect 20535 1739 20587 1748
rect 20535 1705 20544 1739
rect 20544 1705 20578 1739
rect 20578 1705 20587 1739
rect 20535 1696 20587 1705
rect 20843 1739 20895 1748
rect 20843 1705 20852 1739
rect 20852 1705 20886 1739
rect 20886 1705 20895 1739
rect 20843 1696 20895 1705
rect 21151 1739 21203 1748
rect 21151 1705 21160 1739
rect 21160 1705 21194 1739
rect 21194 1705 21203 1739
rect 21151 1696 21203 1705
rect 21459 1739 21511 1748
rect 21459 1705 21468 1739
rect 21468 1705 21502 1739
rect 21502 1705 21511 1739
rect 21459 1696 21511 1705
rect 21767 1739 21819 1748
rect 21767 1705 21776 1739
rect 21776 1705 21810 1739
rect 21810 1705 21819 1739
rect 21767 1696 21819 1705
rect 22075 1739 22127 1748
rect 22075 1705 22084 1739
rect 22084 1705 22118 1739
rect 22118 1705 22127 1739
rect 22075 1696 22127 1705
rect 22383 1739 22435 1748
rect 22383 1705 22392 1739
rect 22392 1705 22426 1739
rect 22426 1705 22435 1739
rect 22383 1696 22435 1705
rect 22691 1739 22743 1748
rect 22691 1705 22700 1739
rect 22700 1705 22734 1739
rect 22734 1705 22743 1739
rect 22691 1696 22743 1705
rect 22999 1739 23051 1748
rect 22999 1705 23008 1739
rect 23008 1705 23042 1739
rect 23042 1705 23051 1739
rect 22999 1696 23051 1705
rect 23307 1739 23359 1748
rect 23307 1705 23316 1739
rect 23316 1705 23350 1739
rect 23350 1705 23359 1739
rect 23307 1696 23359 1705
rect 23615 1739 23667 1748
rect 23615 1705 23624 1739
rect 23624 1705 23658 1739
rect 23658 1705 23667 1739
rect 23615 1696 23667 1705
rect 23923 1739 23975 1748
rect 23923 1705 23932 1739
rect 23932 1705 23966 1739
rect 23966 1705 23975 1739
rect 23923 1696 23975 1705
rect 24231 1739 24283 1748
rect 24231 1705 24240 1739
rect 24240 1705 24274 1739
rect 24274 1705 24283 1739
rect 24231 1696 24283 1705
rect 4826 1624 4878 1633
rect 4826 1590 4835 1624
rect 4835 1590 4869 1624
rect 4869 1590 4878 1624
rect 4826 1581 4878 1590
rect 5234 1624 5286 1633
rect 5234 1590 5243 1624
rect 5243 1590 5277 1624
rect 5277 1590 5286 1624
rect 5234 1581 5286 1590
rect 5642 1624 5694 1633
rect 5642 1590 5651 1624
rect 5651 1590 5685 1624
rect 5685 1590 5694 1624
rect 5642 1581 5694 1590
rect 14515 1426 14567 1478
rect 24351 1426 24403 1478
rect 14515 510 14567 562
rect 24351 510 24403 562
rect 14683 34 14735 43
rect 14683 0 14692 34
rect 14692 0 14726 34
rect 14726 0 14735 34
rect 14683 -9 14735 0
rect 14991 34 15043 43
rect 14991 0 15000 34
rect 15000 0 15034 34
rect 15034 0 15043 34
rect 14991 -9 15043 0
rect 15299 34 15351 43
rect 15299 0 15308 34
rect 15308 0 15342 34
rect 15342 0 15351 34
rect 15299 -9 15351 0
rect 15607 34 15659 43
rect 15607 0 15616 34
rect 15616 0 15650 34
rect 15650 0 15659 34
rect 15607 -9 15659 0
rect 15915 34 15967 43
rect 15915 0 15924 34
rect 15924 0 15958 34
rect 15958 0 15967 34
rect 15915 -9 15967 0
rect 16223 34 16275 43
rect 16223 0 16232 34
rect 16232 0 16266 34
rect 16266 0 16275 34
rect 16223 -9 16275 0
rect 16531 34 16583 43
rect 16531 0 16540 34
rect 16540 0 16574 34
rect 16574 0 16583 34
rect 16531 -9 16583 0
rect 16839 34 16891 43
rect 16839 0 16848 34
rect 16848 0 16882 34
rect 16882 0 16891 34
rect 16839 -9 16891 0
rect 17147 34 17199 43
rect 17147 0 17156 34
rect 17156 0 17190 34
rect 17190 0 17199 34
rect 17147 -9 17199 0
rect 17455 34 17507 43
rect 17455 0 17464 34
rect 17464 0 17498 34
rect 17498 0 17507 34
rect 17455 -9 17507 0
rect 17763 34 17815 43
rect 17763 0 17772 34
rect 17772 0 17806 34
rect 17806 0 17815 34
rect 17763 -9 17815 0
rect 18071 34 18123 43
rect 18071 0 18080 34
rect 18080 0 18114 34
rect 18114 0 18123 34
rect 18071 -9 18123 0
rect 18379 34 18431 43
rect 18379 0 18388 34
rect 18388 0 18422 34
rect 18422 0 18431 34
rect 18379 -9 18431 0
rect 18687 34 18739 43
rect 18687 0 18696 34
rect 18696 0 18730 34
rect 18730 0 18739 34
rect 18687 -9 18739 0
rect 18995 34 19047 43
rect 18995 0 19004 34
rect 19004 0 19038 34
rect 19038 0 19047 34
rect 18995 -9 19047 0
rect 19303 34 19355 43
rect 19303 0 19312 34
rect 19312 0 19346 34
rect 19346 0 19355 34
rect 19303 -9 19355 0
rect 19611 34 19663 43
rect 19611 0 19620 34
rect 19620 0 19654 34
rect 19654 0 19663 34
rect 19611 -9 19663 0
rect 19919 34 19971 43
rect 19919 0 19928 34
rect 19928 0 19962 34
rect 19962 0 19971 34
rect 19919 -9 19971 0
rect 20227 34 20279 43
rect 20227 0 20236 34
rect 20236 0 20270 34
rect 20270 0 20279 34
rect 20227 -9 20279 0
rect 20535 34 20587 43
rect 20535 0 20544 34
rect 20544 0 20578 34
rect 20578 0 20587 34
rect 20535 -9 20587 0
rect 20843 34 20895 43
rect 20843 0 20852 34
rect 20852 0 20886 34
rect 20886 0 20895 34
rect 20843 -9 20895 0
rect 21151 34 21203 43
rect 21151 0 21160 34
rect 21160 0 21194 34
rect 21194 0 21203 34
rect 21151 -9 21203 0
rect 21459 34 21511 43
rect 21459 0 21468 34
rect 21468 0 21502 34
rect 21502 0 21511 34
rect 21459 -9 21511 0
rect 21767 34 21819 43
rect 21767 0 21776 34
rect 21776 0 21810 34
rect 21810 0 21819 34
rect 21767 -9 21819 0
rect 22075 34 22127 43
rect 22075 0 22084 34
rect 22084 0 22118 34
rect 22118 0 22127 34
rect 22075 -9 22127 0
rect 22383 34 22435 43
rect 22383 0 22392 34
rect 22392 0 22426 34
rect 22426 0 22435 34
rect 22383 -9 22435 0
rect 22691 34 22743 43
rect 22691 0 22700 34
rect 22700 0 22734 34
rect 22734 0 22743 34
rect 22691 -9 22743 0
rect 22999 34 23051 43
rect 22999 0 23008 34
rect 23008 0 23042 34
rect 23042 0 23051 34
rect 22999 -9 23051 0
rect 23307 34 23359 43
rect 23307 0 23316 34
rect 23316 0 23350 34
rect 23350 0 23359 34
rect 23307 -9 23359 0
rect 23615 34 23667 43
rect 23615 0 23624 34
rect 23624 0 23658 34
rect 23658 0 23667 34
rect 23615 -9 23667 0
rect 23923 34 23975 43
rect 23923 0 23932 34
rect 23932 0 23966 34
rect 23966 0 23975 34
rect 23923 -9 23975 0
rect 24231 34 24283 43
rect 24231 0 24240 34
rect 24240 0 24274 34
rect 24274 0 24283 34
rect 24231 -9 24283 0
<< metal2 >>
rect 8205 12224 8261 12233
rect 8205 12159 8261 12168
rect 60253 12224 60309 12233
rect 60253 12159 60309 12168
rect 2735 12013 2791 12022
rect 2735 11948 2791 11957
rect 3983 12013 4039 12022
rect 3983 11948 4039 11957
rect 5581 12013 5637 12022
rect 5581 11948 5637 11957
rect 7229 12013 7285 12022
rect 7229 11948 7285 11957
rect 8112 11891 8164 11897
rect 8106 11844 8112 11887
rect 8164 11844 8170 11887
rect 8112 11833 8164 11839
rect 8112 11687 8164 11693
rect 8106 11640 8112 11683
rect 8164 11640 8170 11683
rect 8112 11629 8164 11635
rect 8112 11483 8164 11489
rect 8106 11436 8112 11479
rect 8164 11436 8170 11479
rect 8112 11425 8164 11431
rect 8112 11279 8164 11285
rect 8106 11232 8112 11275
rect 8164 11232 8170 11275
rect 8112 11221 8164 11227
rect 8112 11075 8164 11081
rect 8106 11028 8112 11071
rect 8164 11028 8170 11071
rect 8112 11017 8164 11023
rect 8112 10871 8164 10877
rect 8106 10824 8112 10867
rect 8164 10824 8170 10867
rect 8112 10813 8164 10819
rect 8112 10667 8164 10673
rect 8106 10620 8112 10663
rect 8164 10620 8170 10663
rect 8112 10609 8164 10615
rect 8112 10463 8164 10469
rect 8106 10416 8112 10459
rect 8164 10416 8170 10459
rect 8112 10405 8164 10411
rect 34338 10311 34394 10320
rect 2735 10297 2791 10306
rect 1421 10252 1905 10280
rect 113 9874 169 9883
rect 113 9809 169 9818
rect 1337 9449 1393 9458
rect 1337 9384 1393 9393
rect 1421 9205 1449 10252
rect 2245 10245 2301 10254
rect 2735 10232 2791 10241
rect 3983 10297 4039 10306
rect 3983 10232 4039 10241
rect 5581 10297 5637 10306
rect 5581 10232 5637 10241
rect 7229 10297 7285 10306
rect 34338 10246 34394 10255
rect 7229 10232 7285 10241
rect 2245 10180 2301 10189
rect 8154 9818 8206 9824
rect 8154 9760 8206 9766
rect 8103 9438 8159 9447
rect 8103 9373 8159 9382
rect 1409 9199 1461 9205
rect 1461 9159 4352 9187
rect 1409 9141 1461 9147
rect 113 8922 169 8931
rect 113 8857 169 8866
rect 1337 8497 1393 8506
rect 1337 8432 1393 8441
rect 113 7885 169 7894
rect 113 7820 169 7829
rect 1337 7263 1393 7272
rect 1337 7198 1393 7207
rect 326 7104 382 7113
rect 326 7039 382 7048
rect 734 7104 790 7113
rect 734 7039 790 7048
rect 1142 7104 1198 7113
rect 1142 7039 1198 7048
rect 42 3004 94 3010
rect -1397 2968 -1341 2977
rect 4324 2992 4352 9159
rect 8099 8782 8155 8791
rect 8099 8717 8155 8726
rect 60323 8782 60379 8791
rect 60323 8717 60379 8726
rect 8099 7866 8155 7875
rect 8099 7801 8155 7810
rect 60323 7866 60379 7875
rect 60323 7801 60379 7810
rect 34270 7364 34326 7373
rect 34270 7299 34326 7308
rect 7007 6544 7063 6553
rect 7007 6479 7063 6488
rect 7629 6544 7685 6553
rect 7629 6479 7685 6488
rect 7950 6422 8002 6428
rect 8002 6382 60377 6410
rect 7950 6364 8002 6370
rect 7950 6218 8002 6224
rect 8002 6178 60377 6206
rect 7950 6160 8002 6166
rect 7950 6014 8002 6020
rect 8002 5974 60377 6002
rect 7950 5956 8002 5962
rect 7950 5810 8002 5816
rect 8002 5770 60377 5798
rect 7950 5752 8002 5758
rect 7950 5606 8002 5612
rect 8002 5566 60377 5594
rect 7950 5548 8002 5554
rect 7950 5402 8002 5408
rect 8002 5362 60377 5390
rect 7950 5344 8002 5350
rect 7950 5198 8002 5204
rect 8002 5158 60377 5186
rect 7950 5140 8002 5146
rect 7950 4994 8002 5000
rect 8002 4954 60377 4982
rect 7950 4936 8002 4942
rect 7007 4828 7063 4837
rect 6743 4776 6799 4785
rect 7007 4763 7063 4772
rect 7629 4828 7685 4837
rect 7629 4763 7685 4772
rect 8221 4776 8273 4782
rect 6743 4711 6799 4720
rect 8221 4718 8273 4724
rect 9853 4776 9905 4782
rect 9853 4718 9905 4724
rect 11485 4776 11537 4782
rect 11485 4718 11537 4724
rect 13117 4776 13169 4782
rect 13117 4718 13169 4724
rect 14749 4776 14801 4782
rect 14749 4718 14801 4724
rect 16381 4776 16433 4782
rect 16381 4718 16433 4724
rect 18013 4776 18065 4782
rect 18013 4718 18065 4724
rect 19645 4776 19697 4782
rect 19645 4718 19697 4724
rect 21277 4776 21329 4782
rect 21277 4718 21329 4724
rect 22909 4776 22961 4782
rect 22909 4718 22961 4724
rect 24541 4776 24593 4782
rect 24541 4718 24593 4724
rect 26173 4776 26225 4782
rect 26173 4718 26225 4724
rect 27805 4776 27857 4782
rect 27805 4718 27857 4724
rect 29437 4776 29489 4782
rect 29437 4718 29489 4724
rect 31069 4776 31121 4782
rect 31069 4718 31121 4724
rect 32701 4776 32753 4782
rect 32701 4718 32753 4724
rect 34333 4776 34385 4782
rect 34333 4718 34385 4724
rect 35965 4776 36017 4782
rect 35965 4718 36017 4724
rect 37597 4776 37649 4782
rect 37597 4718 37649 4724
rect 39229 4776 39281 4782
rect 39229 4718 39281 4724
rect 40861 4776 40913 4782
rect 40861 4718 40913 4724
rect 42493 4776 42545 4782
rect 42493 4718 42545 4724
rect 44125 4776 44177 4782
rect 44125 4718 44177 4724
rect 45757 4776 45809 4782
rect 45757 4718 45809 4724
rect 47389 4776 47441 4782
rect 47389 4718 47441 4724
rect 49021 4776 49073 4782
rect 49021 4718 49073 4724
rect 50653 4776 50705 4782
rect 50653 4718 50705 4724
rect 52285 4776 52337 4782
rect 52285 4718 52337 4724
rect 53917 4776 53969 4782
rect 53917 4718 53969 4724
rect 55549 4776 55601 4782
rect 55549 4718 55601 4724
rect 57181 4776 57233 4782
rect 57181 4718 57233 4724
rect 58813 4776 58865 4782
rect 58813 4718 58865 4724
rect 4611 4405 4667 4414
rect 4611 4340 4667 4349
rect 5835 3980 5891 3989
rect 5835 3915 5891 3924
rect 4611 3453 4667 3462
rect 4611 3388 4667 3397
rect 94 2964 4352 2992
rect 5835 3028 5891 3037
rect 5835 2963 5891 2972
rect 42 2946 94 2952
rect -1397 2903 -1341 2912
rect 4611 2416 4667 2425
rect 4611 2351 4667 2360
rect 8233 1977 8261 4718
rect 9865 2079 9893 4718
rect 11497 2181 11525 4718
rect 13129 2283 13157 4718
rect 14761 2385 14789 4718
rect 14749 2379 14801 2385
rect 14749 2321 14801 2327
rect 15915 2379 15967 2385
rect 15915 2321 15967 2327
rect 13117 2277 13169 2283
rect 13117 2219 13169 2225
rect 15607 2277 15659 2283
rect 15607 2219 15659 2225
rect 11485 2175 11537 2181
rect 11485 2117 11537 2123
rect 15299 2175 15351 2181
rect 15299 2117 15351 2123
rect 9853 2073 9905 2079
rect 9853 2015 9905 2021
rect 14991 2073 15043 2079
rect 14991 2015 15043 2021
rect 8221 1971 8273 1977
rect 447 1961 503 1970
rect 8221 1913 8273 1919
rect 14683 1971 14735 1977
rect 14683 1913 14735 1919
rect 447 1896 503 1905
rect 5835 1794 5891 1803
rect 14695 1754 14723 1913
rect 15003 1754 15031 2015
rect 15311 1754 15339 2117
rect 15619 1754 15647 2219
rect 15927 1754 15955 2321
rect 16393 1977 16421 4718
rect 17455 3807 17507 3813
rect 17455 3749 17507 3755
rect 16839 2787 16891 2793
rect 16839 2729 16891 2735
rect 16531 2277 16583 2283
rect 16531 2219 16583 2225
rect 16223 1971 16275 1977
rect 16223 1913 16275 1919
rect 16381 1971 16433 1977
rect 16381 1913 16433 1919
rect 16235 1754 16263 1913
rect 16543 1754 16571 2219
rect 16851 1754 16879 2729
rect 17147 1971 17199 1977
rect 17147 1913 17199 1919
rect 17159 1754 17187 1913
rect 17467 1754 17495 3749
rect 18025 2283 18053 4718
rect 19657 2793 19685 4718
rect 21151 3195 21203 3201
rect 21151 3137 21203 3143
rect 20843 3093 20895 3099
rect 20843 3035 20895 3041
rect 20535 2991 20587 2997
rect 20535 2933 20587 2939
rect 20227 2889 20279 2895
rect 20227 2831 20279 2837
rect 19645 2787 19697 2793
rect 19645 2729 19697 2735
rect 19919 2787 19971 2793
rect 19919 2729 19971 2735
rect 19611 2685 19663 2691
rect 19611 2627 19663 2633
rect 19303 2583 19355 2589
rect 19303 2525 19355 2531
rect 18995 2481 19047 2487
rect 18995 2423 19047 2429
rect 18687 2379 18739 2385
rect 18687 2321 18739 2327
rect 18013 2277 18065 2283
rect 18013 2219 18065 2225
rect 18379 2277 18431 2283
rect 18379 2219 18431 2225
rect 18071 2175 18123 2181
rect 18071 2117 18123 2123
rect 17763 2073 17815 2079
rect 17763 2015 17815 2021
rect 17775 1754 17803 2015
rect 18083 1754 18111 2117
rect 18391 1754 18419 2219
rect 18699 1754 18727 2321
rect 19007 1754 19035 2423
rect 19315 1754 19343 2525
rect 19623 1754 19651 2627
rect 19931 1754 19959 2729
rect 20239 1754 20267 2831
rect 20547 1754 20575 2933
rect 20855 1754 20883 3035
rect 21163 1754 21191 3137
rect 21289 1977 21317 4718
rect 22921 3813 22949 4718
rect 24231 4113 24283 4119
rect 24231 4055 24283 4061
rect 23923 4011 23975 4017
rect 23923 3953 23975 3959
rect 23615 3909 23667 3915
rect 23615 3851 23667 3857
rect 22909 3807 22961 3813
rect 22909 3749 22961 3755
rect 23307 3807 23359 3813
rect 23307 3749 23359 3755
rect 22999 3705 23051 3711
rect 22999 3647 23051 3653
rect 22691 3603 22743 3609
rect 22691 3545 22743 3551
rect 22383 3501 22435 3507
rect 22383 3443 22435 3449
rect 22075 3399 22127 3405
rect 22075 3341 22127 3347
rect 21767 3297 21819 3303
rect 21767 3239 21819 3245
rect 21277 1971 21329 1977
rect 21277 1913 21329 1919
rect 21459 1971 21511 1977
rect 21459 1913 21511 1919
rect 21471 1754 21499 1913
rect 21779 1754 21807 3239
rect 22087 1754 22115 3341
rect 22395 1754 22423 3443
rect 22703 1754 22731 3545
rect 23011 1754 23039 3647
rect 23319 1754 23347 3749
rect 23627 1754 23655 3851
rect 23935 1754 23963 3953
rect 24243 1754 24271 4055
rect 24553 2079 24581 4718
rect 26185 2181 26213 4718
rect 27817 2283 27845 4718
rect 29449 2385 29477 4718
rect 31081 2487 31109 4718
rect 32713 2589 32741 4718
rect 34345 2691 34373 4718
rect 35977 2793 36005 4718
rect 37609 2895 37637 4718
rect 39241 2997 39269 4718
rect 40873 3099 40901 4718
rect 42505 3201 42533 4718
rect 42493 3195 42545 3201
rect 42493 3137 42545 3143
rect 40861 3093 40913 3099
rect 40861 3035 40913 3041
rect 39229 2991 39281 2997
rect 39229 2933 39281 2939
rect 37597 2889 37649 2895
rect 37597 2831 37649 2837
rect 35965 2787 36017 2793
rect 35965 2729 36017 2735
rect 34333 2685 34385 2691
rect 34333 2627 34385 2633
rect 32701 2583 32753 2589
rect 32701 2525 32753 2531
rect 31069 2481 31121 2487
rect 31069 2423 31121 2429
rect 29437 2379 29489 2385
rect 29437 2321 29489 2327
rect 27805 2277 27857 2283
rect 27805 2219 27857 2225
rect 26173 2175 26225 2181
rect 26173 2117 26225 2123
rect 24541 2073 24593 2079
rect 24541 2015 24593 2021
rect 44137 1977 44165 4718
rect 45769 3303 45797 4718
rect 47401 3405 47429 4718
rect 49033 3507 49061 4718
rect 50665 3609 50693 4718
rect 52297 3711 52325 4718
rect 53929 3813 53957 4718
rect 55561 3915 55589 4718
rect 57193 4017 57221 4718
rect 58825 4119 58853 4718
rect 58813 4113 58865 4119
rect 58813 4055 58865 4061
rect 57181 4011 57233 4017
rect 57181 3953 57233 3959
rect 55549 3909 55601 3915
rect 55549 3851 55601 3857
rect 53917 3807 53969 3813
rect 53917 3749 53969 3755
rect 52285 3705 52337 3711
rect 52285 3647 52337 3653
rect 50653 3603 50705 3609
rect 50653 3545 50705 3551
rect 49021 3501 49073 3507
rect 49021 3443 49073 3449
rect 47389 3399 47441 3405
rect 47389 3341 47441 3347
rect 45757 3297 45809 3303
rect 45757 3239 45809 3245
rect 44125 1971 44177 1977
rect 44125 1913 44177 1919
rect 5835 1729 5891 1738
rect 14683 1748 14735 1754
rect 14683 1690 14735 1696
rect 14991 1748 15043 1754
rect 14991 1690 15043 1696
rect 15299 1748 15351 1754
rect 15299 1690 15351 1696
rect 15607 1748 15659 1754
rect 15607 1690 15659 1696
rect 15915 1748 15967 1754
rect 15915 1690 15967 1696
rect 16223 1748 16275 1754
rect 16223 1690 16275 1696
rect 16531 1748 16583 1754
rect 16531 1690 16583 1696
rect 16839 1748 16891 1754
rect 16839 1690 16891 1696
rect 17147 1748 17199 1754
rect 17147 1690 17199 1696
rect 17455 1748 17507 1754
rect 17455 1690 17507 1696
rect 17763 1748 17815 1754
rect 17763 1690 17815 1696
rect 18071 1748 18123 1754
rect 18071 1690 18123 1696
rect 18379 1748 18431 1754
rect 18379 1690 18431 1696
rect 18687 1748 18739 1754
rect 18687 1690 18739 1696
rect 18995 1748 19047 1754
rect 18995 1690 19047 1696
rect 19303 1748 19355 1754
rect 19303 1690 19355 1696
rect 19611 1748 19663 1754
rect 19611 1690 19663 1696
rect 19919 1748 19971 1754
rect 19919 1690 19971 1696
rect 20227 1748 20279 1754
rect 20227 1690 20279 1696
rect 20535 1748 20587 1754
rect 20535 1690 20587 1696
rect 20843 1748 20895 1754
rect 20843 1690 20895 1696
rect 21151 1748 21203 1754
rect 21151 1690 21203 1696
rect 21459 1748 21511 1754
rect 21459 1690 21511 1696
rect 21767 1748 21819 1754
rect 21767 1690 21819 1696
rect 22075 1748 22127 1754
rect 22075 1690 22127 1696
rect 22383 1748 22435 1754
rect 22383 1690 22435 1696
rect 22691 1748 22743 1754
rect 22691 1690 22743 1696
rect 22999 1748 23051 1754
rect 22999 1690 23051 1696
rect 23307 1748 23359 1754
rect 23307 1690 23359 1696
rect 23615 1748 23667 1754
rect 23615 1690 23667 1696
rect 23923 1748 23975 1754
rect 23923 1690 23975 1696
rect 24231 1748 24283 1754
rect 24231 1690 24283 1696
rect 4824 1635 4880 1644
rect 4824 1570 4880 1579
rect 5232 1635 5288 1644
rect 5232 1570 5288 1579
rect 5640 1635 5696 1644
rect 5640 1570 5696 1579
rect 14513 1480 14569 1489
rect 14513 1415 14569 1424
rect 24349 1480 24405 1489
rect 24349 1415 24405 1424
rect 14513 564 14569 573
rect 14513 499 14569 508
rect 24349 564 24405 573
rect 24349 499 24405 508
rect 14672 -11 14681 45
rect 14737 -11 14746 45
rect 14980 -11 14989 45
rect 15045 -11 15054 45
rect 15288 -11 15297 45
rect 15353 -11 15362 45
rect 15596 -11 15605 45
rect 15661 -11 15670 45
rect 15904 -11 15913 45
rect 15969 -11 15978 45
rect 16212 -11 16221 45
rect 16277 -11 16286 45
rect 16520 -11 16529 45
rect 16585 -11 16594 45
rect 16828 -11 16837 45
rect 16893 -11 16902 45
rect 17136 -11 17145 45
rect 17201 -11 17210 45
rect 17444 -11 17453 45
rect 17509 -11 17518 45
rect 17752 -11 17761 45
rect 17817 -11 17826 45
rect 18060 -11 18069 45
rect 18125 -11 18134 45
rect 18368 -11 18377 45
rect 18433 -11 18442 45
rect 18676 -11 18685 45
rect 18741 -11 18750 45
rect 18984 -11 18993 45
rect 19049 -11 19058 45
rect 19292 -11 19301 45
rect 19357 -11 19366 45
rect 19600 -11 19609 45
rect 19665 -11 19674 45
rect 19908 -11 19917 45
rect 19973 -11 19982 45
rect 20216 -11 20225 45
rect 20281 -11 20290 45
rect 20524 -11 20533 45
rect 20589 -11 20598 45
rect 20832 -11 20841 45
rect 20897 -11 20906 45
rect 21140 -11 21149 45
rect 21205 -11 21214 45
rect 21448 -11 21457 45
rect 21513 -11 21522 45
rect 21756 -11 21765 45
rect 21821 -11 21830 45
rect 22064 -11 22073 45
rect 22129 -11 22138 45
rect 22372 -11 22381 45
rect 22437 -11 22446 45
rect 22680 -11 22689 45
rect 22745 -11 22754 45
rect 22988 -11 22997 45
rect 23053 -11 23062 45
rect 23296 -11 23305 45
rect 23361 -11 23370 45
rect 23604 -11 23613 45
rect 23669 -11 23678 45
rect 23912 -11 23921 45
rect 23977 -11 23986 45
rect 24220 -11 24229 45
rect 24285 -11 24294 45
<< via2 >>
rect 8205 12222 8261 12224
rect 8205 12170 8207 12222
rect 8207 12170 8259 12222
rect 8259 12170 8261 12222
rect 8205 12168 8261 12170
rect 60253 12222 60309 12224
rect 60253 12170 60255 12222
rect 60255 12170 60307 12222
rect 60307 12170 60309 12222
rect 60253 12168 60309 12170
rect 2735 12011 2791 12013
rect 2735 11959 2737 12011
rect 2737 11959 2789 12011
rect 2789 11959 2791 12011
rect 2735 11957 2791 11959
rect 3983 12011 4039 12013
rect 3983 11959 3985 12011
rect 3985 11959 4037 12011
rect 4037 11959 4039 12011
rect 3983 11957 4039 11959
rect 5581 12011 5637 12013
rect 5581 11959 5583 12011
rect 5583 11959 5635 12011
rect 5635 11959 5637 12011
rect 5581 11957 5637 11959
rect 7229 12011 7285 12013
rect 7229 11959 7231 12011
rect 7231 11959 7283 12011
rect 7283 11959 7285 12011
rect 7229 11957 7285 11959
rect 2735 10295 2791 10297
rect 113 9872 169 9874
rect 113 9820 115 9872
rect 115 9820 167 9872
rect 167 9820 169 9872
rect 113 9818 169 9820
rect 1337 9447 1393 9449
rect 1337 9395 1339 9447
rect 1339 9395 1391 9447
rect 1391 9395 1393 9447
rect 1337 9393 1393 9395
rect 2245 10189 2301 10245
rect 2735 10243 2737 10295
rect 2737 10243 2789 10295
rect 2789 10243 2791 10295
rect 2735 10241 2791 10243
rect 3983 10295 4039 10297
rect 3983 10243 3985 10295
rect 3985 10243 4037 10295
rect 4037 10243 4039 10295
rect 3983 10241 4039 10243
rect 5581 10295 5637 10297
rect 5581 10243 5583 10295
rect 5583 10243 5635 10295
rect 5635 10243 5637 10295
rect 5581 10241 5637 10243
rect 7229 10295 7285 10297
rect 7229 10243 7231 10295
rect 7231 10243 7283 10295
rect 7283 10243 7285 10295
rect 34338 10255 34394 10311
rect 7229 10241 7285 10243
rect 8103 9382 8159 9438
rect 113 8920 169 8922
rect 113 8868 115 8920
rect 115 8868 167 8920
rect 167 8868 169 8920
rect 113 8866 169 8868
rect 1337 8495 1393 8497
rect 1337 8443 1339 8495
rect 1339 8443 1391 8495
rect 1391 8443 1393 8495
rect 1337 8441 1393 8443
rect 113 7883 169 7885
rect 113 7831 115 7883
rect 115 7831 167 7883
rect 167 7831 169 7883
rect 113 7829 169 7831
rect 1337 7261 1393 7263
rect 1337 7209 1339 7261
rect 1339 7209 1391 7261
rect 1391 7209 1393 7261
rect 1337 7207 1393 7209
rect 326 7102 382 7104
rect 326 7050 328 7102
rect 328 7050 380 7102
rect 380 7050 382 7102
rect 326 7048 382 7050
rect 734 7102 790 7104
rect 734 7050 736 7102
rect 736 7050 788 7102
rect 788 7050 790 7102
rect 734 7048 790 7050
rect 1142 7102 1198 7104
rect 1142 7050 1144 7102
rect 1144 7050 1196 7102
rect 1196 7050 1198 7102
rect 1142 7048 1198 7050
rect -1397 2966 -1341 2968
rect -1397 2914 -1395 2966
rect -1395 2914 -1343 2966
rect -1343 2914 -1341 2966
rect 8099 8780 8155 8782
rect 8099 8728 8101 8780
rect 8101 8728 8153 8780
rect 8153 8728 8155 8780
rect 8099 8726 8155 8728
rect 60323 8780 60379 8782
rect 60323 8728 60325 8780
rect 60325 8728 60377 8780
rect 60377 8728 60379 8780
rect 60323 8726 60379 8728
rect 8099 7864 8155 7866
rect 8099 7812 8101 7864
rect 8101 7812 8153 7864
rect 8153 7812 8155 7864
rect 8099 7810 8155 7812
rect 60323 7864 60379 7866
rect 60323 7812 60325 7864
rect 60325 7812 60377 7864
rect 60377 7812 60379 7864
rect 60323 7810 60379 7812
rect 34270 7308 34326 7364
rect 7007 6542 7063 6544
rect 7007 6490 7009 6542
rect 7009 6490 7061 6542
rect 7061 6490 7063 6542
rect 7007 6488 7063 6490
rect 7629 6542 7685 6544
rect 7629 6490 7631 6542
rect 7631 6490 7683 6542
rect 7683 6490 7685 6542
rect 7629 6488 7685 6490
rect 7007 4826 7063 4828
rect 6743 4720 6799 4776
rect 7007 4774 7009 4826
rect 7009 4774 7061 4826
rect 7061 4774 7063 4826
rect 7007 4772 7063 4774
rect 7629 4826 7685 4828
rect 7629 4774 7631 4826
rect 7631 4774 7683 4826
rect 7683 4774 7685 4826
rect 7629 4772 7685 4774
rect 4611 4403 4667 4405
rect 4611 4351 4613 4403
rect 4613 4351 4665 4403
rect 4665 4351 4667 4403
rect 4611 4349 4667 4351
rect 5835 3978 5891 3980
rect 5835 3926 5837 3978
rect 5837 3926 5889 3978
rect 5889 3926 5891 3978
rect 5835 3924 5891 3926
rect 4611 3451 4667 3453
rect 4611 3399 4613 3451
rect 4613 3399 4665 3451
rect 4665 3399 4667 3451
rect 4611 3397 4667 3399
rect 5835 3026 5891 3028
rect 5835 2974 5837 3026
rect 5837 2974 5889 3026
rect 5889 2974 5891 3026
rect 5835 2972 5891 2974
rect -1397 2912 -1341 2914
rect 4611 2414 4667 2416
rect 4611 2362 4613 2414
rect 4613 2362 4665 2414
rect 4665 2362 4667 2414
rect 4611 2360 4667 2362
rect 447 1959 503 1961
rect 447 1907 449 1959
rect 449 1907 501 1959
rect 501 1907 503 1959
rect 447 1905 503 1907
rect 5835 1792 5891 1794
rect 5835 1740 5837 1792
rect 5837 1740 5889 1792
rect 5889 1740 5891 1792
rect 5835 1738 5891 1740
rect 4824 1633 4880 1635
rect 4824 1581 4826 1633
rect 4826 1581 4878 1633
rect 4878 1581 4880 1633
rect 4824 1579 4880 1581
rect 5232 1633 5288 1635
rect 5232 1581 5234 1633
rect 5234 1581 5286 1633
rect 5286 1581 5288 1633
rect 5232 1579 5288 1581
rect 5640 1633 5696 1635
rect 5640 1581 5642 1633
rect 5642 1581 5694 1633
rect 5694 1581 5696 1633
rect 5640 1579 5696 1581
rect 14513 1478 14569 1480
rect 14513 1426 14515 1478
rect 14515 1426 14567 1478
rect 14567 1426 14569 1478
rect 14513 1424 14569 1426
rect 24349 1478 24405 1480
rect 24349 1426 24351 1478
rect 24351 1426 24403 1478
rect 24403 1426 24405 1478
rect 24349 1424 24405 1426
rect 14513 562 14569 564
rect 14513 510 14515 562
rect 14515 510 14567 562
rect 14567 510 14569 562
rect 14513 508 14569 510
rect 24349 562 24405 564
rect 24349 510 24351 562
rect 24351 510 24403 562
rect 24403 510 24405 562
rect 24349 508 24405 510
rect 14681 43 14737 45
rect 14681 -9 14683 43
rect 14683 -9 14735 43
rect 14735 -9 14737 43
rect 14681 -11 14737 -9
rect 14989 43 15045 45
rect 14989 -9 14991 43
rect 14991 -9 15043 43
rect 15043 -9 15045 43
rect 14989 -11 15045 -9
rect 15297 43 15353 45
rect 15297 -9 15299 43
rect 15299 -9 15351 43
rect 15351 -9 15353 43
rect 15297 -11 15353 -9
rect 15605 43 15661 45
rect 15605 -9 15607 43
rect 15607 -9 15659 43
rect 15659 -9 15661 43
rect 15605 -11 15661 -9
rect 15913 43 15969 45
rect 15913 -9 15915 43
rect 15915 -9 15967 43
rect 15967 -9 15969 43
rect 15913 -11 15969 -9
rect 16221 43 16277 45
rect 16221 -9 16223 43
rect 16223 -9 16275 43
rect 16275 -9 16277 43
rect 16221 -11 16277 -9
rect 16529 43 16585 45
rect 16529 -9 16531 43
rect 16531 -9 16583 43
rect 16583 -9 16585 43
rect 16529 -11 16585 -9
rect 16837 43 16893 45
rect 16837 -9 16839 43
rect 16839 -9 16891 43
rect 16891 -9 16893 43
rect 16837 -11 16893 -9
rect 17145 43 17201 45
rect 17145 -9 17147 43
rect 17147 -9 17199 43
rect 17199 -9 17201 43
rect 17145 -11 17201 -9
rect 17453 43 17509 45
rect 17453 -9 17455 43
rect 17455 -9 17507 43
rect 17507 -9 17509 43
rect 17453 -11 17509 -9
rect 17761 43 17817 45
rect 17761 -9 17763 43
rect 17763 -9 17815 43
rect 17815 -9 17817 43
rect 17761 -11 17817 -9
rect 18069 43 18125 45
rect 18069 -9 18071 43
rect 18071 -9 18123 43
rect 18123 -9 18125 43
rect 18069 -11 18125 -9
rect 18377 43 18433 45
rect 18377 -9 18379 43
rect 18379 -9 18431 43
rect 18431 -9 18433 43
rect 18377 -11 18433 -9
rect 18685 43 18741 45
rect 18685 -9 18687 43
rect 18687 -9 18739 43
rect 18739 -9 18741 43
rect 18685 -11 18741 -9
rect 18993 43 19049 45
rect 18993 -9 18995 43
rect 18995 -9 19047 43
rect 19047 -9 19049 43
rect 18993 -11 19049 -9
rect 19301 43 19357 45
rect 19301 -9 19303 43
rect 19303 -9 19355 43
rect 19355 -9 19357 43
rect 19301 -11 19357 -9
rect 19609 43 19665 45
rect 19609 -9 19611 43
rect 19611 -9 19663 43
rect 19663 -9 19665 43
rect 19609 -11 19665 -9
rect 19917 43 19973 45
rect 19917 -9 19919 43
rect 19919 -9 19971 43
rect 19971 -9 19973 43
rect 19917 -11 19973 -9
rect 20225 43 20281 45
rect 20225 -9 20227 43
rect 20227 -9 20279 43
rect 20279 -9 20281 43
rect 20225 -11 20281 -9
rect 20533 43 20589 45
rect 20533 -9 20535 43
rect 20535 -9 20587 43
rect 20587 -9 20589 43
rect 20533 -11 20589 -9
rect 20841 43 20897 45
rect 20841 -9 20843 43
rect 20843 -9 20895 43
rect 20895 -9 20897 43
rect 20841 -11 20897 -9
rect 21149 43 21205 45
rect 21149 -9 21151 43
rect 21151 -9 21203 43
rect 21203 -9 21205 43
rect 21149 -11 21205 -9
rect 21457 43 21513 45
rect 21457 -9 21459 43
rect 21459 -9 21511 43
rect 21511 -9 21513 43
rect 21457 -11 21513 -9
rect 21765 43 21821 45
rect 21765 -9 21767 43
rect 21767 -9 21819 43
rect 21819 -9 21821 43
rect 21765 -11 21821 -9
rect 22073 43 22129 45
rect 22073 -9 22075 43
rect 22075 -9 22127 43
rect 22127 -9 22129 43
rect 22073 -11 22129 -9
rect 22381 43 22437 45
rect 22381 -9 22383 43
rect 22383 -9 22435 43
rect 22435 -9 22437 43
rect 22381 -11 22437 -9
rect 22689 43 22745 45
rect 22689 -9 22691 43
rect 22691 -9 22743 43
rect 22743 -9 22745 43
rect 22689 -11 22745 -9
rect 22997 43 23053 45
rect 22997 -9 22999 43
rect 22999 -9 23051 43
rect 23051 -9 23053 43
rect 22997 -11 23053 -9
rect 23305 43 23361 45
rect 23305 -9 23307 43
rect 23307 -9 23359 43
rect 23359 -9 23361 43
rect 23305 -11 23361 -9
rect 23613 43 23669 45
rect 23613 -9 23615 43
rect 23615 -9 23667 43
rect 23667 -9 23669 43
rect 23613 -11 23669 -9
rect 23921 43 23977 45
rect 23921 -9 23923 43
rect 23923 -9 23975 43
rect 23975 -9 23977 43
rect 23921 -11 23977 -9
rect 24229 43 24285 45
rect 24229 -9 24231 43
rect 24231 -9 24283 43
rect 24283 -9 24285 43
rect 24229 -11 24285 -9
<< metal3 >>
rect -1496 13746 62074 13752
rect -1496 13682 -1490 13746
rect -1426 13682 -1354 13746
rect -1290 13682 -1218 13746
rect -1154 13682 61732 13746
rect 61796 13682 61868 13746
rect 61932 13682 62004 13746
rect 62068 13682 62074 13746
rect -1496 13610 62074 13682
rect -1496 13546 -1490 13610
rect -1426 13546 -1354 13610
rect -1290 13546 -1218 13610
rect -1154 13546 61732 13610
rect 61796 13546 61868 13610
rect 61932 13546 62004 13610
rect 62068 13546 62074 13610
rect -1496 13474 62074 13546
rect -1496 13410 -1490 13474
rect -1426 13410 -1354 13474
rect -1290 13410 -1218 13474
rect -1154 13410 11372 13474
rect 11436 13410 24345 13474
rect 24409 13410 49142 13474
rect 49206 13410 60319 13474
rect 60383 13410 61732 13474
rect 61796 13410 61868 13474
rect 61932 13410 62004 13474
rect 62068 13410 62074 13474
rect -1496 13404 62074 13410
rect -800 13050 61378 13056
rect -800 12986 -794 13050
rect -730 12986 -658 13050
rect -594 12986 -522 13050
rect -458 12986 61036 13050
rect 61100 12986 61172 13050
rect 61236 12986 61308 13050
rect 61372 12986 61378 13050
rect -800 12914 61378 12986
rect -800 12850 -794 12914
rect -730 12850 -658 12914
rect -594 12850 -522 12914
rect -458 12850 61036 12914
rect 61100 12850 61172 12914
rect 61236 12850 61308 12914
rect 61372 12850 61378 12914
rect -800 12778 61378 12850
rect -800 12714 -794 12778
rect -730 12714 -658 12778
rect -594 12714 -522 12778
rect -458 12714 11790 12778
rect 11854 12714 24101 12778
rect 24165 12714 34334 12778
rect 34398 12714 36413 12778
rect 36477 12714 48724 12778
rect 48788 12714 60100 12778
rect 60164 12714 61036 12778
rect 61100 12714 61172 12778
rect 61236 12714 61308 12778
rect 61372 12714 61378 12778
rect -800 12708 61378 12714
rect 8184 12234 8282 12245
rect 60232 12234 60330 12245
rect 7070 12228 11860 12234
rect 7070 12224 11790 12228
rect 7070 12168 8205 12224
rect 8261 12168 11790 12224
rect 7070 12164 11790 12168
rect 11854 12164 11860 12228
rect 7070 12158 11860 12164
rect 60094 12228 61106 12234
rect 60094 12164 60100 12228
rect 60164 12224 61036 12228
rect 60164 12168 60253 12224
rect 60309 12168 61036 12224
rect 60164 12164 61036 12168
rect 61100 12164 61106 12228
rect 60094 12158 61106 12164
rect 2714 12026 2812 12034
rect -40 12017 2950 12026
rect -40 11953 2731 12017
rect 2795 11953 2950 12017
rect -40 11950 2950 11953
rect 2576 11947 2950 11950
rect 3962 12017 4060 12034
rect 3962 11953 3979 12017
rect 4043 11953 4060 12017
rect 2714 11936 2812 11947
rect 3962 11936 4060 11953
rect 5560 12023 5658 12034
rect 7070 12023 7146 12158
rect 8184 12147 8282 12158
rect 60232 12147 60330 12158
rect 5560 12017 7146 12023
rect 5560 11953 5577 12017
rect 5641 11953 7146 12017
rect 5560 11947 7146 11953
rect 7208 12023 7306 12034
rect 7208 12017 11442 12023
rect 7208 11953 7225 12017
rect 7289 11953 11372 12017
rect 11436 11953 11442 12017
rect 7208 11947 11442 11953
rect 5560 11936 5658 11947
rect 7208 11936 7306 11947
rect 1219 10352 2598 10428
rect 1219 10290 1295 10352
rect -528 10284 45 10290
rect -528 10220 -522 10284
rect -458 10220 45 10284
rect -528 10214 45 10220
rect 1006 10284 1295 10290
rect 1006 10220 1012 10284
rect 1076 10220 1225 10284
rect 1289 10220 1295 10284
rect 2522 10307 2598 10352
rect 2725 10380 5647 10456
rect 2725 10318 2801 10380
rect 5571 10318 5647 10380
rect 34317 10321 34415 10332
rect 2714 10307 2812 10318
rect 3962 10307 4060 10318
rect 2522 10301 2812 10307
rect 2224 10255 2322 10266
rect 1006 10214 1295 10220
rect 1365 10249 2460 10255
rect 1365 10185 1371 10249
rect 1435 10245 2460 10249
rect 1435 10189 2245 10245
rect 2301 10189 2460 10245
rect 2522 10237 2731 10301
rect 2795 10237 2812 10301
rect 2522 10231 2812 10237
rect 2714 10220 2812 10231
rect 2874 10301 4060 10307
rect 2874 10237 3979 10301
rect 4043 10237 4060 10301
rect 2874 10231 4060 10237
rect 1435 10185 2460 10189
rect 1365 10179 2460 10185
rect 2224 10168 2322 10179
rect 2384 10158 2460 10179
rect 2874 10158 2950 10231
rect 3962 10220 4060 10231
rect 5560 10301 5658 10318
rect 7208 10307 7306 10318
rect 5560 10237 5577 10301
rect 5641 10237 5658 10301
rect 5560 10220 5658 10237
rect 5720 10301 7306 10307
rect 5720 10237 7225 10301
rect 7289 10237 7306 10301
rect 5720 10231 7306 10237
rect 34317 10315 48794 10321
rect 34317 10251 34334 10315
rect 34398 10251 36413 10315
rect 36477 10251 48724 10315
rect 48788 10251 48794 10315
rect 34317 10245 48794 10251
rect 34317 10234 34415 10245
rect 2384 10082 2950 10158
rect 3973 10158 4049 10220
rect 5720 10158 5796 10231
rect 7208 10220 7306 10231
rect 3973 10082 5796 10158
rect 92 9884 190 9895
rect -1224 9878 1441 9884
rect -1224 9814 -1218 9878
rect -1154 9814 109 9878
rect 173 9814 1371 9878
rect 1435 9814 1441 9878
rect -1224 9808 1441 9814
rect 92 9797 190 9808
rect 1316 9459 1414 9470
rect 1006 9453 1552 9459
rect 1006 9389 1012 9453
rect 1076 9389 1184 9453
rect 1248 9449 1482 9453
rect 1248 9393 1337 9449
rect 1393 9393 1482 9449
rect 1248 9389 1482 9393
rect 1546 9389 1552 9453
rect 8082 9448 8180 9459
rect 1006 9383 1552 9389
rect 7219 9442 8180 9448
rect 1316 9372 1414 9383
rect 7219 9378 7225 9442
rect 7289 9378 8099 9442
rect 8163 9378 8180 9442
rect 7219 9372 8180 9378
rect 8082 9361 8180 9372
rect 92 8926 190 8943
rect 92 8862 109 8926
rect 173 8862 190 8926
rect 92 8845 190 8862
rect 8078 8786 8176 8803
rect 60302 8792 60400 8803
rect 8078 8722 8095 8786
rect 8159 8722 8176 8786
rect 8078 8705 8176 8722
rect 49136 8786 61802 8792
rect 49136 8722 49142 8786
rect 49206 8722 60319 8786
rect 60383 8722 61732 8786
rect 61796 8722 61802 8786
rect 49136 8716 61802 8722
rect 60302 8705 60400 8716
rect 1316 8507 1414 8518
rect 1316 8501 1552 8507
rect 1316 8437 1333 8501
rect 1397 8437 1482 8501
rect 1546 8437 1552 8501
rect 1316 8431 1552 8437
rect 1316 8420 1414 8431
rect 92 7895 190 7906
rect -1224 7889 190 7895
rect -1224 7825 -1218 7889
rect -1154 7825 109 7889
rect 173 7825 190 7889
rect 8078 7876 8176 7887
rect 60302 7876 60400 7887
rect -1224 7819 190 7825
rect 92 7808 190 7819
rect 6997 7870 8176 7876
rect 6997 7806 7003 7870
rect 7067 7866 8176 7870
rect 7067 7810 8099 7866
rect 8155 7810 8176 7866
rect 7067 7806 8176 7810
rect 6997 7800 8176 7806
rect 48718 7870 61106 7876
rect 48718 7806 48724 7870
rect 48788 7866 61036 7870
rect 48788 7810 60323 7866
rect 60379 7810 61036 7866
rect 48788 7806 61036 7810
rect 61100 7806 61106 7870
rect 48718 7800 61106 7806
rect 8078 7789 8176 7800
rect 60302 7789 60400 7800
rect -1496 7405 949 7411
rect -1496 7341 879 7405
rect 943 7341 949 7405
rect -1496 7335 949 7341
rect 34249 7374 34347 7385
rect 34249 7368 36483 7374
rect 34249 7304 34266 7368
rect 34330 7304 36413 7368
rect 36477 7304 36483 7368
rect 34249 7298 36483 7304
rect 34249 7287 34347 7298
rect 1316 7273 1414 7284
rect -528 7267 1414 7273
rect -528 7203 -522 7267
rect -458 7203 1333 7267
rect 1397 7203 1414 7267
rect -528 7197 1414 7203
rect 1316 7186 1414 7197
rect 305 7114 403 7125
rect 713 7114 811 7125
rect 1121 7114 1219 7125
rect -1496 7104 403 7114
rect -1496 7048 326 7104
rect 382 7048 403 7104
rect -1496 7038 403 7048
rect 465 7108 811 7114
rect 465 7044 471 7108
rect 535 7104 811 7108
rect 535 7048 734 7104
rect 790 7048 811 7104
rect 535 7044 811 7048
rect 465 7038 811 7044
rect 873 7108 1219 7114
rect 873 7044 879 7108
rect 943 7104 1219 7108
rect 943 7048 1142 7104
rect 1198 7048 1219 7104
rect 943 7044 1219 7048
rect 873 7038 1219 7044
rect 305 7027 403 7038
rect 713 7027 811 7038
rect 1121 7027 1219 7038
rect 1355 6958 1453 6969
rect -528 6952 4534 6958
rect -528 6888 -522 6952
rect -458 6888 1372 6952
rect 1436 6888 4464 6952
rect 4528 6888 4534 6952
rect -528 6882 4534 6888
rect 1355 6871 1453 6882
rect -1496 6814 541 6820
rect -1496 6750 471 6814
rect 535 6750 541 6814
rect -1496 6744 541 6750
rect 6986 6557 7084 6565
rect 4458 6551 7222 6557
rect 4458 6487 4464 6551
rect 4528 6548 7222 6551
rect 4528 6487 7003 6548
rect 4458 6484 7003 6487
rect 7067 6484 7222 6548
rect 4458 6481 7222 6484
rect 6848 6478 7222 6481
rect 7608 6554 7706 6565
rect 7608 6548 8165 6554
rect 7608 6484 7625 6548
rect 7689 6484 8095 6548
rect 8159 6484 8165 6548
rect 7608 6478 8165 6484
rect 6986 6467 7084 6478
rect 7608 6467 7706 6478
rect 5717 4911 7073 4987
rect 5717 4821 5793 4911
rect 6997 4849 7073 4911
rect 4458 4815 5793 4821
rect 4458 4751 5510 4815
rect 5574 4751 5723 4815
rect 5787 4751 5793 4815
rect 6986 4832 7084 4849
rect 7608 4838 7706 4849
rect 6722 4786 6820 4797
rect 4458 4745 5793 4751
rect 5863 4780 6820 4786
rect 5863 4716 5869 4780
rect 5933 4776 6820 4780
rect 5933 4720 6743 4776
rect 6799 4720 6820 4776
rect 6986 4768 7003 4832
rect 7067 4768 7084 4832
rect 6986 4751 7084 4768
rect 7146 4832 7706 4838
rect 7146 4768 7625 4832
rect 7689 4768 7706 4832
rect 7146 4762 7706 4768
rect 5933 4716 6820 4720
rect 5863 4710 6820 4716
rect 6722 4699 6820 4710
rect 6733 4637 6809 4699
rect 7146 4637 7222 4762
rect 7608 4751 7706 4762
rect 6733 4561 7222 4637
rect 4590 4415 4688 4426
rect 4590 4409 5939 4415
rect 4590 4345 4607 4409
rect 4671 4345 5869 4409
rect 5933 4345 5939 4409
rect -601 4329 -503 4340
rect -1224 4323 -503 4329
rect 4590 4339 5939 4345
rect 4590 4328 4688 4339
rect -1224 4259 -1218 4323
rect -1154 4259 -503 4323
rect -1224 4253 -503 4259
rect -601 4242 -503 4253
rect 5814 3990 5912 4001
rect 5504 3984 6050 3990
rect 5504 3920 5510 3984
rect 5574 3920 5682 3984
rect 5746 3980 5980 3984
rect 5746 3924 5835 3980
rect 5891 3924 5980 3980
rect 5746 3920 5980 3924
rect 6044 3920 6050 3984
rect 5504 3914 6050 3920
rect 5814 3903 5912 3914
rect 4590 3457 4688 3474
rect 4590 3393 4607 3457
rect 4671 3393 4688 3457
rect 4590 3376 4688 3393
rect 5814 3038 5912 3049
rect 5814 3032 6050 3038
rect -1418 2978 -1320 2989
rect -1496 2968 -1320 2978
rect -1496 2912 -1397 2968
rect -1341 2912 -1320 2968
rect 5814 2968 5831 3032
rect 5895 2968 5980 3032
rect 6044 2968 6050 3032
rect 5814 2962 6050 2968
rect 5814 2951 5912 2962
rect -1496 2902 -1320 2912
rect -1418 2891 -1320 2902
rect 4590 2420 4688 2437
rect 4590 2356 4607 2420
rect 4671 2356 4688 2420
rect 4590 2339 4688 2356
rect 426 1971 524 1982
rect -1496 1961 524 1971
rect -1496 1905 447 1961
rect 503 1905 524 1961
rect -1496 1895 524 1905
rect 426 1884 524 1895
rect 5814 1804 5912 1815
rect 5814 1798 11860 1804
rect 5814 1734 5831 1798
rect 5895 1734 11790 1798
rect 11854 1734 11860 1798
rect 5814 1728 11860 1734
rect 5814 1717 5912 1728
rect -601 1701 -503 1712
rect -800 1695 -503 1701
rect -800 1631 -794 1695
rect -730 1631 -503 1695
rect -800 1625 -503 1631
rect -601 1614 -503 1625
rect 4803 1639 4901 1656
rect 4803 1575 4820 1639
rect 4884 1575 4901 1639
rect 4803 1558 4901 1575
rect 5211 1639 5309 1656
rect 5211 1575 5228 1639
rect 5292 1575 5309 1639
rect 5211 1558 5309 1575
rect 5619 1639 5717 1656
rect 5619 1575 5636 1639
rect 5700 1575 5717 1639
rect 5619 1558 5717 1575
rect 14492 1490 14590 1501
rect 24328 1490 24426 1501
rect 14354 1484 24426 1490
rect 14354 1420 14360 1484
rect 14424 1480 24101 1484
rect 14424 1424 14513 1480
rect 14569 1424 24101 1480
rect 14424 1420 24101 1424
rect 24165 1480 24426 1484
rect 24165 1424 24349 1480
rect 24405 1424 24426 1480
rect 24165 1420 24426 1424
rect 14354 1414 24426 1420
rect 14492 1403 14590 1414
rect 24328 1403 24426 1414
rect 14492 574 14590 585
rect 24328 574 24426 585
rect 14492 568 24032 574
rect 14492 504 14509 568
rect 14573 504 23962 568
rect 24026 504 24032 568
rect 14492 498 24032 504
rect 24328 568 36622 574
rect 24328 504 24345 568
rect 24409 504 36552 568
rect 36616 504 36622 568
rect 24328 498 36622 504
rect 14492 487 14590 498
rect 24328 487 24426 498
rect 14660 49 14758 66
rect 14660 -15 14677 49
rect 14741 -15 14758 49
rect 14660 -32 14758 -15
rect 14968 49 15066 66
rect 14968 -15 14985 49
rect 15049 -15 15066 49
rect 14968 -32 15066 -15
rect 15276 49 15374 66
rect 15276 -15 15293 49
rect 15357 -15 15374 49
rect 15276 -32 15374 -15
rect 15584 49 15682 66
rect 15584 -15 15601 49
rect 15665 -15 15682 49
rect 15584 -32 15682 -15
rect 15892 49 15990 66
rect 15892 -15 15909 49
rect 15973 -15 15990 49
rect 15892 -32 15990 -15
rect 16200 49 16298 66
rect 16200 -15 16217 49
rect 16281 -15 16298 49
rect 16200 -32 16298 -15
rect 16508 49 16606 66
rect 16508 -15 16525 49
rect 16589 -15 16606 49
rect 16508 -32 16606 -15
rect 16816 49 16914 66
rect 16816 -15 16833 49
rect 16897 -15 16914 49
rect 16816 -32 16914 -15
rect 17124 49 17222 66
rect 17124 -15 17141 49
rect 17205 -15 17222 49
rect 17124 -32 17222 -15
rect 17432 49 17530 66
rect 17432 -15 17449 49
rect 17513 -15 17530 49
rect 17432 -32 17530 -15
rect 17740 49 17838 66
rect 17740 -15 17757 49
rect 17821 -15 17838 49
rect 17740 -32 17838 -15
rect 18048 49 18146 66
rect 18048 -15 18065 49
rect 18129 -15 18146 49
rect 18048 -32 18146 -15
rect 18356 49 18454 66
rect 18356 -15 18373 49
rect 18437 -15 18454 49
rect 18356 -32 18454 -15
rect 18664 49 18762 66
rect 18664 -15 18681 49
rect 18745 -15 18762 49
rect 18664 -32 18762 -15
rect 18972 49 19070 66
rect 18972 -15 18989 49
rect 19053 -15 19070 49
rect 18972 -32 19070 -15
rect 19280 49 19378 66
rect 19280 -15 19297 49
rect 19361 -15 19378 49
rect 19280 -32 19378 -15
rect 19588 49 19686 66
rect 19588 -15 19605 49
rect 19669 -15 19686 49
rect 19588 -32 19686 -15
rect 19896 49 19994 66
rect 19896 -15 19913 49
rect 19977 -15 19994 49
rect 19896 -32 19994 -15
rect 20204 49 20302 66
rect 20204 -15 20221 49
rect 20285 -15 20302 49
rect 20204 -32 20302 -15
rect 20512 49 20610 66
rect 20512 -15 20529 49
rect 20593 -15 20610 49
rect 20512 -32 20610 -15
rect 20820 49 20918 66
rect 20820 -15 20837 49
rect 20901 -15 20918 49
rect 20820 -32 20918 -15
rect 21128 49 21226 66
rect 21128 -15 21145 49
rect 21209 -15 21226 49
rect 21128 -32 21226 -15
rect 21436 49 21534 66
rect 21436 -15 21453 49
rect 21517 -15 21534 49
rect 21436 -32 21534 -15
rect 21744 49 21842 66
rect 21744 -15 21761 49
rect 21825 -15 21842 49
rect 21744 -32 21842 -15
rect 22052 49 22150 66
rect 22052 -15 22069 49
rect 22133 -15 22150 49
rect 22052 -32 22150 -15
rect 22360 49 22458 66
rect 22360 -15 22377 49
rect 22441 -15 22458 49
rect 22360 -32 22458 -15
rect 22668 49 22766 66
rect 22668 -15 22685 49
rect 22749 -15 22766 49
rect 22668 -32 22766 -15
rect 22976 49 23074 66
rect 22976 -15 22993 49
rect 23057 -15 23074 49
rect 22976 -32 23074 -15
rect 23284 49 23382 66
rect 23284 -15 23301 49
rect 23365 -15 23382 49
rect 23284 -32 23382 -15
rect 23592 49 23690 66
rect 23900 55 23998 66
rect 23592 -15 23609 49
rect 23673 -15 23690 49
rect 23592 -32 23690 -15
rect 23762 49 23998 55
rect 23762 -15 23768 49
rect 23832 45 23998 49
rect 23832 -11 23921 45
rect 23977 -11 23998 45
rect 23832 -15 23998 -11
rect 23762 -21 23998 -15
rect 23900 -32 23998 -21
rect 24208 55 24306 66
rect 24208 49 24553 55
rect 24208 45 24483 49
rect 24208 -11 24229 45
rect 24285 -11 24483 45
rect 24208 -15 24483 -11
rect 24547 -15 24553 49
rect 24208 -21 24553 -15
rect 24208 -32 24306 -21
rect -800 -458 61378 -452
rect -800 -522 -794 -458
rect -730 -522 -658 -458
rect -594 -522 -522 -458
rect -458 -522 11790 -458
rect 11854 -522 14360 -458
rect 14424 -522 24101 -458
rect 24165 -522 36413 -458
rect 36477 -522 48724 -458
rect 48788 -522 61036 -458
rect 61100 -522 61172 -458
rect 61236 -522 61308 -458
rect 61372 -522 61378 -458
rect -800 -594 61378 -522
rect -800 -658 -794 -594
rect -730 -658 -658 -594
rect -594 -658 -522 -594
rect -458 -658 61036 -594
rect 61100 -658 61172 -594
rect 61236 -658 61308 -594
rect 61372 -658 61378 -594
rect -800 -730 61378 -658
rect -800 -794 -794 -730
rect -730 -794 -658 -730
rect -594 -794 -522 -730
rect -458 -794 61036 -730
rect 61100 -794 61172 -730
rect 61236 -794 61308 -730
rect 61372 -794 61378 -730
rect -800 -800 61378 -794
rect -1496 -1154 62074 -1148
rect -1496 -1218 -1490 -1154
rect -1426 -1218 -1354 -1154
rect -1290 -1218 -1218 -1154
rect -1154 -1218 7625 -1154
rect 7689 -1218 14509 -1154
rect 14573 -1218 23962 -1154
rect 24026 -1218 24345 -1154
rect 24409 -1218 36552 -1154
rect 36616 -1218 49142 -1154
rect 49206 -1218 61732 -1154
rect 61796 -1218 61868 -1154
rect 61932 -1218 62004 -1154
rect 62068 -1218 62074 -1154
rect -1496 -1290 62074 -1218
rect -1496 -1354 -1490 -1290
rect -1426 -1354 -1354 -1290
rect -1290 -1354 -1218 -1290
rect -1154 -1354 61732 -1290
rect 61796 -1354 61868 -1290
rect 61932 -1354 62004 -1290
rect 62068 -1354 62074 -1290
rect -1496 -1426 62074 -1354
rect -1496 -1490 -1490 -1426
rect -1426 -1490 -1354 -1426
rect -1290 -1490 -1218 -1426
rect -1154 -1490 61732 -1426
rect 61796 -1490 61868 -1426
rect 61932 -1490 62004 -1426
rect 62068 -1490 62074 -1426
rect -1496 -1496 62074 -1490
<< via3 >>
rect -1490 13682 -1426 13746
rect -1354 13682 -1290 13746
rect -1218 13682 -1154 13746
rect 61732 13682 61796 13746
rect 61868 13682 61932 13746
rect 62004 13682 62068 13746
rect -1490 13546 -1426 13610
rect -1354 13546 -1290 13610
rect -1218 13546 -1154 13610
rect 61732 13546 61796 13610
rect 61868 13546 61932 13610
rect 62004 13546 62068 13610
rect -1490 13410 -1426 13474
rect -1354 13410 -1290 13474
rect -1218 13410 -1154 13474
rect 11372 13410 11436 13474
rect 24345 13410 24409 13474
rect 49142 13410 49206 13474
rect 60319 13410 60383 13474
rect 61732 13410 61796 13474
rect 61868 13410 61932 13474
rect 62004 13410 62068 13474
rect -794 12986 -730 13050
rect -658 12986 -594 13050
rect -522 12986 -458 13050
rect 61036 12986 61100 13050
rect 61172 12986 61236 13050
rect 61308 12986 61372 13050
rect -794 12850 -730 12914
rect -658 12850 -594 12914
rect -522 12850 -458 12914
rect 61036 12850 61100 12914
rect 61172 12850 61236 12914
rect 61308 12850 61372 12914
rect -794 12714 -730 12778
rect -658 12714 -594 12778
rect -522 12714 -458 12778
rect 11790 12714 11854 12778
rect 24101 12714 24165 12778
rect 34334 12714 34398 12778
rect 36413 12714 36477 12778
rect 48724 12714 48788 12778
rect 60100 12714 60164 12778
rect 61036 12714 61100 12778
rect 61172 12714 61236 12778
rect 61308 12714 61372 12778
rect 11790 12164 11854 12228
rect 60100 12164 60164 12228
rect 61036 12164 61100 12228
rect 2731 12013 2795 12017
rect 2731 11957 2735 12013
rect 2735 11957 2791 12013
rect 2791 11957 2795 12013
rect 2731 11953 2795 11957
rect 3979 12013 4043 12017
rect 3979 11957 3983 12013
rect 3983 11957 4039 12013
rect 4039 11957 4043 12013
rect 3979 11953 4043 11957
rect 5577 12013 5641 12017
rect 5577 11957 5581 12013
rect 5581 11957 5637 12013
rect 5637 11957 5641 12013
rect 5577 11953 5641 11957
rect 7225 12013 7289 12017
rect 7225 11957 7229 12013
rect 7229 11957 7285 12013
rect 7285 11957 7289 12013
rect 7225 11953 7289 11957
rect 11372 11953 11436 12017
rect -522 10220 -458 10284
rect 1012 10220 1076 10284
rect 1225 10220 1289 10284
rect 1371 10185 1435 10249
rect 2731 10297 2795 10301
rect 2731 10241 2735 10297
rect 2735 10241 2791 10297
rect 2791 10241 2795 10297
rect 2731 10237 2795 10241
rect 3979 10297 4043 10301
rect 3979 10241 3983 10297
rect 3983 10241 4039 10297
rect 4039 10241 4043 10297
rect 3979 10237 4043 10241
rect 5577 10297 5641 10301
rect 5577 10241 5581 10297
rect 5581 10241 5637 10297
rect 5637 10241 5641 10297
rect 5577 10237 5641 10241
rect 7225 10297 7289 10301
rect 7225 10241 7229 10297
rect 7229 10241 7285 10297
rect 7285 10241 7289 10297
rect 7225 10237 7289 10241
rect 34334 10311 34398 10315
rect 34334 10255 34338 10311
rect 34338 10255 34394 10311
rect 34394 10255 34398 10311
rect 34334 10251 34398 10255
rect 36413 10251 36477 10315
rect 48724 10251 48788 10315
rect -1218 9814 -1154 9878
rect 109 9874 173 9878
rect 109 9818 113 9874
rect 113 9818 169 9874
rect 169 9818 173 9874
rect 109 9814 173 9818
rect 1371 9814 1435 9878
rect 1012 9389 1076 9453
rect 1184 9389 1248 9453
rect 1482 9389 1546 9453
rect 7225 9378 7289 9442
rect 8099 9438 8163 9442
rect 8099 9382 8103 9438
rect 8103 9382 8159 9438
rect 8159 9382 8163 9438
rect 8099 9378 8163 9382
rect 109 8922 173 8926
rect 109 8866 113 8922
rect 113 8866 169 8922
rect 169 8866 173 8922
rect 109 8862 173 8866
rect 8095 8782 8159 8786
rect 8095 8726 8099 8782
rect 8099 8726 8155 8782
rect 8155 8726 8159 8782
rect 8095 8722 8159 8726
rect 49142 8722 49206 8786
rect 60319 8782 60383 8786
rect 60319 8726 60323 8782
rect 60323 8726 60379 8782
rect 60379 8726 60383 8782
rect 60319 8722 60383 8726
rect 61732 8722 61796 8786
rect 1333 8497 1397 8501
rect 1333 8441 1337 8497
rect 1337 8441 1393 8497
rect 1393 8441 1397 8497
rect 1333 8437 1397 8441
rect 1482 8437 1546 8501
rect -1218 7825 -1154 7889
rect 109 7885 173 7889
rect 109 7829 113 7885
rect 113 7829 169 7885
rect 169 7829 173 7885
rect 109 7825 173 7829
rect 7003 7806 7067 7870
rect 48724 7806 48788 7870
rect 61036 7806 61100 7870
rect 879 7341 943 7405
rect 34266 7364 34330 7368
rect 34266 7308 34270 7364
rect 34270 7308 34326 7364
rect 34326 7308 34330 7364
rect 34266 7304 34330 7308
rect 36413 7304 36477 7368
rect -522 7203 -458 7267
rect 1333 7263 1397 7267
rect 1333 7207 1337 7263
rect 1337 7207 1393 7263
rect 1393 7207 1397 7263
rect 1333 7203 1397 7207
rect 471 7044 535 7108
rect 879 7044 943 7108
rect -522 6888 -458 6952
rect 1372 6888 1436 6952
rect 4464 6888 4528 6952
rect 471 6750 535 6814
rect 4464 6487 4528 6551
rect 7003 6544 7067 6548
rect 7003 6488 7007 6544
rect 7007 6488 7063 6544
rect 7063 6488 7067 6544
rect 7003 6484 7067 6488
rect 7625 6544 7689 6548
rect 7625 6488 7629 6544
rect 7629 6488 7685 6544
rect 7685 6488 7689 6544
rect 7625 6484 7689 6488
rect 8095 6484 8159 6548
rect 5510 4751 5574 4815
rect 5723 4751 5787 4815
rect 5869 4716 5933 4780
rect 7003 4828 7067 4832
rect 7003 4772 7007 4828
rect 7007 4772 7063 4828
rect 7063 4772 7067 4828
rect 7003 4768 7067 4772
rect 7625 4828 7689 4832
rect 7625 4772 7629 4828
rect 7629 4772 7685 4828
rect 7685 4772 7689 4828
rect 7625 4768 7689 4772
rect 4607 4405 4671 4409
rect 4607 4349 4611 4405
rect 4611 4349 4667 4405
rect 4667 4349 4671 4405
rect 4607 4345 4671 4349
rect 5869 4345 5933 4409
rect -1218 4259 -1154 4323
rect 5510 3920 5574 3984
rect 5682 3920 5746 3984
rect 5980 3920 6044 3984
rect 4607 3453 4671 3457
rect 4607 3397 4611 3453
rect 4611 3397 4667 3453
rect 4667 3397 4671 3453
rect 4607 3393 4671 3397
rect 5831 3028 5895 3032
rect 5831 2972 5835 3028
rect 5835 2972 5891 3028
rect 5891 2972 5895 3028
rect 5831 2968 5895 2972
rect 5980 2968 6044 3032
rect 4607 2416 4671 2420
rect 4607 2360 4611 2416
rect 4611 2360 4667 2416
rect 4667 2360 4671 2416
rect 4607 2356 4671 2360
rect 5831 1794 5895 1798
rect 5831 1738 5835 1794
rect 5835 1738 5891 1794
rect 5891 1738 5895 1794
rect 5831 1734 5895 1738
rect 11790 1734 11854 1798
rect -794 1631 -730 1695
rect 4820 1635 4884 1639
rect 4820 1579 4824 1635
rect 4824 1579 4880 1635
rect 4880 1579 4884 1635
rect 4820 1575 4884 1579
rect 5228 1635 5292 1639
rect 5228 1579 5232 1635
rect 5232 1579 5288 1635
rect 5288 1579 5292 1635
rect 5228 1575 5292 1579
rect 5636 1635 5700 1639
rect 5636 1579 5640 1635
rect 5640 1579 5696 1635
rect 5696 1579 5700 1635
rect 5636 1575 5700 1579
rect 14360 1420 14424 1484
rect 24101 1420 24165 1484
rect 14509 564 14573 568
rect 14509 508 14513 564
rect 14513 508 14569 564
rect 14569 508 14573 564
rect 14509 504 14573 508
rect 23962 504 24026 568
rect 24345 564 24409 568
rect 24345 508 24349 564
rect 24349 508 24405 564
rect 24405 508 24409 564
rect 24345 504 24409 508
rect 36552 504 36616 568
rect 14677 45 14741 49
rect 14677 -11 14681 45
rect 14681 -11 14737 45
rect 14737 -11 14741 45
rect 14677 -15 14741 -11
rect 14985 45 15049 49
rect 14985 -11 14989 45
rect 14989 -11 15045 45
rect 15045 -11 15049 45
rect 14985 -15 15049 -11
rect 15293 45 15357 49
rect 15293 -11 15297 45
rect 15297 -11 15353 45
rect 15353 -11 15357 45
rect 15293 -15 15357 -11
rect 15601 45 15665 49
rect 15601 -11 15605 45
rect 15605 -11 15661 45
rect 15661 -11 15665 45
rect 15601 -15 15665 -11
rect 15909 45 15973 49
rect 15909 -11 15913 45
rect 15913 -11 15969 45
rect 15969 -11 15973 45
rect 15909 -15 15973 -11
rect 16217 45 16281 49
rect 16217 -11 16221 45
rect 16221 -11 16277 45
rect 16277 -11 16281 45
rect 16217 -15 16281 -11
rect 16525 45 16589 49
rect 16525 -11 16529 45
rect 16529 -11 16585 45
rect 16585 -11 16589 45
rect 16525 -15 16589 -11
rect 16833 45 16897 49
rect 16833 -11 16837 45
rect 16837 -11 16893 45
rect 16893 -11 16897 45
rect 16833 -15 16897 -11
rect 17141 45 17205 49
rect 17141 -11 17145 45
rect 17145 -11 17201 45
rect 17201 -11 17205 45
rect 17141 -15 17205 -11
rect 17449 45 17513 49
rect 17449 -11 17453 45
rect 17453 -11 17509 45
rect 17509 -11 17513 45
rect 17449 -15 17513 -11
rect 17757 45 17821 49
rect 17757 -11 17761 45
rect 17761 -11 17817 45
rect 17817 -11 17821 45
rect 17757 -15 17821 -11
rect 18065 45 18129 49
rect 18065 -11 18069 45
rect 18069 -11 18125 45
rect 18125 -11 18129 45
rect 18065 -15 18129 -11
rect 18373 45 18437 49
rect 18373 -11 18377 45
rect 18377 -11 18433 45
rect 18433 -11 18437 45
rect 18373 -15 18437 -11
rect 18681 45 18745 49
rect 18681 -11 18685 45
rect 18685 -11 18741 45
rect 18741 -11 18745 45
rect 18681 -15 18745 -11
rect 18989 45 19053 49
rect 18989 -11 18993 45
rect 18993 -11 19049 45
rect 19049 -11 19053 45
rect 18989 -15 19053 -11
rect 19297 45 19361 49
rect 19297 -11 19301 45
rect 19301 -11 19357 45
rect 19357 -11 19361 45
rect 19297 -15 19361 -11
rect 19605 45 19669 49
rect 19605 -11 19609 45
rect 19609 -11 19665 45
rect 19665 -11 19669 45
rect 19605 -15 19669 -11
rect 19913 45 19977 49
rect 19913 -11 19917 45
rect 19917 -11 19973 45
rect 19973 -11 19977 45
rect 19913 -15 19977 -11
rect 20221 45 20285 49
rect 20221 -11 20225 45
rect 20225 -11 20281 45
rect 20281 -11 20285 45
rect 20221 -15 20285 -11
rect 20529 45 20593 49
rect 20529 -11 20533 45
rect 20533 -11 20589 45
rect 20589 -11 20593 45
rect 20529 -15 20593 -11
rect 20837 45 20901 49
rect 20837 -11 20841 45
rect 20841 -11 20897 45
rect 20897 -11 20901 45
rect 20837 -15 20901 -11
rect 21145 45 21209 49
rect 21145 -11 21149 45
rect 21149 -11 21205 45
rect 21205 -11 21209 45
rect 21145 -15 21209 -11
rect 21453 45 21517 49
rect 21453 -11 21457 45
rect 21457 -11 21513 45
rect 21513 -11 21517 45
rect 21453 -15 21517 -11
rect 21761 45 21825 49
rect 21761 -11 21765 45
rect 21765 -11 21821 45
rect 21821 -11 21825 45
rect 21761 -15 21825 -11
rect 22069 45 22133 49
rect 22069 -11 22073 45
rect 22073 -11 22129 45
rect 22129 -11 22133 45
rect 22069 -15 22133 -11
rect 22377 45 22441 49
rect 22377 -11 22381 45
rect 22381 -11 22437 45
rect 22437 -11 22441 45
rect 22377 -15 22441 -11
rect 22685 45 22749 49
rect 22685 -11 22689 45
rect 22689 -11 22745 45
rect 22745 -11 22749 45
rect 22685 -15 22749 -11
rect 22993 45 23057 49
rect 22993 -11 22997 45
rect 22997 -11 23053 45
rect 23053 -11 23057 45
rect 22993 -15 23057 -11
rect 23301 45 23365 49
rect 23301 -11 23305 45
rect 23305 -11 23361 45
rect 23361 -11 23365 45
rect 23301 -15 23365 -11
rect 23609 45 23673 49
rect 23609 -11 23613 45
rect 23613 -11 23669 45
rect 23669 -11 23673 45
rect 23609 -15 23673 -11
rect 23768 -15 23832 49
rect 24483 -15 24547 49
rect -794 -522 -730 -458
rect -658 -522 -594 -458
rect -522 -522 -458 -458
rect 11790 -522 11854 -458
rect 14360 -522 14424 -458
rect 24101 -522 24165 -458
rect 36413 -522 36477 -458
rect 48724 -522 48788 -458
rect 61036 -522 61100 -458
rect 61172 -522 61236 -458
rect 61308 -522 61372 -458
rect -794 -658 -730 -594
rect -658 -658 -594 -594
rect -522 -658 -458 -594
rect 61036 -658 61100 -594
rect 61172 -658 61236 -594
rect 61308 -658 61372 -594
rect -794 -794 -730 -730
rect -658 -794 -594 -730
rect -522 -794 -458 -730
rect 61036 -794 61100 -730
rect 61172 -794 61236 -730
rect 61308 -794 61372 -730
rect -1490 -1218 -1426 -1154
rect -1354 -1218 -1290 -1154
rect -1218 -1218 -1154 -1154
rect 7625 -1218 7689 -1154
rect 14509 -1218 14573 -1154
rect 23962 -1218 24026 -1154
rect 24345 -1218 24409 -1154
rect 36552 -1218 36616 -1154
rect 49142 -1218 49206 -1154
rect 61732 -1218 61796 -1154
rect 61868 -1218 61932 -1154
rect 62004 -1218 62068 -1154
rect -1490 -1354 -1426 -1290
rect -1354 -1354 -1290 -1290
rect -1218 -1354 -1154 -1290
rect 61732 -1354 61796 -1290
rect 61868 -1354 61932 -1290
rect 62004 -1354 62068 -1290
rect -1490 -1490 -1426 -1426
rect -1354 -1490 -1290 -1426
rect -1218 -1490 -1154 -1426
rect 61732 -1490 61796 -1426
rect 61868 -1490 61932 -1426
rect 62004 -1490 62068 -1426
<< metal4 >>
rect -1496 13746 -1148 13752
rect -1496 13682 -1490 13746
rect -1426 13682 -1354 13746
rect -1290 13682 -1218 13746
rect -1154 13682 -1148 13746
rect -1496 13610 -1148 13682
rect -1496 13546 -1490 13610
rect -1426 13546 -1354 13610
rect -1290 13546 -1218 13610
rect -1154 13546 -1148 13610
rect -1496 13474 -1148 13546
rect 61726 13746 62074 13752
rect 61726 13682 61732 13746
rect 61796 13682 61868 13746
rect 61932 13682 62004 13746
rect 62068 13682 62074 13746
rect 61726 13610 62074 13682
rect 61726 13546 61732 13610
rect 61796 13546 61868 13610
rect 61932 13546 62004 13610
rect 62068 13546 62074 13610
rect -1496 13410 -1490 13474
rect -1426 13410 -1354 13474
rect -1290 13410 -1218 13474
rect -1154 13410 -1148 13474
rect -1496 9878 -1148 13410
rect 11366 13474 11442 13480
rect 11366 13410 11372 13474
rect 11436 13410 11442 13474
rect -1496 9814 -1218 9878
rect -1154 9814 -1148 9878
rect -1496 7889 -1148 9814
rect -1496 7825 -1218 7889
rect -1154 7825 -1148 7889
rect -1496 4323 -1148 7825
rect -1496 4259 -1218 4323
rect -1154 4259 -1148 4323
rect -1496 -1154 -1148 4259
rect -800 13050 -452 13056
rect -800 12986 -794 13050
rect -730 12986 -658 13050
rect -594 12986 -522 13050
rect -458 12986 -452 13050
rect -800 12914 -452 12986
rect -800 12850 -794 12914
rect -730 12850 -658 12914
rect -594 12850 -522 12914
rect -458 12850 -452 12914
rect -800 12778 -452 12850
rect -800 12714 -794 12778
rect -730 12714 -658 12778
rect -594 12714 -522 12778
rect -458 12714 -452 12778
rect -800 10284 -452 12714
rect 2725 12017 2801 12023
rect 2725 11953 2731 12017
rect 2795 11953 2801 12017
rect 2725 10301 2801 11953
rect -800 10220 -522 10284
rect -458 10220 -452 10284
rect -800 7267 -452 10220
rect 1006 10284 1082 10290
rect 1006 10220 1012 10284
rect 1076 10220 1082 10284
rect 103 9878 179 9884
rect 103 9814 109 9878
rect 173 9814 179 9878
rect 103 8926 179 9814
rect 1006 9453 1082 10220
rect 1219 10284 1295 10290
rect 1219 10220 1225 10284
rect 1289 10220 1295 10284
rect 1219 9459 1295 10220
rect 1365 10249 1441 10255
rect 1365 10185 1371 10249
rect 1435 10185 1441 10249
rect 2725 10237 2731 10301
rect 2795 10237 2801 10301
rect 2725 10231 2801 10237
rect 3973 12017 4049 12023
rect 3973 11953 3979 12017
rect 4043 11953 4049 12017
rect 3973 10301 4049 11953
rect 3973 10237 3979 10301
rect 4043 10237 4049 10301
rect 3973 10231 4049 10237
rect 5571 12017 5647 12023
rect 5571 11953 5577 12017
rect 5641 11953 5647 12017
rect 5571 10301 5647 11953
rect 5571 10237 5577 10301
rect 5641 10237 5647 10301
rect 5571 10231 5647 10237
rect 7219 12017 7295 12023
rect 7219 11953 7225 12017
rect 7289 11953 7295 12017
rect 7219 10301 7295 11953
rect 11366 12017 11442 13410
rect 24339 13474 24415 13480
rect 24339 13410 24345 13474
rect 24409 13410 24415 13474
rect 11784 12778 11860 12784
rect 11784 12714 11790 12778
rect 11854 12714 11860 12778
rect 11784 12228 11860 12714
rect 11784 12164 11790 12228
rect 11854 12164 11860 12228
rect 11784 12158 11860 12164
rect 24095 12778 24171 12784
rect 24095 12714 24101 12778
rect 24165 12714 24171 12778
rect 11366 11953 11372 12017
rect 11436 11953 11442 12017
rect 11366 11947 11442 11953
rect 7219 10237 7225 10301
rect 7289 10237 7295 10301
rect 1365 9878 1441 10185
rect 1365 9814 1371 9878
rect 1435 9814 1441 9878
rect 1365 9808 1441 9814
rect 1006 9389 1012 9453
rect 1076 9389 1082 9453
rect 1006 9383 1082 9389
rect 1178 9453 1295 9459
rect 1178 9389 1184 9453
rect 1248 9389 1295 9453
rect 1178 9383 1295 9389
rect 1476 9453 1552 9459
rect 1476 9389 1482 9453
rect 1546 9389 1552 9453
rect 103 8862 109 8926
rect 173 8862 179 8926
rect 103 7889 179 8862
rect 103 7825 109 7889
rect 173 7825 179 7889
rect 103 7819 179 7825
rect 1327 8501 1403 8507
rect 1327 8437 1333 8501
rect 1397 8437 1403 8501
rect -800 7203 -522 7267
rect -458 7203 -452 7267
rect -800 6952 -452 7203
rect 873 7405 949 7411
rect 873 7341 879 7405
rect 943 7341 949 7405
rect -800 6888 -522 6952
rect -458 6888 -452 6952
rect -800 1695 -452 6888
rect 465 7108 541 7114
rect 465 7044 471 7108
rect 535 7044 541 7108
rect 465 6814 541 7044
rect 873 7108 949 7341
rect 873 7044 879 7108
rect 943 7044 949 7108
rect 873 7038 949 7044
rect 1327 7267 1403 8437
rect 1476 8501 1552 9389
rect 7219 9442 7295 10237
rect 7219 9378 7225 9442
rect 7289 9378 7295 9442
rect 7219 9372 7295 9378
rect 8089 9442 8169 9448
rect 8089 9378 8099 9442
rect 8163 9378 8169 9442
rect 8089 9372 8169 9378
rect 1476 8437 1482 8501
rect 1546 8437 1552 8501
rect 1476 8431 1552 8437
rect 8089 8786 8165 9372
rect 8089 8722 8095 8786
rect 8159 8722 8165 8786
rect 1327 7203 1333 7267
rect 1397 7203 1403 7267
rect 1327 6958 1403 7203
rect 6997 7870 7073 7876
rect 6997 7806 7003 7870
rect 7067 7806 7073 7870
rect 1327 6952 1442 6958
rect 1327 6888 1372 6952
rect 1436 6888 1442 6952
rect 1327 6882 1442 6888
rect 4458 6952 4534 6958
rect 4458 6888 4464 6952
rect 4528 6888 4534 6952
rect 465 6750 471 6814
rect 535 6750 541 6814
rect 465 6744 541 6750
rect 4458 6551 4534 6888
rect 4458 6487 4464 6551
rect 4528 6487 4534 6551
rect 4458 6481 4534 6487
rect 6997 6548 7073 7806
rect 6997 6484 7003 6548
rect 7067 6484 7073 6548
rect 6997 4832 7073 6484
rect 5504 4815 5580 4821
rect 5504 4751 5510 4815
rect 5574 4751 5580 4815
rect 4601 4409 4677 4415
rect 4601 4345 4607 4409
rect 4671 4345 4677 4409
rect 4601 3457 4677 4345
rect 5504 3984 5580 4751
rect 5717 4815 5793 4821
rect 5717 4751 5723 4815
rect 5787 4751 5793 4815
rect 5717 3990 5793 4751
rect 5863 4780 5939 4786
rect 5863 4716 5869 4780
rect 5933 4716 5939 4780
rect 6997 4768 7003 4832
rect 7067 4768 7073 4832
rect 6997 4762 7073 4768
rect 7619 6548 7695 6554
rect 7619 6484 7625 6548
rect 7689 6484 7695 6548
rect 7619 4832 7695 6484
rect 8089 6548 8165 8722
rect 8089 6484 8095 6548
rect 8159 6484 8165 6548
rect 8089 6478 8165 6484
rect 7619 4768 7625 4832
rect 7689 4768 7695 4832
rect 5863 4409 5939 4716
rect 5863 4345 5869 4409
rect 5933 4345 5939 4409
rect 5863 4339 5939 4345
rect 5504 3920 5510 3984
rect 5574 3920 5580 3984
rect 5504 3914 5580 3920
rect 5676 3984 5793 3990
rect 5676 3920 5682 3984
rect 5746 3920 5793 3984
rect 5676 3914 5793 3920
rect 5974 3984 6050 3990
rect 5974 3920 5980 3984
rect 6044 3920 6050 3984
rect 4601 3393 4607 3457
rect 4671 3393 4677 3457
rect 4601 2420 4677 3393
rect 4601 2356 4607 2420
rect 4671 2356 4677 2420
rect 4601 2350 4677 2356
rect 5825 3032 5901 3038
rect 5825 2968 5831 3032
rect 5895 2968 5901 3032
rect 5825 1798 5901 2968
rect 5974 3032 6050 3920
rect 5974 2968 5980 3032
rect 6044 2968 6050 3032
rect 5974 2962 6050 2968
rect 5825 1734 5831 1798
rect 5895 1734 5901 1798
rect 5825 1728 5901 1734
rect -800 1631 -794 1695
rect -730 1631 -452 1695
rect -800 -458 -452 1631
rect -800 -522 -794 -458
rect -730 -522 -658 -458
rect -594 -522 -522 -458
rect -458 -522 -452 -458
rect -800 -594 -452 -522
rect -800 -658 -794 -594
rect -730 -658 -658 -594
rect -594 -658 -522 -594
rect -458 -658 -452 -594
rect -800 -730 -452 -658
rect -800 -794 -794 -730
rect -730 -794 -658 -730
rect -594 -794 -522 -730
rect -458 -794 -452 -730
rect -800 -800 -452 -794
rect 4814 1639 4890 1645
rect 4814 1575 4820 1639
rect 4884 1575 4890 1639
rect -1496 -1218 -1490 -1154
rect -1426 -1218 -1354 -1154
rect -1290 -1218 -1218 -1154
rect -1154 -1218 -1148 -1154
rect -1496 -1290 -1148 -1218
rect -1496 -1354 -1490 -1290
rect -1426 -1354 -1354 -1290
rect -1290 -1354 -1218 -1290
rect -1154 -1354 -1148 -1290
rect -1496 -1426 -1148 -1354
rect -1496 -1490 -1490 -1426
rect -1426 -1490 -1354 -1426
rect -1290 -1490 -1218 -1426
rect -1154 -1490 -1148 -1426
rect -1496 -1496 -1148 -1490
rect 4814 -1496 4890 1575
rect 5222 1639 5298 1645
rect 5222 1575 5228 1639
rect 5292 1575 5298 1639
rect 5222 -1496 5298 1575
rect 5630 1639 5706 1645
rect 5630 1575 5636 1639
rect 5700 1575 5706 1639
rect 5630 -1496 5706 1575
rect 7619 -1154 7695 4768
rect 11784 1798 11860 1804
rect 11784 1734 11790 1798
rect 11854 1734 11860 1798
rect 11784 -458 11860 1734
rect 11784 -522 11790 -458
rect 11854 -522 11860 -458
rect 11784 -528 11860 -522
rect 14354 1484 14430 1490
rect 14354 1420 14360 1484
rect 14424 1420 14430 1484
rect 14354 -458 14430 1420
rect 24095 1484 24171 12714
rect 24095 1420 24101 1484
rect 24165 1420 24171 1484
rect 14354 -522 14360 -458
rect 14424 -522 14430 -458
rect 14354 -528 14430 -522
rect 14503 568 14579 574
rect 14503 504 14509 568
rect 14573 504 14579 568
rect 7619 -1218 7625 -1154
rect 7689 -1218 7695 -1154
rect 7619 -1224 7695 -1218
rect 14503 -1154 14579 504
rect 23956 568 24032 574
rect 23956 504 23962 568
rect 24026 504 24032 568
rect 14503 -1218 14509 -1154
rect 14573 -1218 14579 -1154
rect 14503 -1224 14579 -1218
rect 14671 49 14747 55
rect 14671 -15 14677 49
rect 14741 -15 14747 49
rect 14671 -1496 14747 -15
rect 14979 49 15055 55
rect 14979 -15 14985 49
rect 15049 -15 15055 49
rect 14979 -1496 15055 -15
rect 15287 49 15363 55
rect 15287 -15 15293 49
rect 15357 -15 15363 49
rect 15287 -1496 15363 -15
rect 15595 49 15671 55
rect 15595 -15 15601 49
rect 15665 -15 15671 49
rect 15595 -1496 15671 -15
rect 15903 49 15979 55
rect 15903 -15 15909 49
rect 15973 -15 15979 49
rect 15903 -1496 15979 -15
rect 16211 49 16287 55
rect 16211 -15 16217 49
rect 16281 -15 16287 49
rect 16211 -1496 16287 -15
rect 16519 49 16595 55
rect 16519 -15 16525 49
rect 16589 -15 16595 49
rect 16519 -1496 16595 -15
rect 16827 49 16903 55
rect 16827 -15 16833 49
rect 16897 -15 16903 49
rect 16827 -1496 16903 -15
rect 17135 49 17211 55
rect 17135 -15 17141 49
rect 17205 -15 17211 49
rect 17135 -1496 17211 -15
rect 17443 49 17519 55
rect 17443 -15 17449 49
rect 17513 -15 17519 49
rect 17443 -1496 17519 -15
rect 17751 49 17827 55
rect 17751 -15 17757 49
rect 17821 -15 17827 49
rect 17751 -1496 17827 -15
rect 18059 49 18135 55
rect 18059 -15 18065 49
rect 18129 -15 18135 49
rect 18059 -1496 18135 -15
rect 18367 49 18443 55
rect 18367 -15 18373 49
rect 18437 -15 18443 49
rect 18367 -1496 18443 -15
rect 18675 49 18751 55
rect 18675 -15 18681 49
rect 18745 -15 18751 49
rect 18675 -1496 18751 -15
rect 18983 49 19059 55
rect 18983 -15 18989 49
rect 19053 -15 19059 49
rect 18983 -1496 19059 -15
rect 19291 49 19367 55
rect 19291 -15 19297 49
rect 19361 -15 19367 49
rect 19291 -1496 19367 -15
rect 19599 49 19675 55
rect 19599 -15 19605 49
rect 19669 -15 19675 49
rect 19599 -1496 19675 -15
rect 19907 49 19983 55
rect 19907 -15 19913 49
rect 19977 -15 19983 49
rect 19907 -1496 19983 -15
rect 20215 49 20291 55
rect 20215 -15 20221 49
rect 20285 -15 20291 49
rect 20215 -1496 20291 -15
rect 20523 49 20599 55
rect 20523 -15 20529 49
rect 20593 -15 20599 49
rect 20523 -1496 20599 -15
rect 20831 49 20907 55
rect 20831 -15 20837 49
rect 20901 -15 20907 49
rect 20831 -1496 20907 -15
rect 21139 49 21215 55
rect 21139 -15 21145 49
rect 21209 -15 21215 49
rect 21139 -1496 21215 -15
rect 21447 49 21523 55
rect 21447 -15 21453 49
rect 21517 -15 21523 49
rect 21447 -1496 21523 -15
rect 21755 49 21831 55
rect 21755 -15 21761 49
rect 21825 -15 21831 49
rect 21755 -1496 21831 -15
rect 22063 49 22139 55
rect 22063 -15 22069 49
rect 22133 -15 22139 49
rect 22063 -1496 22139 -15
rect 22371 49 22447 55
rect 22371 -15 22377 49
rect 22441 -15 22447 49
rect 22371 -1496 22447 -15
rect 22679 49 22755 55
rect 22679 -15 22685 49
rect 22749 -15 22755 49
rect 22679 -1496 22755 -15
rect 22987 49 23063 55
rect 22987 -15 22993 49
rect 23057 -15 23063 49
rect 22987 -1496 23063 -15
rect 23295 49 23371 55
rect 23295 -15 23301 49
rect 23365 -15 23371 49
rect 23295 -1496 23371 -15
rect 23603 49 23679 55
rect 23603 -15 23609 49
rect 23673 -15 23679 49
rect 23603 -1496 23679 -15
rect 23762 49 23838 55
rect 23762 -15 23768 49
rect 23832 -15 23838 49
rect 23762 -1496 23838 -15
rect 23956 -1154 24032 504
rect 24095 -458 24171 1420
rect 24095 -522 24101 -458
rect 24165 -522 24171 -458
rect 24095 -528 24171 -522
rect 24339 568 24415 13410
rect 49136 13474 49212 13480
rect 49136 13410 49142 13474
rect 49206 13410 49212 13474
rect 34328 12778 34404 12784
rect 34328 12714 34334 12778
rect 34398 12714 34404 12778
rect 34328 10315 34404 12714
rect 34328 10251 34334 10315
rect 34398 10251 34404 10315
rect 34328 7374 34404 10251
rect 36407 12778 36483 12784
rect 36407 12714 36413 12778
rect 36477 12714 36483 12778
rect 36407 10315 36483 12714
rect 36407 10251 36413 10315
rect 36477 10251 36483 10315
rect 36407 10245 36483 10251
rect 48718 12778 48794 12784
rect 48718 12714 48724 12778
rect 48788 12714 48794 12778
rect 48718 10315 48794 12714
rect 48718 10251 48724 10315
rect 48788 10251 48794 10315
rect 48718 10245 48794 10251
rect 49136 8786 49212 13410
rect 60313 13474 60389 13480
rect 60313 13410 60319 13474
rect 60383 13410 60389 13474
rect 60094 12778 60170 12784
rect 60094 12714 60100 12778
rect 60164 12714 60170 12778
rect 60094 12228 60170 12714
rect 60094 12164 60100 12228
rect 60164 12164 60170 12228
rect 60094 12158 60170 12164
rect 49136 8722 49142 8786
rect 49206 8722 49212 8786
rect 48718 7870 48794 7876
rect 48718 7806 48724 7870
rect 48788 7806 48794 7870
rect 34260 7368 34404 7374
rect 34260 7304 34266 7368
rect 34330 7304 34404 7368
rect 34260 7298 34404 7304
rect 36407 7368 36483 7374
rect 36407 7304 36413 7368
rect 36477 7304 36483 7368
rect 24339 504 24345 568
rect 24409 504 24415 568
rect 23956 -1218 23962 -1154
rect 24026 -1218 24032 -1154
rect 23956 -1224 24032 -1218
rect 24339 -1154 24415 504
rect 24339 -1218 24345 -1154
rect 24409 -1218 24415 -1154
rect 24339 -1224 24415 -1218
rect 24477 49 24553 55
rect 24477 -15 24483 49
rect 24547 -15 24553 49
rect 24477 -1496 24553 -15
rect 36407 -458 36483 7304
rect 36407 -522 36413 -458
rect 36477 -522 36483 -458
rect 36407 -528 36483 -522
rect 36546 568 36622 574
rect 36546 504 36552 568
rect 36616 504 36622 568
rect 36546 -1154 36622 504
rect 48718 -458 48794 7806
rect 48718 -522 48724 -458
rect 48788 -522 48794 -458
rect 48718 -528 48794 -522
rect 36546 -1218 36552 -1154
rect 36616 -1218 36622 -1154
rect 36546 -1224 36622 -1218
rect 49136 -1154 49212 8722
rect 60313 8786 60389 13410
rect 61726 13474 62074 13546
rect 61726 13410 61732 13474
rect 61796 13410 61868 13474
rect 61932 13410 62004 13474
rect 62068 13410 62074 13474
rect 60313 8722 60319 8786
rect 60383 8722 60389 8786
rect 60313 8716 60389 8722
rect 61030 13050 61378 13056
rect 61030 12986 61036 13050
rect 61100 12986 61172 13050
rect 61236 12986 61308 13050
rect 61372 12986 61378 13050
rect 61030 12914 61378 12986
rect 61030 12850 61036 12914
rect 61100 12850 61172 12914
rect 61236 12850 61308 12914
rect 61372 12850 61378 12914
rect 61030 12778 61378 12850
rect 61030 12714 61036 12778
rect 61100 12714 61172 12778
rect 61236 12714 61308 12778
rect 61372 12714 61378 12778
rect 61030 12228 61378 12714
rect 61030 12164 61036 12228
rect 61100 12164 61378 12228
rect 61030 7870 61378 12164
rect 61030 7806 61036 7870
rect 61100 7806 61378 7870
rect 61030 -458 61378 7806
rect 61030 -522 61036 -458
rect 61100 -522 61172 -458
rect 61236 -522 61308 -458
rect 61372 -522 61378 -458
rect 61030 -594 61378 -522
rect 61030 -658 61036 -594
rect 61100 -658 61172 -594
rect 61236 -658 61308 -594
rect 61372 -658 61378 -594
rect 61030 -730 61378 -658
rect 61030 -794 61036 -730
rect 61100 -794 61172 -730
rect 61236 -794 61308 -730
rect 61372 -794 61378 -730
rect 61030 -800 61378 -794
rect 61726 8786 62074 13410
rect 61726 8722 61732 8786
rect 61796 8722 62074 8786
rect 49136 -1218 49142 -1154
rect 49206 -1218 49212 -1154
rect 49136 -1224 49212 -1218
rect 61726 -1154 62074 8722
rect 61726 -1218 61732 -1154
rect 61796 -1218 61868 -1154
rect 61932 -1218 62004 -1154
rect 62068 -1218 62074 -1154
rect 61726 -1290 62074 -1218
rect 61726 -1354 61732 -1290
rect 61796 -1354 61868 -1290
rect 61932 -1354 62004 -1290
rect 62068 -1354 62074 -1290
rect 61726 -1426 62074 -1354
rect 61726 -1490 61732 -1426
rect 61796 -1490 61868 -1426
rect 61932 -1490 62004 -1426
rect 62068 -1490 62074 -1426
rect 61726 -1496 62074 -1490
use sky130_rom_krom_rom_base_array  sky130_rom_krom_rom_base_array_0
timestamp 1581365160
transform 1 0 8105 0 1 9410
box 0 -84 52473 2813
use sky130_rom_krom_rom_bitline_inverter  sky130_rom_krom_rom_bitline_inverter_0
timestamp 1581365163
transform 0 -1 60351 1 0 7508
box 136 -79 1879 52319
use sky130_rom_krom_rom_column_decode  sky130_rom_krom_rom_column_decode_0
timestamp 1581365163
transform 1 0 4498 0 1 1530
box -39 44 3513 5257
use sky130_rom_krom_rom_column_mux_array  sky130_rom_krom_rom_column_mux_array_0
timestamp 1581365163
transform 1 0 8153 0 1 4342
box 0 382 52275 3061
use sky130_rom_krom_rom_control_logic  sky130_rom_krom_rom_control_logic_0
timestamp 1581365163
transform 1 0 -1450 0 1 1663
box -36 -49 5744 5306
use sky130_rom_krom_rom_output_buffer  sky130_rom_krom_rom_output_buffer_0
timestamp 1581365163
transform 0 1 14521 -1 0 1782
box 44 -50 1800 9951
use sky130_rom_krom_rom_row_decode  sky130_rom_krom_rom_row_decode_0
timestamp 1581365162
transform 1 0 0 0 1 6999
box -39 44 8011 5257
<< labels >>
rlabel metal3 s -1496 1895 -1420 1971 4 cs0
port 3 nsew
rlabel metal3 s -1496 2902 -1420 2978 4 clk0
port 5 nsew
rlabel metal4 s 14671 -1496 14747 -1420 4 dout0[0]
port 7 nsew
rlabel metal4 s 14979 -1496 15055 -1420 4 dout0[1]
port 9 nsew
rlabel metal4 s 15287 -1496 15363 -1420 4 dout0[2]
port 11 nsew
rlabel metal4 s 15595 -1496 15671 -1420 4 dout0[3]
port 13 nsew
rlabel metal4 s 15903 -1496 15979 -1420 4 dout0[4]
port 15 nsew
rlabel metal4 s 16211 -1496 16287 -1420 4 dout0[5]
port 17 nsew
rlabel metal4 s 16519 -1496 16595 -1420 4 dout0[6]
port 19 nsew
rlabel metal4 s 16827 -1496 16903 -1420 4 dout0[7]
port 21 nsew
rlabel metal4 s 17135 -1496 17211 -1420 4 dout0[8]
port 23 nsew
rlabel metal4 s 17443 -1496 17519 -1420 4 dout0[9]
port 25 nsew
rlabel metal4 s 17751 -1496 17827 -1420 4 dout0[10]
port 27 nsew
rlabel metal4 s 18059 -1496 18135 -1420 4 dout0[11]
port 29 nsew
rlabel metal4 s 18367 -1496 18443 -1420 4 dout0[12]
port 31 nsew
rlabel metal4 s 18675 -1496 18751 -1420 4 dout0[13]
port 33 nsew
rlabel metal4 s 18983 -1496 19059 -1420 4 dout0[14]
port 35 nsew
rlabel metal4 s 19291 -1496 19367 -1420 4 dout0[15]
port 37 nsew
rlabel metal4 s 19599 -1496 19675 -1420 4 dout0[16]
port 39 nsew
rlabel metal4 s 19907 -1496 19983 -1420 4 dout0[17]
port 41 nsew
rlabel metal4 s 20215 -1496 20291 -1420 4 dout0[18]
port 43 nsew
rlabel metal4 s 20523 -1496 20599 -1420 4 dout0[19]
port 45 nsew
rlabel metal4 s 20831 -1496 20907 -1420 4 dout0[20]
port 47 nsew
rlabel metal4 s 21139 -1496 21215 -1420 4 dout0[21]
port 49 nsew
rlabel metal4 s 21447 -1496 21523 -1420 4 dout0[22]
port 51 nsew
rlabel metal4 s 21755 -1496 21831 -1420 4 dout0[23]
port 53 nsew
rlabel metal4 s 22063 -1496 22139 -1420 4 dout0[24]
port 55 nsew
rlabel metal4 s 22371 -1496 22447 -1420 4 dout0[25]
port 57 nsew
rlabel metal4 s 22679 -1496 22755 -1420 4 dout0[26]
port 59 nsew
rlabel metal4 s 22987 -1496 23063 -1420 4 dout0[27]
port 61 nsew
rlabel metal4 s 23295 -1496 23371 -1420 4 dout0[28]
port 63 nsew
rlabel metal4 s 23603 -1496 23679 -1420 4 dout0[29]
port 65 nsew
rlabel metal4 s 23762 -1496 23838 -1420 4 dout0[30]
port 67 nsew
rlabel metal4 s 24477 -1496 24553 -1420 4 dout0[31]
port 69 nsew
rlabel metal4 s 4814 -1496 4890 -1420 4 addr0[0]
port 71 nsew
rlabel metal4 s 5222 -1496 5298 -1420 4 addr0[1]
port 73 nsew
rlabel metal4 s 5630 -1496 5706 -1420 4 addr0[2]
port 75 nsew
rlabel metal3 s -1496 7038 -1420 7114 4 addr0[3]
port 77 nsew
rlabel metal3 s -1496 6744 -1420 6820 4 addr0[4]
port 79 nsew
rlabel metal3 s -1496 7335 -1420 7411 4 addr0[5]
port 81 nsew
rlabel metal3 s -1496 13404 62074 13752 4 vccd1
port 83 nsew
rlabel metal3 s -1496 -1496 62074 -1148 4 vccd1
port 83 nsew
rlabel metal4 s 61726 -1496 62074 13752 4 vccd1
port 83 nsew
rlabel metal4 s -1496 -1496 -1148 13752 4 vccd1
port 83 nsew
rlabel metal3 s -800 -800 61378 -452 4 vssd1
port 85 nsew
rlabel metal3 s -800 12708 61378 13056 4 vssd1
port 85 nsew
rlabel metal4 s -800 -800 -452 13056 4 vssd1
port 85 nsew
rlabel metal4 s 61030 -800 61378 13056 4 vssd1
port 85 nsew
<< properties >>
string FIXED_BBOX 61998 -1491 62074 -1425
<< end >>
