magic
tech sky130A
magscale 1 2
timestamp 1581365163
<< checkpaint >>
rect -1296 -1277 1772 3946
<< nwell >>
rect -36 1262 512 2686
<< pwell >>
rect 28 159 338 225
rect 28 25 442 159
<< scnmos >>
rect 114 51 144 199
rect 222 51 252 199
<< scpmos >>
rect 114 2326 144 2578
rect 222 2326 252 2578
<< ndiff >>
rect 54 142 114 199
rect 54 108 62 142
rect 96 108 114 142
rect 54 51 114 108
rect 144 142 222 199
rect 144 108 166 142
rect 200 108 222 142
rect 144 51 222 108
rect 252 142 312 199
rect 252 108 270 142
rect 304 108 312 142
rect 252 51 312 108
<< pdiff >>
rect 54 2469 114 2578
rect 54 2435 62 2469
rect 96 2435 114 2469
rect 54 2326 114 2435
rect 144 2469 222 2578
rect 144 2435 166 2469
rect 200 2435 222 2469
rect 144 2326 222 2435
rect 252 2469 312 2578
rect 252 2435 270 2469
rect 304 2435 312 2469
rect 252 2326 312 2435
<< ndiffc >>
rect 62 108 96 142
rect 166 108 200 142
rect 270 108 304 142
<< pdiffc >>
rect 62 2435 96 2469
rect 166 2435 200 2469
rect 270 2435 304 2469
<< psubdiff >>
rect 366 109 416 133
rect 366 75 374 109
rect 408 75 416 109
rect 366 51 416 75
<< nsubdiff >>
rect 366 2541 416 2565
rect 366 2507 374 2541
rect 408 2507 416 2541
rect 366 2483 416 2507
<< psubdiffcont >>
rect 374 75 408 109
<< nsubdiffcont >>
rect 374 2507 408 2541
<< poly >>
rect 114 2578 144 2604
rect 222 2578 252 2604
rect 114 2300 144 2326
rect 222 2300 252 2326
rect 114 2270 252 2300
rect 114 1322 144 2270
rect 48 1306 144 1322
rect 48 1272 64 1306
rect 98 1272 144 1306
rect 48 1256 144 1272
rect 114 255 144 1256
rect 114 225 252 255
rect 114 199 144 225
rect 222 199 252 225
rect 114 25 144 51
rect 222 25 252 51
<< polycont >>
rect 64 1272 98 1306
<< locali >>
rect 0 2612 476 2646
rect 62 2469 96 2612
rect 62 2419 96 2435
rect 166 2469 200 2485
rect 64 1306 98 1322
rect 64 1256 98 1272
rect 166 1306 200 2435
rect 270 2469 304 2612
rect 374 2541 408 2612
rect 374 2491 408 2507
rect 270 2419 304 2435
rect 166 1272 217 1306
rect 62 142 96 158
rect 62 17 96 108
rect 166 142 200 1272
rect 166 92 200 108
rect 270 142 304 158
rect 270 17 304 108
rect 374 109 408 125
rect 374 17 408 75
rect 0 -17 476 17
<< labels >>
rlabel locali s 81 1289 81 1289 4 A
port 1 nsew
rlabel locali s 200 1289 200 1289 4 Z
port 2 nsew
rlabel locali s 238 0 238 0 4 gnd
port 3 nsew
rlabel locali s 238 2629 238 2629 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 476 2368
<< end >>
