magic
tech sky130A
magscale 1 2
timestamp 1581479693
<< checkpaint >>
rect -1296 -1277 1880 3946
<< nwell >>
rect -36 1262 620 2686
<< pwell >>
rect 28 159 446 677
rect 28 25 550 159
<< scnmos >>
rect 114 51 144 651
rect 222 51 252 651
rect 330 51 360 651
<< scpmos >>
rect 114 1978 144 2578
rect 222 1978 252 2578
rect 330 1978 360 2578
<< ndiff >>
rect 54 368 114 651
rect 54 334 62 368
rect 96 334 114 368
rect 54 51 114 334
rect 144 368 222 651
rect 144 334 166 368
rect 200 334 222 368
rect 144 51 222 334
rect 252 368 330 651
rect 252 334 274 368
rect 308 334 330 368
rect 252 51 330 334
rect 360 368 420 651
rect 360 334 378 368
rect 412 334 420 368
rect 360 51 420 334
<< pdiff >>
rect 54 2295 114 2578
rect 54 2261 62 2295
rect 96 2261 114 2295
rect 54 1978 114 2261
rect 144 2295 222 2578
rect 144 2261 166 2295
rect 200 2261 222 2295
rect 144 1978 222 2261
rect 252 2295 330 2578
rect 252 2261 274 2295
rect 308 2261 330 2295
rect 252 1978 330 2261
rect 360 2295 420 2578
rect 360 2261 378 2295
rect 412 2261 420 2295
rect 360 1978 420 2261
<< ndiffc >>
rect 62 334 96 368
rect 166 334 200 368
rect 274 334 308 368
rect 378 334 412 368
<< pdiffc >>
rect 62 2261 96 2295
rect 166 2261 200 2295
rect 274 2261 308 2295
rect 378 2261 412 2295
<< psubdiff >>
rect 474 109 524 133
rect 474 75 482 109
rect 516 75 524 109
rect 474 51 524 75
<< nsubdiff >>
rect 474 2541 524 2565
rect 474 2507 482 2541
rect 516 2507 524 2541
rect 474 2483 524 2507
<< psubdiffcont >>
rect 482 75 516 109
<< nsubdiffcont >>
rect 482 2507 516 2541
<< poly >>
rect 114 2578 144 2604
rect 222 2578 252 2604
rect 330 2578 360 2604
rect 114 1952 144 1978
rect 222 1952 252 1978
rect 330 1952 360 1978
rect 114 1922 360 1952
rect 114 1348 144 1922
rect 48 1332 144 1348
rect 48 1298 64 1332
rect 98 1298 144 1332
rect 48 1282 144 1298
rect 114 707 144 1282
rect 114 677 360 707
rect 114 651 144 677
rect 222 651 252 677
rect 330 651 360 677
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
<< polycont >>
rect 64 1298 98 1332
<< locali >>
rect 0 2612 584 2646
rect 62 2295 96 2612
rect 62 2245 96 2261
rect 166 2295 200 2311
rect 166 2211 200 2261
rect 274 2295 308 2612
rect 482 2541 516 2612
rect 482 2491 516 2507
rect 274 2245 308 2261
rect 378 2295 412 2311
rect 378 2211 412 2261
rect 166 2177 412 2211
rect 64 1332 98 1348
rect 64 1282 98 1298
rect 272 1332 306 2177
rect 272 1298 323 1332
rect 272 452 306 1298
rect 166 418 412 452
rect 62 368 96 384
rect 62 17 96 334
rect 166 368 200 418
rect 166 318 200 334
rect 274 368 308 384
rect 274 17 308 334
rect 378 368 412 418
rect 378 318 412 334
rect 482 109 516 125
rect 482 17 516 75
rect 0 -17 584 17
<< labels >>
rlabel locali s 81 1315 81 1315 4 A
port 1 nsew
rlabel locali s 306 1315 306 1315 4 Z
port 2 nsew
rlabel locali s 292 0 292 0 4 gnd
port 3 nsew
rlabel locali s 292 2629 292 2629 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 584 2194
<< end >>
