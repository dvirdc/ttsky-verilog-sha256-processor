magic
tech sky130A
magscale 1 2
timestamp 1581449086
<< checkpaint >>
rect -1260 -1260 1261 1261
<< end >>
