magic
tech sky130A
magscale 1 2
timestamp 1581449086
<< checkpaint >>
rect -1260 -1472 53592 1668
<< nwell >>
rect 0 -196 52332 408
<< poly >>
rect 60 65 90 240
rect 1692 65 1722 240
rect 3324 65 3354 240
rect 4956 65 4986 240
rect 6588 65 6618 240
rect 8220 65 8250 240
rect 9852 65 9882 240
rect 11484 65 11514 240
rect 13116 65 13146 240
rect 14748 65 14778 240
rect 16380 65 16410 240
rect 18012 65 18042 240
rect 19644 65 19674 240
rect 21276 65 21306 240
rect 22908 65 22938 240
rect 24540 65 24570 240
rect 26172 65 26202 240
rect 27804 65 27834 240
rect 29436 65 29466 240
rect 31068 65 31098 240
rect 32700 65 32730 240
rect 34332 65 34362 240
rect 35964 65 35994 240
rect 37596 65 37626 240
rect 39228 65 39258 240
rect 40860 65 40890 240
rect 42492 65 42522 240
rect 44124 65 44154 240
rect 45756 65 45786 240
rect 47388 65 47418 240
rect 49020 65 49050 240
rect 50652 65 50682 240
rect 52284 65 52314 240
rect 60 50 52314 65
rect 61 35 52314 50
<< locali >>
rect 35 -111 69 -95
rect 35 -161 69 -145
rect 239 -111 273 -95
rect 239 -161 273 -145
rect 443 -111 477 -95
rect 443 -161 477 -145
rect 647 -111 681 -95
rect 647 -161 681 -145
rect 851 -111 885 -95
rect 851 -161 885 -145
rect 1055 -111 1089 -95
rect 1055 -161 1089 -145
rect 1259 -111 1293 -95
rect 1259 -161 1293 -145
rect 1463 -111 1497 -95
rect 1463 -161 1497 -145
rect 1667 -111 1701 -95
rect 1667 -161 1701 -145
rect 1871 -111 1905 -95
rect 1871 -161 1905 -145
rect 2075 -111 2109 -95
rect 2075 -161 2109 -145
rect 2279 -111 2313 -95
rect 2279 -161 2313 -145
rect 2483 -111 2517 -95
rect 2483 -161 2517 -145
rect 2687 -111 2721 -95
rect 2687 -161 2721 -145
rect 2891 -111 2925 -95
rect 2891 -161 2925 -145
rect 3095 -111 3129 -95
rect 3095 -161 3129 -145
rect 3299 -111 3333 -95
rect 3299 -161 3333 -145
rect 3503 -111 3537 -95
rect 3503 -161 3537 -145
rect 3707 -111 3741 -95
rect 3707 -161 3741 -145
rect 3911 -111 3945 -95
rect 3911 -161 3945 -145
rect 4115 -111 4149 -95
rect 4115 -161 4149 -145
rect 4319 -111 4353 -95
rect 4319 -161 4353 -145
rect 4523 -111 4557 -95
rect 4523 -161 4557 -145
rect 4727 -111 4761 -95
rect 4727 -161 4761 -145
rect 4931 -111 4965 -95
rect 4931 -161 4965 -145
rect 5135 -111 5169 -95
rect 5135 -161 5169 -145
rect 5339 -111 5373 -95
rect 5339 -161 5373 -145
rect 5543 -111 5577 -95
rect 5543 -161 5577 -145
rect 5747 -111 5781 -95
rect 5747 -161 5781 -145
rect 5951 -111 5985 -95
rect 5951 -161 5985 -145
rect 6155 -111 6189 -95
rect 6155 -161 6189 -145
rect 6359 -111 6393 -95
rect 6359 -161 6393 -145
rect 6563 -111 6597 -95
rect 6563 -161 6597 -145
rect 6767 -111 6801 -95
rect 6767 -161 6801 -145
rect 6971 -111 7005 -95
rect 6971 -161 7005 -145
rect 7175 -111 7209 -95
rect 7175 -161 7209 -145
rect 7379 -111 7413 -95
rect 7379 -161 7413 -145
rect 7583 -111 7617 -95
rect 7583 -161 7617 -145
rect 7787 -111 7821 -95
rect 7787 -161 7821 -145
rect 7991 -111 8025 -95
rect 7991 -161 8025 -145
rect 8195 -111 8229 -95
rect 8195 -161 8229 -145
rect 8399 -111 8433 -95
rect 8399 -161 8433 -145
rect 8603 -111 8637 -95
rect 8603 -161 8637 -145
rect 8807 -111 8841 -95
rect 8807 -161 8841 -145
rect 9011 -111 9045 -95
rect 9011 -161 9045 -145
rect 9215 -111 9249 -95
rect 9215 -161 9249 -145
rect 9419 -111 9453 -95
rect 9419 -161 9453 -145
rect 9623 -111 9657 -95
rect 9623 -161 9657 -145
rect 9827 -111 9861 -95
rect 9827 -161 9861 -145
rect 10031 -111 10065 -95
rect 10031 -161 10065 -145
rect 10235 -111 10269 -95
rect 10235 -161 10269 -145
rect 10439 -111 10473 -95
rect 10439 -161 10473 -145
rect 10643 -111 10677 -95
rect 10643 -161 10677 -145
rect 10847 -111 10881 -95
rect 10847 -161 10881 -145
rect 11051 -111 11085 -95
rect 11051 -161 11085 -145
rect 11255 -111 11289 -95
rect 11255 -161 11289 -145
rect 11459 -111 11493 -95
rect 11459 -161 11493 -145
rect 11663 -111 11697 -95
rect 11663 -161 11697 -145
rect 11867 -111 11901 -95
rect 11867 -161 11901 -145
rect 12071 -111 12105 -95
rect 12071 -161 12105 -145
rect 12275 -111 12309 -95
rect 12275 -161 12309 -145
rect 12479 -111 12513 -95
rect 12479 -161 12513 -145
rect 12683 -111 12717 -95
rect 12683 -161 12717 -145
rect 12887 -111 12921 -95
rect 12887 -161 12921 -145
rect 13091 -111 13125 -95
rect 13091 -161 13125 -145
rect 13295 -111 13329 -95
rect 13295 -161 13329 -145
rect 13499 -111 13533 -95
rect 13499 -161 13533 -145
rect 13703 -111 13737 -95
rect 13703 -161 13737 -145
rect 13907 -111 13941 -95
rect 13907 -161 13941 -145
rect 14111 -111 14145 -95
rect 14111 -161 14145 -145
rect 14315 -111 14349 -95
rect 14315 -161 14349 -145
rect 14519 -111 14553 -95
rect 14519 -161 14553 -145
rect 14723 -111 14757 -95
rect 14723 -161 14757 -145
rect 14927 -111 14961 -95
rect 14927 -161 14961 -145
rect 15131 -111 15165 -95
rect 15131 -161 15165 -145
rect 15335 -111 15369 -95
rect 15335 -161 15369 -145
rect 15539 -111 15573 -95
rect 15539 -161 15573 -145
rect 15743 -111 15777 -95
rect 15743 -161 15777 -145
rect 15947 -111 15981 -95
rect 15947 -161 15981 -145
rect 16151 -111 16185 -95
rect 16151 -161 16185 -145
rect 16355 -111 16389 -95
rect 16355 -161 16389 -145
rect 16559 -111 16593 -95
rect 16559 -161 16593 -145
rect 16763 -111 16797 -95
rect 16763 -161 16797 -145
rect 16967 -111 17001 -95
rect 16967 -161 17001 -145
rect 17171 -111 17205 -95
rect 17171 -161 17205 -145
rect 17375 -111 17409 -95
rect 17375 -161 17409 -145
rect 17579 -111 17613 -95
rect 17579 -161 17613 -145
rect 17783 -111 17817 -95
rect 17783 -161 17817 -145
rect 17987 -111 18021 -95
rect 17987 -161 18021 -145
rect 18191 -111 18225 -95
rect 18191 -161 18225 -145
rect 18395 -111 18429 -95
rect 18395 -161 18429 -145
rect 18599 -111 18633 -95
rect 18599 -161 18633 -145
rect 18803 -111 18837 -95
rect 18803 -161 18837 -145
rect 19007 -111 19041 -95
rect 19007 -161 19041 -145
rect 19211 -111 19245 -95
rect 19211 -161 19245 -145
rect 19415 -111 19449 -95
rect 19415 -161 19449 -145
rect 19619 -111 19653 -95
rect 19619 -161 19653 -145
rect 19823 -111 19857 -95
rect 19823 -161 19857 -145
rect 20027 -111 20061 -95
rect 20027 -161 20061 -145
rect 20231 -111 20265 -95
rect 20231 -161 20265 -145
rect 20435 -111 20469 -95
rect 20435 -161 20469 -145
rect 20639 -111 20673 -95
rect 20639 -161 20673 -145
rect 20843 -111 20877 -95
rect 20843 -161 20877 -145
rect 21047 -111 21081 -95
rect 21047 -161 21081 -145
rect 21251 -111 21285 -95
rect 21251 -161 21285 -145
rect 21455 -111 21489 -95
rect 21455 -161 21489 -145
rect 21659 -111 21693 -95
rect 21659 -161 21693 -145
rect 21863 -111 21897 -95
rect 21863 -161 21897 -145
rect 22067 -111 22101 -95
rect 22067 -161 22101 -145
rect 22271 -111 22305 -95
rect 22271 -161 22305 -145
rect 22475 -111 22509 -95
rect 22475 -161 22509 -145
rect 22679 -111 22713 -95
rect 22679 -161 22713 -145
rect 22883 -111 22917 -95
rect 22883 -161 22917 -145
rect 23087 -111 23121 -95
rect 23087 -161 23121 -145
rect 23291 -111 23325 -95
rect 23291 -161 23325 -145
rect 23495 -111 23529 -95
rect 23495 -161 23529 -145
rect 23699 -111 23733 -95
rect 23699 -161 23733 -145
rect 23903 -111 23937 -95
rect 23903 -161 23937 -145
rect 24107 -111 24141 -95
rect 24107 -161 24141 -145
rect 24311 -111 24345 -95
rect 24311 -161 24345 -145
rect 24515 -111 24549 -95
rect 24515 -161 24549 -145
rect 24719 -111 24753 -95
rect 24719 -161 24753 -145
rect 24923 -111 24957 -95
rect 24923 -161 24957 -145
rect 25127 -111 25161 -95
rect 25127 -161 25161 -145
rect 25331 -111 25365 -95
rect 25331 -161 25365 -145
rect 25535 -111 25569 -95
rect 25535 -161 25569 -145
rect 25739 -111 25773 -95
rect 25739 -161 25773 -145
rect 25943 -111 25977 -95
rect 25943 -161 25977 -145
rect 26147 -111 26181 -95
rect 26147 -161 26181 -145
rect 26351 -111 26385 -95
rect 26351 -161 26385 -145
rect 26555 -111 26589 -95
rect 26555 -161 26589 -145
rect 26759 -111 26793 -95
rect 26759 -161 26793 -145
rect 26963 -111 26997 -95
rect 26963 -161 26997 -145
rect 27167 -111 27201 -95
rect 27167 -161 27201 -145
rect 27371 -111 27405 -95
rect 27371 -161 27405 -145
rect 27575 -111 27609 -95
rect 27575 -161 27609 -145
rect 27779 -111 27813 -95
rect 27779 -161 27813 -145
rect 27983 -111 28017 -95
rect 27983 -161 28017 -145
rect 28187 -111 28221 -95
rect 28187 -161 28221 -145
rect 28391 -111 28425 -95
rect 28391 -161 28425 -145
rect 28595 -111 28629 -95
rect 28595 -161 28629 -145
rect 28799 -111 28833 -95
rect 28799 -161 28833 -145
rect 29003 -111 29037 -95
rect 29003 -161 29037 -145
rect 29207 -111 29241 -95
rect 29207 -161 29241 -145
rect 29411 -111 29445 -95
rect 29411 -161 29445 -145
rect 29615 -111 29649 -95
rect 29615 -161 29649 -145
rect 29819 -111 29853 -95
rect 29819 -161 29853 -145
rect 30023 -111 30057 -95
rect 30023 -161 30057 -145
rect 30227 -111 30261 -95
rect 30227 -161 30261 -145
rect 30431 -111 30465 -95
rect 30431 -161 30465 -145
rect 30635 -111 30669 -95
rect 30635 -161 30669 -145
rect 30839 -111 30873 -95
rect 30839 -161 30873 -145
rect 31043 -111 31077 -95
rect 31043 -161 31077 -145
rect 31247 -111 31281 -95
rect 31247 -161 31281 -145
rect 31451 -111 31485 -95
rect 31451 -161 31485 -145
rect 31655 -111 31689 -95
rect 31655 -161 31689 -145
rect 31859 -111 31893 -95
rect 31859 -161 31893 -145
rect 32063 -111 32097 -95
rect 32063 -161 32097 -145
rect 32267 -111 32301 -95
rect 32267 -161 32301 -145
rect 32471 -111 32505 -95
rect 32471 -161 32505 -145
rect 32675 -111 32709 -95
rect 32675 -161 32709 -145
rect 32879 -111 32913 -95
rect 32879 -161 32913 -145
rect 33083 -111 33117 -95
rect 33083 -161 33117 -145
rect 33287 -111 33321 -95
rect 33287 -161 33321 -145
rect 33491 -111 33525 -95
rect 33491 -161 33525 -145
rect 33695 -111 33729 -95
rect 33695 -161 33729 -145
rect 33899 -111 33933 -95
rect 33899 -161 33933 -145
rect 34103 -111 34137 -95
rect 34103 -161 34137 -145
rect 34307 -111 34341 -95
rect 34307 -161 34341 -145
rect 34511 -111 34545 -95
rect 34511 -161 34545 -145
rect 34715 -111 34749 -95
rect 34715 -161 34749 -145
rect 34919 -111 34953 -95
rect 34919 -161 34953 -145
rect 35123 -111 35157 -95
rect 35123 -161 35157 -145
rect 35327 -111 35361 -95
rect 35327 -161 35361 -145
rect 35531 -111 35565 -95
rect 35531 -161 35565 -145
rect 35735 -111 35769 -95
rect 35735 -161 35769 -145
rect 35939 -111 35973 -95
rect 35939 -161 35973 -145
rect 36143 -111 36177 -95
rect 36143 -161 36177 -145
rect 36347 -111 36381 -95
rect 36347 -161 36381 -145
rect 36551 -111 36585 -95
rect 36551 -161 36585 -145
rect 36755 -111 36789 -95
rect 36755 -161 36789 -145
rect 36959 -111 36993 -95
rect 36959 -161 36993 -145
rect 37163 -111 37197 -95
rect 37163 -161 37197 -145
rect 37367 -111 37401 -95
rect 37367 -161 37401 -145
rect 37571 -111 37605 -95
rect 37571 -161 37605 -145
rect 37775 -111 37809 -95
rect 37775 -161 37809 -145
rect 37979 -111 38013 -95
rect 37979 -161 38013 -145
rect 38183 -111 38217 -95
rect 38183 -161 38217 -145
rect 38387 -111 38421 -95
rect 38387 -161 38421 -145
rect 38591 -111 38625 -95
rect 38591 -161 38625 -145
rect 38795 -111 38829 -95
rect 38795 -161 38829 -145
rect 38999 -111 39033 -95
rect 38999 -161 39033 -145
rect 39203 -111 39237 -95
rect 39203 -161 39237 -145
rect 39407 -111 39441 -95
rect 39407 -161 39441 -145
rect 39611 -111 39645 -95
rect 39611 -161 39645 -145
rect 39815 -111 39849 -95
rect 39815 -161 39849 -145
rect 40019 -111 40053 -95
rect 40019 -161 40053 -145
rect 40223 -111 40257 -95
rect 40223 -161 40257 -145
rect 40427 -111 40461 -95
rect 40427 -161 40461 -145
rect 40631 -111 40665 -95
rect 40631 -161 40665 -145
rect 40835 -111 40869 -95
rect 40835 -161 40869 -145
rect 41039 -111 41073 -95
rect 41039 -161 41073 -145
rect 41243 -111 41277 -95
rect 41243 -161 41277 -145
rect 41447 -111 41481 -95
rect 41447 -161 41481 -145
rect 41651 -111 41685 -95
rect 41651 -161 41685 -145
rect 41855 -111 41889 -95
rect 41855 -161 41889 -145
rect 42059 -111 42093 -95
rect 42059 -161 42093 -145
rect 42263 -111 42297 -95
rect 42263 -161 42297 -145
rect 42467 -111 42501 -95
rect 42467 -161 42501 -145
rect 42671 -111 42705 -95
rect 42671 -161 42705 -145
rect 42875 -111 42909 -95
rect 42875 -161 42909 -145
rect 43079 -111 43113 -95
rect 43079 -161 43113 -145
rect 43283 -111 43317 -95
rect 43283 -161 43317 -145
rect 43487 -111 43521 -95
rect 43487 -161 43521 -145
rect 43691 -111 43725 -95
rect 43691 -161 43725 -145
rect 43895 -111 43929 -95
rect 43895 -161 43929 -145
rect 44099 -111 44133 -95
rect 44099 -161 44133 -145
rect 44303 -111 44337 -95
rect 44303 -161 44337 -145
rect 44507 -111 44541 -95
rect 44507 -161 44541 -145
rect 44711 -111 44745 -95
rect 44711 -161 44745 -145
rect 44915 -111 44949 -95
rect 44915 -161 44949 -145
rect 45119 -111 45153 -95
rect 45119 -161 45153 -145
rect 45323 -111 45357 -95
rect 45323 -161 45357 -145
rect 45527 -111 45561 -95
rect 45527 -161 45561 -145
rect 45731 -111 45765 -95
rect 45731 -161 45765 -145
rect 45935 -111 45969 -95
rect 45935 -161 45969 -145
rect 46139 -111 46173 -95
rect 46139 -161 46173 -145
rect 46343 -111 46377 -95
rect 46343 -161 46377 -145
rect 46547 -111 46581 -95
rect 46547 -161 46581 -145
rect 46751 -111 46785 -95
rect 46751 -161 46785 -145
rect 46955 -111 46989 -95
rect 46955 -161 46989 -145
rect 47159 -111 47193 -95
rect 47159 -161 47193 -145
rect 47363 -111 47397 -95
rect 47363 -161 47397 -145
rect 47567 -111 47601 -95
rect 47567 -161 47601 -145
rect 47771 -111 47805 -95
rect 47771 -161 47805 -145
rect 47975 -111 48009 -95
rect 47975 -161 48009 -145
rect 48179 -111 48213 -95
rect 48179 -161 48213 -145
rect 48383 -111 48417 -95
rect 48383 -161 48417 -145
rect 48587 -111 48621 -95
rect 48587 -161 48621 -145
rect 48791 -111 48825 -95
rect 48791 -161 48825 -145
rect 48995 -111 49029 -95
rect 48995 -161 49029 -145
rect 49199 -111 49233 -95
rect 49199 -161 49233 -145
rect 49403 -111 49437 -95
rect 49403 -161 49437 -145
rect 49607 -111 49641 -95
rect 49607 -161 49641 -145
rect 49811 -111 49845 -95
rect 49811 -161 49845 -145
rect 50015 -111 50049 -95
rect 50015 -161 50049 -145
rect 50219 -111 50253 -95
rect 50219 -161 50253 -145
rect 50423 -111 50457 -95
rect 50423 -161 50457 -145
rect 50627 -111 50661 -95
rect 50627 -161 50661 -145
rect 50831 -111 50865 -95
rect 50831 -161 50865 -145
rect 51035 -111 51069 -95
rect 51035 -161 51069 -145
rect 51239 -111 51273 -95
rect 51239 -161 51273 -145
rect 51443 -111 51477 -95
rect 51443 -161 51477 -145
rect 51647 -111 51681 -95
rect 51647 -161 51681 -145
rect 51851 -111 51885 -95
rect 51851 -161 51885 -145
rect 52055 -111 52089 -95
rect 52055 -161 52089 -145
<< viali >>
rect 35 -145 69 -111
rect 239 -145 273 -111
rect 443 -145 477 -111
rect 647 -145 681 -111
rect 851 -145 885 -111
rect 1055 -145 1089 -111
rect 1259 -145 1293 -111
rect 1463 -145 1497 -111
rect 1667 -145 1701 -111
rect 1871 -145 1905 -111
rect 2075 -145 2109 -111
rect 2279 -145 2313 -111
rect 2483 -145 2517 -111
rect 2687 -145 2721 -111
rect 2891 -145 2925 -111
rect 3095 -145 3129 -111
rect 3299 -145 3333 -111
rect 3503 -145 3537 -111
rect 3707 -145 3741 -111
rect 3911 -145 3945 -111
rect 4115 -145 4149 -111
rect 4319 -145 4353 -111
rect 4523 -145 4557 -111
rect 4727 -145 4761 -111
rect 4931 -145 4965 -111
rect 5135 -145 5169 -111
rect 5339 -145 5373 -111
rect 5543 -145 5577 -111
rect 5747 -145 5781 -111
rect 5951 -145 5985 -111
rect 6155 -145 6189 -111
rect 6359 -145 6393 -111
rect 6563 -145 6597 -111
rect 6767 -145 6801 -111
rect 6971 -145 7005 -111
rect 7175 -145 7209 -111
rect 7379 -145 7413 -111
rect 7583 -145 7617 -111
rect 7787 -145 7821 -111
rect 7991 -145 8025 -111
rect 8195 -145 8229 -111
rect 8399 -145 8433 -111
rect 8603 -145 8637 -111
rect 8807 -145 8841 -111
rect 9011 -145 9045 -111
rect 9215 -145 9249 -111
rect 9419 -145 9453 -111
rect 9623 -145 9657 -111
rect 9827 -145 9861 -111
rect 10031 -145 10065 -111
rect 10235 -145 10269 -111
rect 10439 -145 10473 -111
rect 10643 -145 10677 -111
rect 10847 -145 10881 -111
rect 11051 -145 11085 -111
rect 11255 -145 11289 -111
rect 11459 -145 11493 -111
rect 11663 -145 11697 -111
rect 11867 -145 11901 -111
rect 12071 -145 12105 -111
rect 12275 -145 12309 -111
rect 12479 -145 12513 -111
rect 12683 -145 12717 -111
rect 12887 -145 12921 -111
rect 13091 -145 13125 -111
rect 13295 -145 13329 -111
rect 13499 -145 13533 -111
rect 13703 -145 13737 -111
rect 13907 -145 13941 -111
rect 14111 -145 14145 -111
rect 14315 -145 14349 -111
rect 14519 -145 14553 -111
rect 14723 -145 14757 -111
rect 14927 -145 14961 -111
rect 15131 -145 15165 -111
rect 15335 -145 15369 -111
rect 15539 -145 15573 -111
rect 15743 -145 15777 -111
rect 15947 -145 15981 -111
rect 16151 -145 16185 -111
rect 16355 -145 16389 -111
rect 16559 -145 16593 -111
rect 16763 -145 16797 -111
rect 16967 -145 17001 -111
rect 17171 -145 17205 -111
rect 17375 -145 17409 -111
rect 17579 -145 17613 -111
rect 17783 -145 17817 -111
rect 17987 -145 18021 -111
rect 18191 -145 18225 -111
rect 18395 -145 18429 -111
rect 18599 -145 18633 -111
rect 18803 -145 18837 -111
rect 19007 -145 19041 -111
rect 19211 -145 19245 -111
rect 19415 -145 19449 -111
rect 19619 -145 19653 -111
rect 19823 -145 19857 -111
rect 20027 -145 20061 -111
rect 20231 -145 20265 -111
rect 20435 -145 20469 -111
rect 20639 -145 20673 -111
rect 20843 -145 20877 -111
rect 21047 -145 21081 -111
rect 21251 -145 21285 -111
rect 21455 -145 21489 -111
rect 21659 -145 21693 -111
rect 21863 -145 21897 -111
rect 22067 -145 22101 -111
rect 22271 -145 22305 -111
rect 22475 -145 22509 -111
rect 22679 -145 22713 -111
rect 22883 -145 22917 -111
rect 23087 -145 23121 -111
rect 23291 -145 23325 -111
rect 23495 -145 23529 -111
rect 23699 -145 23733 -111
rect 23903 -145 23937 -111
rect 24107 -145 24141 -111
rect 24311 -145 24345 -111
rect 24515 -145 24549 -111
rect 24719 -145 24753 -111
rect 24923 -145 24957 -111
rect 25127 -145 25161 -111
rect 25331 -145 25365 -111
rect 25535 -145 25569 -111
rect 25739 -145 25773 -111
rect 25943 -145 25977 -111
rect 26147 -145 26181 -111
rect 26351 -145 26385 -111
rect 26555 -145 26589 -111
rect 26759 -145 26793 -111
rect 26963 -145 26997 -111
rect 27167 -145 27201 -111
rect 27371 -145 27405 -111
rect 27575 -145 27609 -111
rect 27779 -145 27813 -111
rect 27983 -145 28017 -111
rect 28187 -145 28221 -111
rect 28391 -145 28425 -111
rect 28595 -145 28629 -111
rect 28799 -145 28833 -111
rect 29003 -145 29037 -111
rect 29207 -145 29241 -111
rect 29411 -145 29445 -111
rect 29615 -145 29649 -111
rect 29819 -145 29853 -111
rect 30023 -145 30057 -111
rect 30227 -145 30261 -111
rect 30431 -145 30465 -111
rect 30635 -145 30669 -111
rect 30839 -145 30873 -111
rect 31043 -145 31077 -111
rect 31247 -145 31281 -111
rect 31451 -145 31485 -111
rect 31655 -145 31689 -111
rect 31859 -145 31893 -111
rect 32063 -145 32097 -111
rect 32267 -145 32301 -111
rect 32471 -145 32505 -111
rect 32675 -145 32709 -111
rect 32879 -145 32913 -111
rect 33083 -145 33117 -111
rect 33287 -145 33321 -111
rect 33491 -145 33525 -111
rect 33695 -145 33729 -111
rect 33899 -145 33933 -111
rect 34103 -145 34137 -111
rect 34307 -145 34341 -111
rect 34511 -145 34545 -111
rect 34715 -145 34749 -111
rect 34919 -145 34953 -111
rect 35123 -145 35157 -111
rect 35327 -145 35361 -111
rect 35531 -145 35565 -111
rect 35735 -145 35769 -111
rect 35939 -145 35973 -111
rect 36143 -145 36177 -111
rect 36347 -145 36381 -111
rect 36551 -145 36585 -111
rect 36755 -145 36789 -111
rect 36959 -145 36993 -111
rect 37163 -145 37197 -111
rect 37367 -145 37401 -111
rect 37571 -145 37605 -111
rect 37775 -145 37809 -111
rect 37979 -145 38013 -111
rect 38183 -145 38217 -111
rect 38387 -145 38421 -111
rect 38591 -145 38625 -111
rect 38795 -145 38829 -111
rect 38999 -145 39033 -111
rect 39203 -145 39237 -111
rect 39407 -145 39441 -111
rect 39611 -145 39645 -111
rect 39815 -145 39849 -111
rect 40019 -145 40053 -111
rect 40223 -145 40257 -111
rect 40427 -145 40461 -111
rect 40631 -145 40665 -111
rect 40835 -145 40869 -111
rect 41039 -145 41073 -111
rect 41243 -145 41277 -111
rect 41447 -145 41481 -111
rect 41651 -145 41685 -111
rect 41855 -145 41889 -111
rect 42059 -145 42093 -111
rect 42263 -145 42297 -111
rect 42467 -145 42501 -111
rect 42671 -145 42705 -111
rect 42875 -145 42909 -111
rect 43079 -145 43113 -111
rect 43283 -145 43317 -111
rect 43487 -145 43521 -111
rect 43691 -145 43725 -111
rect 43895 -145 43929 -111
rect 44099 -145 44133 -111
rect 44303 -145 44337 -111
rect 44507 -145 44541 -111
rect 44711 -145 44745 -111
rect 44915 -145 44949 -111
rect 45119 -145 45153 -111
rect 45323 -145 45357 -111
rect 45527 -145 45561 -111
rect 45731 -145 45765 -111
rect 45935 -145 45969 -111
rect 46139 -145 46173 -111
rect 46343 -145 46377 -111
rect 46547 -145 46581 -111
rect 46751 -145 46785 -111
rect 46955 -145 46989 -111
rect 47159 -145 47193 -111
rect 47363 -145 47397 -111
rect 47567 -145 47601 -111
rect 47771 -145 47805 -111
rect 47975 -145 48009 -111
rect 48179 -145 48213 -111
rect 48383 -145 48417 -111
rect 48587 -145 48621 -111
rect 48791 -145 48825 -111
rect 48995 -145 49029 -111
rect 49199 -145 49233 -111
rect 49403 -145 49437 -111
rect 49607 -145 49641 -111
rect 49811 -145 49845 -111
rect 50015 -145 50049 -111
rect 50219 -145 50253 -111
rect 50423 -145 50457 -111
rect 50627 -145 50661 -111
rect 50831 -145 50865 -111
rect 51035 -145 51069 -111
rect 51239 -145 51273 -111
rect 51443 -145 51477 -111
rect 51647 -145 51681 -111
rect 51851 -145 51885 -111
rect 52055 -145 52089 -111
<< metal1 >>
rect 122 86 150 114
rect 326 86 354 114
rect 530 86 558 114
rect 734 86 762 114
rect 938 86 966 114
rect 1142 86 1170 114
rect 1346 86 1374 114
rect 1550 86 1578 114
rect 1754 86 1782 114
rect 1958 86 1986 114
rect 2162 86 2190 114
rect 2366 86 2394 114
rect 2570 86 2598 114
rect 2774 86 2802 114
rect 2978 86 3006 114
rect 3182 86 3210 114
rect 3386 86 3414 114
rect 3590 86 3618 114
rect 3794 86 3822 114
rect 3998 86 4026 114
rect 4202 86 4230 114
rect 4406 86 4434 114
rect 4610 86 4638 114
rect 4814 86 4842 114
rect 5018 86 5046 114
rect 5222 86 5250 114
rect 5426 86 5454 114
rect 5630 86 5658 114
rect 5834 86 5862 114
rect 6038 86 6066 114
rect 6242 86 6270 114
rect 6446 86 6474 114
rect 6650 86 6678 114
rect 6854 86 6882 114
rect 7058 86 7086 114
rect 7262 86 7290 114
rect 7466 86 7494 114
rect 7670 86 7698 114
rect 7874 86 7902 114
rect 8078 86 8106 114
rect 8282 86 8310 114
rect 8486 86 8514 114
rect 8690 86 8718 114
rect 8894 86 8922 114
rect 9098 86 9126 114
rect 9302 86 9330 114
rect 9506 86 9534 114
rect 9710 86 9738 114
rect 9914 86 9942 114
rect 10118 86 10146 114
rect 10322 86 10350 114
rect 10526 86 10554 114
rect 10730 86 10758 114
rect 10934 86 10962 114
rect 11138 86 11166 114
rect 11342 86 11370 114
rect 11546 86 11574 114
rect 11750 86 11778 114
rect 11954 86 11982 114
rect 12158 86 12186 114
rect 12362 86 12390 114
rect 12566 86 12594 114
rect 12770 86 12798 114
rect 12974 86 13002 114
rect 13178 86 13206 114
rect 13382 86 13410 114
rect 13586 86 13614 114
rect 13790 86 13818 114
rect 13994 86 14022 114
rect 14198 86 14226 114
rect 14402 86 14430 114
rect 14606 86 14634 114
rect 14810 86 14838 114
rect 15014 86 15042 114
rect 15218 86 15246 114
rect 15422 86 15450 114
rect 15626 86 15654 114
rect 15830 86 15858 114
rect 16034 86 16062 114
rect 16238 86 16266 114
rect 16442 86 16470 114
rect 16646 86 16674 114
rect 16850 86 16878 114
rect 17054 86 17082 114
rect 17258 86 17286 114
rect 17462 86 17490 114
rect 17666 86 17694 114
rect 17870 86 17898 114
rect 18074 86 18102 114
rect 18278 86 18306 114
rect 18482 86 18510 114
rect 18686 86 18714 114
rect 18890 86 18918 114
rect 19094 86 19122 114
rect 19298 86 19326 114
rect 19502 86 19530 114
rect 19706 86 19734 114
rect 19910 86 19938 114
rect 20114 86 20142 114
rect 20318 86 20346 114
rect 20522 86 20550 114
rect 20726 86 20754 114
rect 20930 86 20958 114
rect 21134 86 21162 114
rect 21338 86 21366 114
rect 21542 86 21570 114
rect 21746 86 21774 114
rect 21950 86 21978 114
rect 22154 86 22182 114
rect 22358 86 22386 114
rect 22562 86 22590 114
rect 22766 86 22794 114
rect 22970 86 22998 114
rect 23174 86 23202 114
rect 23378 86 23406 114
rect 23582 86 23610 114
rect 23786 86 23814 114
rect 23990 86 24018 114
rect 24194 86 24222 114
rect 24398 86 24426 114
rect 24602 86 24630 114
rect 24806 86 24834 114
rect 25010 86 25038 114
rect 25214 86 25242 114
rect 25418 86 25446 114
rect 25622 86 25650 114
rect 25826 86 25854 114
rect 26030 86 26058 114
rect 26234 86 26262 114
rect 26438 86 26466 114
rect 26642 86 26670 114
rect 26846 86 26874 114
rect 27050 86 27078 114
rect 27254 86 27282 114
rect 27458 86 27486 114
rect 27662 86 27690 114
rect 27866 86 27894 114
rect 28070 86 28098 114
rect 28274 86 28302 114
rect 28478 86 28506 114
rect 28682 86 28710 114
rect 28886 86 28914 114
rect 29090 86 29118 114
rect 29294 86 29322 114
rect 29498 86 29526 114
rect 29702 86 29730 114
rect 29906 86 29934 114
rect 30110 86 30138 114
rect 30314 86 30342 114
rect 30518 86 30546 114
rect 30722 86 30750 114
rect 30926 86 30954 114
rect 31130 86 31158 114
rect 31334 86 31362 114
rect 31538 86 31566 114
rect 31742 86 31770 114
rect 31946 86 31974 114
rect 32150 86 32178 114
rect 32354 86 32382 114
rect 32558 86 32586 114
rect 32762 86 32790 114
rect 32966 86 32994 114
rect 33170 86 33198 114
rect 33374 86 33402 114
rect 33578 86 33606 114
rect 33782 86 33810 114
rect 33986 86 34014 114
rect 34190 86 34218 114
rect 34394 86 34422 114
rect 34598 86 34626 114
rect 34802 86 34830 114
rect 35006 86 35034 114
rect 35210 86 35238 114
rect 35414 86 35442 114
rect 35618 86 35646 114
rect 35822 86 35850 114
rect 36026 86 36054 114
rect 36230 86 36258 114
rect 36434 86 36462 114
rect 36638 86 36666 114
rect 36842 86 36870 114
rect 37046 86 37074 114
rect 37250 86 37278 114
rect 37454 86 37482 114
rect 37658 86 37686 114
rect 37862 86 37890 114
rect 38066 86 38094 114
rect 38270 86 38298 114
rect 38474 86 38502 114
rect 38678 86 38706 114
rect 38882 86 38910 114
rect 39086 86 39114 114
rect 39290 86 39318 114
rect 39494 86 39522 114
rect 39698 86 39726 114
rect 39902 86 39930 114
rect 40106 86 40134 114
rect 40310 86 40338 114
rect 40514 86 40542 114
rect 40718 86 40746 114
rect 40922 86 40950 114
rect 41126 86 41154 114
rect 41330 86 41358 114
rect 41534 86 41562 114
rect 41738 86 41766 114
rect 41942 86 41970 114
rect 42146 86 42174 114
rect 42350 86 42378 114
rect 42554 86 42582 114
rect 42758 86 42786 114
rect 42962 86 42990 114
rect 43166 86 43194 114
rect 43370 86 43398 114
rect 43574 86 43602 114
rect 43778 86 43806 114
rect 43982 86 44010 114
rect 44186 86 44214 114
rect 44390 86 44418 114
rect 44594 86 44622 114
rect 44798 86 44826 114
rect 45002 86 45030 114
rect 45206 86 45234 114
rect 45410 86 45438 114
rect 45614 86 45642 114
rect 45818 86 45846 114
rect 46022 86 46050 114
rect 46226 86 46254 114
rect 46430 86 46458 114
rect 46634 86 46662 114
rect 46838 86 46866 114
rect 47042 86 47070 114
rect 47246 86 47274 114
rect 47450 86 47478 114
rect 47654 86 47682 114
rect 47858 86 47886 114
rect 48062 86 48090 114
rect 48266 86 48294 114
rect 48470 86 48498 114
rect 48674 86 48702 114
rect 48878 86 48906 114
rect 49082 86 49110 114
rect 49286 86 49314 114
rect 49490 86 49518 114
rect 49694 86 49722 114
rect 49898 86 49926 114
rect 50102 86 50130 114
rect 50306 86 50334 114
rect 50510 86 50538 114
rect 50714 86 50742 114
rect 50918 86 50946 114
rect 51122 86 51150 114
rect 51326 86 51354 114
rect 51530 86 51558 114
rect 51734 86 51762 114
rect 51938 86 51966 114
rect 52142 86 52170 114
rect 20 -154 26 -102
rect 78 -154 84 -102
rect 224 -154 230 -102
rect 282 -154 288 -102
rect 428 -154 434 -102
rect 486 -154 492 -102
rect 632 -154 638 -102
rect 690 -154 696 -102
rect 836 -154 842 -102
rect 894 -154 900 -102
rect 1040 -154 1046 -102
rect 1098 -154 1104 -102
rect 1244 -154 1250 -102
rect 1302 -154 1308 -102
rect 1448 -154 1454 -102
rect 1506 -154 1512 -102
rect 1652 -154 1658 -102
rect 1710 -154 1716 -102
rect 1856 -154 1862 -102
rect 1914 -154 1920 -102
rect 2060 -154 2066 -102
rect 2118 -154 2124 -102
rect 2264 -154 2270 -102
rect 2322 -154 2328 -102
rect 2468 -154 2474 -102
rect 2526 -154 2532 -102
rect 2672 -154 2678 -102
rect 2730 -154 2736 -102
rect 2876 -154 2882 -102
rect 2934 -154 2940 -102
rect 3080 -154 3086 -102
rect 3138 -154 3144 -102
rect 3284 -154 3290 -102
rect 3342 -154 3348 -102
rect 3488 -154 3494 -102
rect 3546 -154 3552 -102
rect 3692 -154 3698 -102
rect 3750 -154 3756 -102
rect 3896 -154 3902 -102
rect 3954 -154 3960 -102
rect 4100 -154 4106 -102
rect 4158 -154 4164 -102
rect 4304 -154 4310 -102
rect 4362 -154 4368 -102
rect 4508 -154 4514 -102
rect 4566 -154 4572 -102
rect 4712 -154 4718 -102
rect 4770 -154 4776 -102
rect 4916 -154 4922 -102
rect 4974 -154 4980 -102
rect 5120 -154 5126 -102
rect 5178 -154 5184 -102
rect 5324 -154 5330 -102
rect 5382 -154 5388 -102
rect 5528 -154 5534 -102
rect 5586 -154 5592 -102
rect 5732 -154 5738 -102
rect 5790 -154 5796 -102
rect 5936 -154 5942 -102
rect 5994 -154 6000 -102
rect 6140 -154 6146 -102
rect 6198 -154 6204 -102
rect 6344 -154 6350 -102
rect 6402 -154 6408 -102
rect 6548 -154 6554 -102
rect 6606 -154 6612 -102
rect 6752 -154 6758 -102
rect 6810 -154 6816 -102
rect 6956 -154 6962 -102
rect 7014 -154 7020 -102
rect 7160 -154 7166 -102
rect 7218 -154 7224 -102
rect 7364 -154 7370 -102
rect 7422 -154 7428 -102
rect 7568 -154 7574 -102
rect 7626 -154 7632 -102
rect 7772 -154 7778 -102
rect 7830 -154 7836 -102
rect 7976 -154 7982 -102
rect 8034 -154 8040 -102
rect 8180 -154 8186 -102
rect 8238 -154 8244 -102
rect 8384 -154 8390 -102
rect 8442 -154 8448 -102
rect 8588 -154 8594 -102
rect 8646 -154 8652 -102
rect 8792 -154 8798 -102
rect 8850 -154 8856 -102
rect 8996 -154 9002 -102
rect 9054 -154 9060 -102
rect 9200 -154 9206 -102
rect 9258 -154 9264 -102
rect 9404 -154 9410 -102
rect 9462 -154 9468 -102
rect 9608 -154 9614 -102
rect 9666 -154 9672 -102
rect 9812 -154 9818 -102
rect 9870 -154 9876 -102
rect 10016 -154 10022 -102
rect 10074 -154 10080 -102
rect 10220 -154 10226 -102
rect 10278 -154 10284 -102
rect 10424 -154 10430 -102
rect 10482 -154 10488 -102
rect 10628 -154 10634 -102
rect 10686 -154 10692 -102
rect 10832 -154 10838 -102
rect 10890 -154 10896 -102
rect 11036 -154 11042 -102
rect 11094 -154 11100 -102
rect 11240 -154 11246 -102
rect 11298 -154 11304 -102
rect 11444 -154 11450 -102
rect 11502 -154 11508 -102
rect 11648 -154 11654 -102
rect 11706 -154 11712 -102
rect 11852 -154 11858 -102
rect 11910 -154 11916 -102
rect 12056 -154 12062 -102
rect 12114 -154 12120 -102
rect 12260 -154 12266 -102
rect 12318 -154 12324 -102
rect 12464 -154 12470 -102
rect 12522 -154 12528 -102
rect 12668 -154 12674 -102
rect 12726 -154 12732 -102
rect 12872 -154 12878 -102
rect 12930 -154 12936 -102
rect 13076 -154 13082 -102
rect 13134 -154 13140 -102
rect 13280 -154 13286 -102
rect 13338 -154 13344 -102
rect 13484 -154 13490 -102
rect 13542 -154 13548 -102
rect 13688 -154 13694 -102
rect 13746 -154 13752 -102
rect 13892 -154 13898 -102
rect 13950 -154 13956 -102
rect 14096 -154 14102 -102
rect 14154 -154 14160 -102
rect 14300 -154 14306 -102
rect 14358 -154 14364 -102
rect 14504 -154 14510 -102
rect 14562 -154 14568 -102
rect 14708 -154 14714 -102
rect 14766 -154 14772 -102
rect 14912 -154 14918 -102
rect 14970 -154 14976 -102
rect 15116 -154 15122 -102
rect 15174 -154 15180 -102
rect 15320 -154 15326 -102
rect 15378 -154 15384 -102
rect 15524 -154 15530 -102
rect 15582 -154 15588 -102
rect 15728 -154 15734 -102
rect 15786 -154 15792 -102
rect 15932 -154 15938 -102
rect 15990 -154 15996 -102
rect 16136 -154 16142 -102
rect 16194 -154 16200 -102
rect 16340 -154 16346 -102
rect 16398 -154 16404 -102
rect 16544 -154 16550 -102
rect 16602 -154 16608 -102
rect 16748 -154 16754 -102
rect 16806 -154 16812 -102
rect 16952 -154 16958 -102
rect 17010 -154 17016 -102
rect 17156 -154 17162 -102
rect 17214 -154 17220 -102
rect 17360 -154 17366 -102
rect 17418 -154 17424 -102
rect 17564 -154 17570 -102
rect 17622 -154 17628 -102
rect 17768 -154 17774 -102
rect 17826 -154 17832 -102
rect 17972 -154 17978 -102
rect 18030 -154 18036 -102
rect 18176 -154 18182 -102
rect 18234 -154 18240 -102
rect 18380 -154 18386 -102
rect 18438 -154 18444 -102
rect 18584 -154 18590 -102
rect 18642 -154 18648 -102
rect 18788 -154 18794 -102
rect 18846 -154 18852 -102
rect 18992 -154 18998 -102
rect 19050 -154 19056 -102
rect 19196 -154 19202 -102
rect 19254 -154 19260 -102
rect 19400 -154 19406 -102
rect 19458 -154 19464 -102
rect 19604 -154 19610 -102
rect 19662 -154 19668 -102
rect 19808 -154 19814 -102
rect 19866 -154 19872 -102
rect 20012 -154 20018 -102
rect 20070 -154 20076 -102
rect 20216 -154 20222 -102
rect 20274 -154 20280 -102
rect 20420 -154 20426 -102
rect 20478 -154 20484 -102
rect 20624 -154 20630 -102
rect 20682 -154 20688 -102
rect 20828 -154 20834 -102
rect 20886 -154 20892 -102
rect 21032 -154 21038 -102
rect 21090 -154 21096 -102
rect 21236 -154 21242 -102
rect 21294 -154 21300 -102
rect 21440 -154 21446 -102
rect 21498 -154 21504 -102
rect 21644 -154 21650 -102
rect 21702 -154 21708 -102
rect 21848 -154 21854 -102
rect 21906 -154 21912 -102
rect 22052 -154 22058 -102
rect 22110 -154 22116 -102
rect 22256 -154 22262 -102
rect 22314 -154 22320 -102
rect 22460 -154 22466 -102
rect 22518 -154 22524 -102
rect 22664 -154 22670 -102
rect 22722 -154 22728 -102
rect 22868 -154 22874 -102
rect 22926 -154 22932 -102
rect 23072 -154 23078 -102
rect 23130 -154 23136 -102
rect 23276 -154 23282 -102
rect 23334 -154 23340 -102
rect 23480 -154 23486 -102
rect 23538 -154 23544 -102
rect 23684 -154 23690 -102
rect 23742 -154 23748 -102
rect 23888 -154 23894 -102
rect 23946 -154 23952 -102
rect 24092 -154 24098 -102
rect 24150 -154 24156 -102
rect 24296 -154 24302 -102
rect 24354 -154 24360 -102
rect 24500 -154 24506 -102
rect 24558 -154 24564 -102
rect 24704 -154 24710 -102
rect 24762 -154 24768 -102
rect 24908 -154 24914 -102
rect 24966 -154 24972 -102
rect 25112 -154 25118 -102
rect 25170 -154 25176 -102
rect 25316 -154 25322 -102
rect 25374 -154 25380 -102
rect 25520 -154 25526 -102
rect 25578 -154 25584 -102
rect 25724 -154 25730 -102
rect 25782 -154 25788 -102
rect 25928 -154 25934 -102
rect 25986 -154 25992 -102
rect 26132 -154 26138 -102
rect 26190 -154 26196 -102
rect 26336 -154 26342 -102
rect 26394 -154 26400 -102
rect 26540 -154 26546 -102
rect 26598 -154 26604 -102
rect 26744 -154 26750 -102
rect 26802 -154 26808 -102
rect 26948 -154 26954 -102
rect 27006 -154 27012 -102
rect 27152 -154 27158 -102
rect 27210 -154 27216 -102
rect 27356 -154 27362 -102
rect 27414 -154 27420 -102
rect 27560 -154 27566 -102
rect 27618 -154 27624 -102
rect 27764 -154 27770 -102
rect 27822 -154 27828 -102
rect 27968 -154 27974 -102
rect 28026 -154 28032 -102
rect 28172 -154 28178 -102
rect 28230 -154 28236 -102
rect 28376 -154 28382 -102
rect 28434 -154 28440 -102
rect 28580 -154 28586 -102
rect 28638 -154 28644 -102
rect 28784 -154 28790 -102
rect 28842 -154 28848 -102
rect 28988 -154 28994 -102
rect 29046 -154 29052 -102
rect 29192 -154 29198 -102
rect 29250 -154 29256 -102
rect 29396 -154 29402 -102
rect 29454 -154 29460 -102
rect 29600 -154 29606 -102
rect 29658 -154 29664 -102
rect 29804 -154 29810 -102
rect 29862 -154 29868 -102
rect 30008 -154 30014 -102
rect 30066 -154 30072 -102
rect 30212 -154 30218 -102
rect 30270 -154 30276 -102
rect 30416 -154 30422 -102
rect 30474 -154 30480 -102
rect 30620 -154 30626 -102
rect 30678 -154 30684 -102
rect 30824 -154 30830 -102
rect 30882 -154 30888 -102
rect 31028 -154 31034 -102
rect 31086 -154 31092 -102
rect 31232 -154 31238 -102
rect 31290 -154 31296 -102
rect 31436 -154 31442 -102
rect 31494 -154 31500 -102
rect 31640 -154 31646 -102
rect 31698 -154 31704 -102
rect 31844 -154 31850 -102
rect 31902 -154 31908 -102
rect 32048 -154 32054 -102
rect 32106 -154 32112 -102
rect 32252 -154 32258 -102
rect 32310 -154 32316 -102
rect 32456 -154 32462 -102
rect 32514 -154 32520 -102
rect 32660 -154 32666 -102
rect 32718 -154 32724 -102
rect 32864 -154 32870 -102
rect 32922 -154 32928 -102
rect 33068 -154 33074 -102
rect 33126 -154 33132 -102
rect 33272 -154 33278 -102
rect 33330 -154 33336 -102
rect 33476 -154 33482 -102
rect 33534 -154 33540 -102
rect 33680 -154 33686 -102
rect 33738 -154 33744 -102
rect 33884 -154 33890 -102
rect 33942 -154 33948 -102
rect 34088 -154 34094 -102
rect 34146 -154 34152 -102
rect 34292 -154 34298 -102
rect 34350 -154 34356 -102
rect 34496 -154 34502 -102
rect 34554 -154 34560 -102
rect 34700 -154 34706 -102
rect 34758 -154 34764 -102
rect 34904 -154 34910 -102
rect 34962 -154 34968 -102
rect 35108 -154 35114 -102
rect 35166 -154 35172 -102
rect 35312 -154 35318 -102
rect 35370 -154 35376 -102
rect 35516 -154 35522 -102
rect 35574 -154 35580 -102
rect 35720 -154 35726 -102
rect 35778 -154 35784 -102
rect 35924 -154 35930 -102
rect 35982 -154 35988 -102
rect 36128 -154 36134 -102
rect 36186 -154 36192 -102
rect 36332 -154 36338 -102
rect 36390 -154 36396 -102
rect 36536 -154 36542 -102
rect 36594 -154 36600 -102
rect 36740 -154 36746 -102
rect 36798 -154 36804 -102
rect 36944 -154 36950 -102
rect 37002 -154 37008 -102
rect 37148 -154 37154 -102
rect 37206 -154 37212 -102
rect 37352 -154 37358 -102
rect 37410 -154 37416 -102
rect 37556 -154 37562 -102
rect 37614 -154 37620 -102
rect 37760 -154 37766 -102
rect 37818 -154 37824 -102
rect 37964 -154 37970 -102
rect 38022 -154 38028 -102
rect 38168 -154 38174 -102
rect 38226 -154 38232 -102
rect 38372 -154 38378 -102
rect 38430 -154 38436 -102
rect 38576 -154 38582 -102
rect 38634 -154 38640 -102
rect 38780 -154 38786 -102
rect 38838 -154 38844 -102
rect 38984 -154 38990 -102
rect 39042 -154 39048 -102
rect 39188 -154 39194 -102
rect 39246 -154 39252 -102
rect 39392 -154 39398 -102
rect 39450 -154 39456 -102
rect 39596 -154 39602 -102
rect 39654 -154 39660 -102
rect 39800 -154 39806 -102
rect 39858 -154 39864 -102
rect 40004 -154 40010 -102
rect 40062 -154 40068 -102
rect 40208 -154 40214 -102
rect 40266 -154 40272 -102
rect 40412 -154 40418 -102
rect 40470 -154 40476 -102
rect 40616 -154 40622 -102
rect 40674 -154 40680 -102
rect 40820 -154 40826 -102
rect 40878 -154 40884 -102
rect 41024 -154 41030 -102
rect 41082 -154 41088 -102
rect 41228 -154 41234 -102
rect 41286 -154 41292 -102
rect 41432 -154 41438 -102
rect 41490 -154 41496 -102
rect 41636 -154 41642 -102
rect 41694 -154 41700 -102
rect 41840 -154 41846 -102
rect 41898 -154 41904 -102
rect 42044 -154 42050 -102
rect 42102 -154 42108 -102
rect 42248 -154 42254 -102
rect 42306 -154 42312 -102
rect 42452 -154 42458 -102
rect 42510 -154 42516 -102
rect 42656 -154 42662 -102
rect 42714 -154 42720 -102
rect 42860 -154 42866 -102
rect 42918 -154 42924 -102
rect 43064 -154 43070 -102
rect 43122 -154 43128 -102
rect 43268 -154 43274 -102
rect 43326 -154 43332 -102
rect 43472 -154 43478 -102
rect 43530 -154 43536 -102
rect 43676 -154 43682 -102
rect 43734 -154 43740 -102
rect 43880 -154 43886 -102
rect 43938 -154 43944 -102
rect 44084 -154 44090 -102
rect 44142 -154 44148 -102
rect 44288 -154 44294 -102
rect 44346 -154 44352 -102
rect 44492 -154 44498 -102
rect 44550 -154 44556 -102
rect 44696 -154 44702 -102
rect 44754 -154 44760 -102
rect 44900 -154 44906 -102
rect 44958 -154 44964 -102
rect 45104 -154 45110 -102
rect 45162 -154 45168 -102
rect 45308 -154 45314 -102
rect 45366 -154 45372 -102
rect 45512 -154 45518 -102
rect 45570 -154 45576 -102
rect 45716 -154 45722 -102
rect 45774 -154 45780 -102
rect 45920 -154 45926 -102
rect 45978 -154 45984 -102
rect 46124 -154 46130 -102
rect 46182 -154 46188 -102
rect 46328 -154 46334 -102
rect 46386 -154 46392 -102
rect 46532 -154 46538 -102
rect 46590 -154 46596 -102
rect 46736 -154 46742 -102
rect 46794 -154 46800 -102
rect 46940 -154 46946 -102
rect 46998 -154 47004 -102
rect 47144 -154 47150 -102
rect 47202 -154 47208 -102
rect 47348 -154 47354 -102
rect 47406 -154 47412 -102
rect 47552 -154 47558 -102
rect 47610 -154 47616 -102
rect 47756 -154 47762 -102
rect 47814 -154 47820 -102
rect 47960 -154 47966 -102
rect 48018 -154 48024 -102
rect 48164 -154 48170 -102
rect 48222 -154 48228 -102
rect 48368 -154 48374 -102
rect 48426 -154 48432 -102
rect 48572 -154 48578 -102
rect 48630 -154 48636 -102
rect 48776 -154 48782 -102
rect 48834 -154 48840 -102
rect 48980 -154 48986 -102
rect 49038 -154 49044 -102
rect 49184 -154 49190 -102
rect 49242 -154 49248 -102
rect 49388 -154 49394 -102
rect 49446 -154 49452 -102
rect 49592 -154 49598 -102
rect 49650 -154 49656 -102
rect 49796 -154 49802 -102
rect 49854 -154 49860 -102
rect 50000 -154 50006 -102
rect 50058 -154 50064 -102
rect 50204 -154 50210 -102
rect 50262 -154 50268 -102
rect 50408 -154 50414 -102
rect 50466 -154 50472 -102
rect 50612 -154 50618 -102
rect 50670 -154 50676 -102
rect 50816 -154 50822 -102
rect 50874 -154 50880 -102
rect 51020 -154 51026 -102
rect 51078 -154 51084 -102
rect 51224 -154 51230 -102
rect 51282 -154 51288 -102
rect 51428 -154 51434 -102
rect 51486 -154 51492 -102
rect 51632 -154 51638 -102
rect 51690 -154 51696 -102
rect 51836 -154 51842 -102
rect 51894 -154 51900 -102
rect 52040 -154 52046 -102
rect 52098 -154 52104 -102
<< via1 >>
rect 26 -111 78 -102
rect 26 -145 35 -111
rect 35 -145 69 -111
rect 69 -145 78 -111
rect 26 -154 78 -145
rect 230 -111 282 -102
rect 230 -145 239 -111
rect 239 -145 273 -111
rect 273 -145 282 -111
rect 230 -154 282 -145
rect 434 -111 486 -102
rect 434 -145 443 -111
rect 443 -145 477 -111
rect 477 -145 486 -111
rect 434 -154 486 -145
rect 638 -111 690 -102
rect 638 -145 647 -111
rect 647 -145 681 -111
rect 681 -145 690 -111
rect 638 -154 690 -145
rect 842 -111 894 -102
rect 842 -145 851 -111
rect 851 -145 885 -111
rect 885 -145 894 -111
rect 842 -154 894 -145
rect 1046 -111 1098 -102
rect 1046 -145 1055 -111
rect 1055 -145 1089 -111
rect 1089 -145 1098 -111
rect 1046 -154 1098 -145
rect 1250 -111 1302 -102
rect 1250 -145 1259 -111
rect 1259 -145 1293 -111
rect 1293 -145 1302 -111
rect 1250 -154 1302 -145
rect 1454 -111 1506 -102
rect 1454 -145 1463 -111
rect 1463 -145 1497 -111
rect 1497 -145 1506 -111
rect 1454 -154 1506 -145
rect 1658 -111 1710 -102
rect 1658 -145 1667 -111
rect 1667 -145 1701 -111
rect 1701 -145 1710 -111
rect 1658 -154 1710 -145
rect 1862 -111 1914 -102
rect 1862 -145 1871 -111
rect 1871 -145 1905 -111
rect 1905 -145 1914 -111
rect 1862 -154 1914 -145
rect 2066 -111 2118 -102
rect 2066 -145 2075 -111
rect 2075 -145 2109 -111
rect 2109 -145 2118 -111
rect 2066 -154 2118 -145
rect 2270 -111 2322 -102
rect 2270 -145 2279 -111
rect 2279 -145 2313 -111
rect 2313 -145 2322 -111
rect 2270 -154 2322 -145
rect 2474 -111 2526 -102
rect 2474 -145 2483 -111
rect 2483 -145 2517 -111
rect 2517 -145 2526 -111
rect 2474 -154 2526 -145
rect 2678 -111 2730 -102
rect 2678 -145 2687 -111
rect 2687 -145 2721 -111
rect 2721 -145 2730 -111
rect 2678 -154 2730 -145
rect 2882 -111 2934 -102
rect 2882 -145 2891 -111
rect 2891 -145 2925 -111
rect 2925 -145 2934 -111
rect 2882 -154 2934 -145
rect 3086 -111 3138 -102
rect 3086 -145 3095 -111
rect 3095 -145 3129 -111
rect 3129 -145 3138 -111
rect 3086 -154 3138 -145
rect 3290 -111 3342 -102
rect 3290 -145 3299 -111
rect 3299 -145 3333 -111
rect 3333 -145 3342 -111
rect 3290 -154 3342 -145
rect 3494 -111 3546 -102
rect 3494 -145 3503 -111
rect 3503 -145 3537 -111
rect 3537 -145 3546 -111
rect 3494 -154 3546 -145
rect 3698 -111 3750 -102
rect 3698 -145 3707 -111
rect 3707 -145 3741 -111
rect 3741 -145 3750 -111
rect 3698 -154 3750 -145
rect 3902 -111 3954 -102
rect 3902 -145 3911 -111
rect 3911 -145 3945 -111
rect 3945 -145 3954 -111
rect 3902 -154 3954 -145
rect 4106 -111 4158 -102
rect 4106 -145 4115 -111
rect 4115 -145 4149 -111
rect 4149 -145 4158 -111
rect 4106 -154 4158 -145
rect 4310 -111 4362 -102
rect 4310 -145 4319 -111
rect 4319 -145 4353 -111
rect 4353 -145 4362 -111
rect 4310 -154 4362 -145
rect 4514 -111 4566 -102
rect 4514 -145 4523 -111
rect 4523 -145 4557 -111
rect 4557 -145 4566 -111
rect 4514 -154 4566 -145
rect 4718 -111 4770 -102
rect 4718 -145 4727 -111
rect 4727 -145 4761 -111
rect 4761 -145 4770 -111
rect 4718 -154 4770 -145
rect 4922 -111 4974 -102
rect 4922 -145 4931 -111
rect 4931 -145 4965 -111
rect 4965 -145 4974 -111
rect 4922 -154 4974 -145
rect 5126 -111 5178 -102
rect 5126 -145 5135 -111
rect 5135 -145 5169 -111
rect 5169 -145 5178 -111
rect 5126 -154 5178 -145
rect 5330 -111 5382 -102
rect 5330 -145 5339 -111
rect 5339 -145 5373 -111
rect 5373 -145 5382 -111
rect 5330 -154 5382 -145
rect 5534 -111 5586 -102
rect 5534 -145 5543 -111
rect 5543 -145 5577 -111
rect 5577 -145 5586 -111
rect 5534 -154 5586 -145
rect 5738 -111 5790 -102
rect 5738 -145 5747 -111
rect 5747 -145 5781 -111
rect 5781 -145 5790 -111
rect 5738 -154 5790 -145
rect 5942 -111 5994 -102
rect 5942 -145 5951 -111
rect 5951 -145 5985 -111
rect 5985 -145 5994 -111
rect 5942 -154 5994 -145
rect 6146 -111 6198 -102
rect 6146 -145 6155 -111
rect 6155 -145 6189 -111
rect 6189 -145 6198 -111
rect 6146 -154 6198 -145
rect 6350 -111 6402 -102
rect 6350 -145 6359 -111
rect 6359 -145 6393 -111
rect 6393 -145 6402 -111
rect 6350 -154 6402 -145
rect 6554 -111 6606 -102
rect 6554 -145 6563 -111
rect 6563 -145 6597 -111
rect 6597 -145 6606 -111
rect 6554 -154 6606 -145
rect 6758 -111 6810 -102
rect 6758 -145 6767 -111
rect 6767 -145 6801 -111
rect 6801 -145 6810 -111
rect 6758 -154 6810 -145
rect 6962 -111 7014 -102
rect 6962 -145 6971 -111
rect 6971 -145 7005 -111
rect 7005 -145 7014 -111
rect 6962 -154 7014 -145
rect 7166 -111 7218 -102
rect 7166 -145 7175 -111
rect 7175 -145 7209 -111
rect 7209 -145 7218 -111
rect 7166 -154 7218 -145
rect 7370 -111 7422 -102
rect 7370 -145 7379 -111
rect 7379 -145 7413 -111
rect 7413 -145 7422 -111
rect 7370 -154 7422 -145
rect 7574 -111 7626 -102
rect 7574 -145 7583 -111
rect 7583 -145 7617 -111
rect 7617 -145 7626 -111
rect 7574 -154 7626 -145
rect 7778 -111 7830 -102
rect 7778 -145 7787 -111
rect 7787 -145 7821 -111
rect 7821 -145 7830 -111
rect 7778 -154 7830 -145
rect 7982 -111 8034 -102
rect 7982 -145 7991 -111
rect 7991 -145 8025 -111
rect 8025 -145 8034 -111
rect 7982 -154 8034 -145
rect 8186 -111 8238 -102
rect 8186 -145 8195 -111
rect 8195 -145 8229 -111
rect 8229 -145 8238 -111
rect 8186 -154 8238 -145
rect 8390 -111 8442 -102
rect 8390 -145 8399 -111
rect 8399 -145 8433 -111
rect 8433 -145 8442 -111
rect 8390 -154 8442 -145
rect 8594 -111 8646 -102
rect 8594 -145 8603 -111
rect 8603 -145 8637 -111
rect 8637 -145 8646 -111
rect 8594 -154 8646 -145
rect 8798 -111 8850 -102
rect 8798 -145 8807 -111
rect 8807 -145 8841 -111
rect 8841 -145 8850 -111
rect 8798 -154 8850 -145
rect 9002 -111 9054 -102
rect 9002 -145 9011 -111
rect 9011 -145 9045 -111
rect 9045 -145 9054 -111
rect 9002 -154 9054 -145
rect 9206 -111 9258 -102
rect 9206 -145 9215 -111
rect 9215 -145 9249 -111
rect 9249 -145 9258 -111
rect 9206 -154 9258 -145
rect 9410 -111 9462 -102
rect 9410 -145 9419 -111
rect 9419 -145 9453 -111
rect 9453 -145 9462 -111
rect 9410 -154 9462 -145
rect 9614 -111 9666 -102
rect 9614 -145 9623 -111
rect 9623 -145 9657 -111
rect 9657 -145 9666 -111
rect 9614 -154 9666 -145
rect 9818 -111 9870 -102
rect 9818 -145 9827 -111
rect 9827 -145 9861 -111
rect 9861 -145 9870 -111
rect 9818 -154 9870 -145
rect 10022 -111 10074 -102
rect 10022 -145 10031 -111
rect 10031 -145 10065 -111
rect 10065 -145 10074 -111
rect 10022 -154 10074 -145
rect 10226 -111 10278 -102
rect 10226 -145 10235 -111
rect 10235 -145 10269 -111
rect 10269 -145 10278 -111
rect 10226 -154 10278 -145
rect 10430 -111 10482 -102
rect 10430 -145 10439 -111
rect 10439 -145 10473 -111
rect 10473 -145 10482 -111
rect 10430 -154 10482 -145
rect 10634 -111 10686 -102
rect 10634 -145 10643 -111
rect 10643 -145 10677 -111
rect 10677 -145 10686 -111
rect 10634 -154 10686 -145
rect 10838 -111 10890 -102
rect 10838 -145 10847 -111
rect 10847 -145 10881 -111
rect 10881 -145 10890 -111
rect 10838 -154 10890 -145
rect 11042 -111 11094 -102
rect 11042 -145 11051 -111
rect 11051 -145 11085 -111
rect 11085 -145 11094 -111
rect 11042 -154 11094 -145
rect 11246 -111 11298 -102
rect 11246 -145 11255 -111
rect 11255 -145 11289 -111
rect 11289 -145 11298 -111
rect 11246 -154 11298 -145
rect 11450 -111 11502 -102
rect 11450 -145 11459 -111
rect 11459 -145 11493 -111
rect 11493 -145 11502 -111
rect 11450 -154 11502 -145
rect 11654 -111 11706 -102
rect 11654 -145 11663 -111
rect 11663 -145 11697 -111
rect 11697 -145 11706 -111
rect 11654 -154 11706 -145
rect 11858 -111 11910 -102
rect 11858 -145 11867 -111
rect 11867 -145 11901 -111
rect 11901 -145 11910 -111
rect 11858 -154 11910 -145
rect 12062 -111 12114 -102
rect 12062 -145 12071 -111
rect 12071 -145 12105 -111
rect 12105 -145 12114 -111
rect 12062 -154 12114 -145
rect 12266 -111 12318 -102
rect 12266 -145 12275 -111
rect 12275 -145 12309 -111
rect 12309 -145 12318 -111
rect 12266 -154 12318 -145
rect 12470 -111 12522 -102
rect 12470 -145 12479 -111
rect 12479 -145 12513 -111
rect 12513 -145 12522 -111
rect 12470 -154 12522 -145
rect 12674 -111 12726 -102
rect 12674 -145 12683 -111
rect 12683 -145 12717 -111
rect 12717 -145 12726 -111
rect 12674 -154 12726 -145
rect 12878 -111 12930 -102
rect 12878 -145 12887 -111
rect 12887 -145 12921 -111
rect 12921 -145 12930 -111
rect 12878 -154 12930 -145
rect 13082 -111 13134 -102
rect 13082 -145 13091 -111
rect 13091 -145 13125 -111
rect 13125 -145 13134 -111
rect 13082 -154 13134 -145
rect 13286 -111 13338 -102
rect 13286 -145 13295 -111
rect 13295 -145 13329 -111
rect 13329 -145 13338 -111
rect 13286 -154 13338 -145
rect 13490 -111 13542 -102
rect 13490 -145 13499 -111
rect 13499 -145 13533 -111
rect 13533 -145 13542 -111
rect 13490 -154 13542 -145
rect 13694 -111 13746 -102
rect 13694 -145 13703 -111
rect 13703 -145 13737 -111
rect 13737 -145 13746 -111
rect 13694 -154 13746 -145
rect 13898 -111 13950 -102
rect 13898 -145 13907 -111
rect 13907 -145 13941 -111
rect 13941 -145 13950 -111
rect 13898 -154 13950 -145
rect 14102 -111 14154 -102
rect 14102 -145 14111 -111
rect 14111 -145 14145 -111
rect 14145 -145 14154 -111
rect 14102 -154 14154 -145
rect 14306 -111 14358 -102
rect 14306 -145 14315 -111
rect 14315 -145 14349 -111
rect 14349 -145 14358 -111
rect 14306 -154 14358 -145
rect 14510 -111 14562 -102
rect 14510 -145 14519 -111
rect 14519 -145 14553 -111
rect 14553 -145 14562 -111
rect 14510 -154 14562 -145
rect 14714 -111 14766 -102
rect 14714 -145 14723 -111
rect 14723 -145 14757 -111
rect 14757 -145 14766 -111
rect 14714 -154 14766 -145
rect 14918 -111 14970 -102
rect 14918 -145 14927 -111
rect 14927 -145 14961 -111
rect 14961 -145 14970 -111
rect 14918 -154 14970 -145
rect 15122 -111 15174 -102
rect 15122 -145 15131 -111
rect 15131 -145 15165 -111
rect 15165 -145 15174 -111
rect 15122 -154 15174 -145
rect 15326 -111 15378 -102
rect 15326 -145 15335 -111
rect 15335 -145 15369 -111
rect 15369 -145 15378 -111
rect 15326 -154 15378 -145
rect 15530 -111 15582 -102
rect 15530 -145 15539 -111
rect 15539 -145 15573 -111
rect 15573 -145 15582 -111
rect 15530 -154 15582 -145
rect 15734 -111 15786 -102
rect 15734 -145 15743 -111
rect 15743 -145 15777 -111
rect 15777 -145 15786 -111
rect 15734 -154 15786 -145
rect 15938 -111 15990 -102
rect 15938 -145 15947 -111
rect 15947 -145 15981 -111
rect 15981 -145 15990 -111
rect 15938 -154 15990 -145
rect 16142 -111 16194 -102
rect 16142 -145 16151 -111
rect 16151 -145 16185 -111
rect 16185 -145 16194 -111
rect 16142 -154 16194 -145
rect 16346 -111 16398 -102
rect 16346 -145 16355 -111
rect 16355 -145 16389 -111
rect 16389 -145 16398 -111
rect 16346 -154 16398 -145
rect 16550 -111 16602 -102
rect 16550 -145 16559 -111
rect 16559 -145 16593 -111
rect 16593 -145 16602 -111
rect 16550 -154 16602 -145
rect 16754 -111 16806 -102
rect 16754 -145 16763 -111
rect 16763 -145 16797 -111
rect 16797 -145 16806 -111
rect 16754 -154 16806 -145
rect 16958 -111 17010 -102
rect 16958 -145 16967 -111
rect 16967 -145 17001 -111
rect 17001 -145 17010 -111
rect 16958 -154 17010 -145
rect 17162 -111 17214 -102
rect 17162 -145 17171 -111
rect 17171 -145 17205 -111
rect 17205 -145 17214 -111
rect 17162 -154 17214 -145
rect 17366 -111 17418 -102
rect 17366 -145 17375 -111
rect 17375 -145 17409 -111
rect 17409 -145 17418 -111
rect 17366 -154 17418 -145
rect 17570 -111 17622 -102
rect 17570 -145 17579 -111
rect 17579 -145 17613 -111
rect 17613 -145 17622 -111
rect 17570 -154 17622 -145
rect 17774 -111 17826 -102
rect 17774 -145 17783 -111
rect 17783 -145 17817 -111
rect 17817 -145 17826 -111
rect 17774 -154 17826 -145
rect 17978 -111 18030 -102
rect 17978 -145 17987 -111
rect 17987 -145 18021 -111
rect 18021 -145 18030 -111
rect 17978 -154 18030 -145
rect 18182 -111 18234 -102
rect 18182 -145 18191 -111
rect 18191 -145 18225 -111
rect 18225 -145 18234 -111
rect 18182 -154 18234 -145
rect 18386 -111 18438 -102
rect 18386 -145 18395 -111
rect 18395 -145 18429 -111
rect 18429 -145 18438 -111
rect 18386 -154 18438 -145
rect 18590 -111 18642 -102
rect 18590 -145 18599 -111
rect 18599 -145 18633 -111
rect 18633 -145 18642 -111
rect 18590 -154 18642 -145
rect 18794 -111 18846 -102
rect 18794 -145 18803 -111
rect 18803 -145 18837 -111
rect 18837 -145 18846 -111
rect 18794 -154 18846 -145
rect 18998 -111 19050 -102
rect 18998 -145 19007 -111
rect 19007 -145 19041 -111
rect 19041 -145 19050 -111
rect 18998 -154 19050 -145
rect 19202 -111 19254 -102
rect 19202 -145 19211 -111
rect 19211 -145 19245 -111
rect 19245 -145 19254 -111
rect 19202 -154 19254 -145
rect 19406 -111 19458 -102
rect 19406 -145 19415 -111
rect 19415 -145 19449 -111
rect 19449 -145 19458 -111
rect 19406 -154 19458 -145
rect 19610 -111 19662 -102
rect 19610 -145 19619 -111
rect 19619 -145 19653 -111
rect 19653 -145 19662 -111
rect 19610 -154 19662 -145
rect 19814 -111 19866 -102
rect 19814 -145 19823 -111
rect 19823 -145 19857 -111
rect 19857 -145 19866 -111
rect 19814 -154 19866 -145
rect 20018 -111 20070 -102
rect 20018 -145 20027 -111
rect 20027 -145 20061 -111
rect 20061 -145 20070 -111
rect 20018 -154 20070 -145
rect 20222 -111 20274 -102
rect 20222 -145 20231 -111
rect 20231 -145 20265 -111
rect 20265 -145 20274 -111
rect 20222 -154 20274 -145
rect 20426 -111 20478 -102
rect 20426 -145 20435 -111
rect 20435 -145 20469 -111
rect 20469 -145 20478 -111
rect 20426 -154 20478 -145
rect 20630 -111 20682 -102
rect 20630 -145 20639 -111
rect 20639 -145 20673 -111
rect 20673 -145 20682 -111
rect 20630 -154 20682 -145
rect 20834 -111 20886 -102
rect 20834 -145 20843 -111
rect 20843 -145 20877 -111
rect 20877 -145 20886 -111
rect 20834 -154 20886 -145
rect 21038 -111 21090 -102
rect 21038 -145 21047 -111
rect 21047 -145 21081 -111
rect 21081 -145 21090 -111
rect 21038 -154 21090 -145
rect 21242 -111 21294 -102
rect 21242 -145 21251 -111
rect 21251 -145 21285 -111
rect 21285 -145 21294 -111
rect 21242 -154 21294 -145
rect 21446 -111 21498 -102
rect 21446 -145 21455 -111
rect 21455 -145 21489 -111
rect 21489 -145 21498 -111
rect 21446 -154 21498 -145
rect 21650 -111 21702 -102
rect 21650 -145 21659 -111
rect 21659 -145 21693 -111
rect 21693 -145 21702 -111
rect 21650 -154 21702 -145
rect 21854 -111 21906 -102
rect 21854 -145 21863 -111
rect 21863 -145 21897 -111
rect 21897 -145 21906 -111
rect 21854 -154 21906 -145
rect 22058 -111 22110 -102
rect 22058 -145 22067 -111
rect 22067 -145 22101 -111
rect 22101 -145 22110 -111
rect 22058 -154 22110 -145
rect 22262 -111 22314 -102
rect 22262 -145 22271 -111
rect 22271 -145 22305 -111
rect 22305 -145 22314 -111
rect 22262 -154 22314 -145
rect 22466 -111 22518 -102
rect 22466 -145 22475 -111
rect 22475 -145 22509 -111
rect 22509 -145 22518 -111
rect 22466 -154 22518 -145
rect 22670 -111 22722 -102
rect 22670 -145 22679 -111
rect 22679 -145 22713 -111
rect 22713 -145 22722 -111
rect 22670 -154 22722 -145
rect 22874 -111 22926 -102
rect 22874 -145 22883 -111
rect 22883 -145 22917 -111
rect 22917 -145 22926 -111
rect 22874 -154 22926 -145
rect 23078 -111 23130 -102
rect 23078 -145 23087 -111
rect 23087 -145 23121 -111
rect 23121 -145 23130 -111
rect 23078 -154 23130 -145
rect 23282 -111 23334 -102
rect 23282 -145 23291 -111
rect 23291 -145 23325 -111
rect 23325 -145 23334 -111
rect 23282 -154 23334 -145
rect 23486 -111 23538 -102
rect 23486 -145 23495 -111
rect 23495 -145 23529 -111
rect 23529 -145 23538 -111
rect 23486 -154 23538 -145
rect 23690 -111 23742 -102
rect 23690 -145 23699 -111
rect 23699 -145 23733 -111
rect 23733 -145 23742 -111
rect 23690 -154 23742 -145
rect 23894 -111 23946 -102
rect 23894 -145 23903 -111
rect 23903 -145 23937 -111
rect 23937 -145 23946 -111
rect 23894 -154 23946 -145
rect 24098 -111 24150 -102
rect 24098 -145 24107 -111
rect 24107 -145 24141 -111
rect 24141 -145 24150 -111
rect 24098 -154 24150 -145
rect 24302 -111 24354 -102
rect 24302 -145 24311 -111
rect 24311 -145 24345 -111
rect 24345 -145 24354 -111
rect 24302 -154 24354 -145
rect 24506 -111 24558 -102
rect 24506 -145 24515 -111
rect 24515 -145 24549 -111
rect 24549 -145 24558 -111
rect 24506 -154 24558 -145
rect 24710 -111 24762 -102
rect 24710 -145 24719 -111
rect 24719 -145 24753 -111
rect 24753 -145 24762 -111
rect 24710 -154 24762 -145
rect 24914 -111 24966 -102
rect 24914 -145 24923 -111
rect 24923 -145 24957 -111
rect 24957 -145 24966 -111
rect 24914 -154 24966 -145
rect 25118 -111 25170 -102
rect 25118 -145 25127 -111
rect 25127 -145 25161 -111
rect 25161 -145 25170 -111
rect 25118 -154 25170 -145
rect 25322 -111 25374 -102
rect 25322 -145 25331 -111
rect 25331 -145 25365 -111
rect 25365 -145 25374 -111
rect 25322 -154 25374 -145
rect 25526 -111 25578 -102
rect 25526 -145 25535 -111
rect 25535 -145 25569 -111
rect 25569 -145 25578 -111
rect 25526 -154 25578 -145
rect 25730 -111 25782 -102
rect 25730 -145 25739 -111
rect 25739 -145 25773 -111
rect 25773 -145 25782 -111
rect 25730 -154 25782 -145
rect 25934 -111 25986 -102
rect 25934 -145 25943 -111
rect 25943 -145 25977 -111
rect 25977 -145 25986 -111
rect 25934 -154 25986 -145
rect 26138 -111 26190 -102
rect 26138 -145 26147 -111
rect 26147 -145 26181 -111
rect 26181 -145 26190 -111
rect 26138 -154 26190 -145
rect 26342 -111 26394 -102
rect 26342 -145 26351 -111
rect 26351 -145 26385 -111
rect 26385 -145 26394 -111
rect 26342 -154 26394 -145
rect 26546 -111 26598 -102
rect 26546 -145 26555 -111
rect 26555 -145 26589 -111
rect 26589 -145 26598 -111
rect 26546 -154 26598 -145
rect 26750 -111 26802 -102
rect 26750 -145 26759 -111
rect 26759 -145 26793 -111
rect 26793 -145 26802 -111
rect 26750 -154 26802 -145
rect 26954 -111 27006 -102
rect 26954 -145 26963 -111
rect 26963 -145 26997 -111
rect 26997 -145 27006 -111
rect 26954 -154 27006 -145
rect 27158 -111 27210 -102
rect 27158 -145 27167 -111
rect 27167 -145 27201 -111
rect 27201 -145 27210 -111
rect 27158 -154 27210 -145
rect 27362 -111 27414 -102
rect 27362 -145 27371 -111
rect 27371 -145 27405 -111
rect 27405 -145 27414 -111
rect 27362 -154 27414 -145
rect 27566 -111 27618 -102
rect 27566 -145 27575 -111
rect 27575 -145 27609 -111
rect 27609 -145 27618 -111
rect 27566 -154 27618 -145
rect 27770 -111 27822 -102
rect 27770 -145 27779 -111
rect 27779 -145 27813 -111
rect 27813 -145 27822 -111
rect 27770 -154 27822 -145
rect 27974 -111 28026 -102
rect 27974 -145 27983 -111
rect 27983 -145 28017 -111
rect 28017 -145 28026 -111
rect 27974 -154 28026 -145
rect 28178 -111 28230 -102
rect 28178 -145 28187 -111
rect 28187 -145 28221 -111
rect 28221 -145 28230 -111
rect 28178 -154 28230 -145
rect 28382 -111 28434 -102
rect 28382 -145 28391 -111
rect 28391 -145 28425 -111
rect 28425 -145 28434 -111
rect 28382 -154 28434 -145
rect 28586 -111 28638 -102
rect 28586 -145 28595 -111
rect 28595 -145 28629 -111
rect 28629 -145 28638 -111
rect 28586 -154 28638 -145
rect 28790 -111 28842 -102
rect 28790 -145 28799 -111
rect 28799 -145 28833 -111
rect 28833 -145 28842 -111
rect 28790 -154 28842 -145
rect 28994 -111 29046 -102
rect 28994 -145 29003 -111
rect 29003 -145 29037 -111
rect 29037 -145 29046 -111
rect 28994 -154 29046 -145
rect 29198 -111 29250 -102
rect 29198 -145 29207 -111
rect 29207 -145 29241 -111
rect 29241 -145 29250 -111
rect 29198 -154 29250 -145
rect 29402 -111 29454 -102
rect 29402 -145 29411 -111
rect 29411 -145 29445 -111
rect 29445 -145 29454 -111
rect 29402 -154 29454 -145
rect 29606 -111 29658 -102
rect 29606 -145 29615 -111
rect 29615 -145 29649 -111
rect 29649 -145 29658 -111
rect 29606 -154 29658 -145
rect 29810 -111 29862 -102
rect 29810 -145 29819 -111
rect 29819 -145 29853 -111
rect 29853 -145 29862 -111
rect 29810 -154 29862 -145
rect 30014 -111 30066 -102
rect 30014 -145 30023 -111
rect 30023 -145 30057 -111
rect 30057 -145 30066 -111
rect 30014 -154 30066 -145
rect 30218 -111 30270 -102
rect 30218 -145 30227 -111
rect 30227 -145 30261 -111
rect 30261 -145 30270 -111
rect 30218 -154 30270 -145
rect 30422 -111 30474 -102
rect 30422 -145 30431 -111
rect 30431 -145 30465 -111
rect 30465 -145 30474 -111
rect 30422 -154 30474 -145
rect 30626 -111 30678 -102
rect 30626 -145 30635 -111
rect 30635 -145 30669 -111
rect 30669 -145 30678 -111
rect 30626 -154 30678 -145
rect 30830 -111 30882 -102
rect 30830 -145 30839 -111
rect 30839 -145 30873 -111
rect 30873 -145 30882 -111
rect 30830 -154 30882 -145
rect 31034 -111 31086 -102
rect 31034 -145 31043 -111
rect 31043 -145 31077 -111
rect 31077 -145 31086 -111
rect 31034 -154 31086 -145
rect 31238 -111 31290 -102
rect 31238 -145 31247 -111
rect 31247 -145 31281 -111
rect 31281 -145 31290 -111
rect 31238 -154 31290 -145
rect 31442 -111 31494 -102
rect 31442 -145 31451 -111
rect 31451 -145 31485 -111
rect 31485 -145 31494 -111
rect 31442 -154 31494 -145
rect 31646 -111 31698 -102
rect 31646 -145 31655 -111
rect 31655 -145 31689 -111
rect 31689 -145 31698 -111
rect 31646 -154 31698 -145
rect 31850 -111 31902 -102
rect 31850 -145 31859 -111
rect 31859 -145 31893 -111
rect 31893 -145 31902 -111
rect 31850 -154 31902 -145
rect 32054 -111 32106 -102
rect 32054 -145 32063 -111
rect 32063 -145 32097 -111
rect 32097 -145 32106 -111
rect 32054 -154 32106 -145
rect 32258 -111 32310 -102
rect 32258 -145 32267 -111
rect 32267 -145 32301 -111
rect 32301 -145 32310 -111
rect 32258 -154 32310 -145
rect 32462 -111 32514 -102
rect 32462 -145 32471 -111
rect 32471 -145 32505 -111
rect 32505 -145 32514 -111
rect 32462 -154 32514 -145
rect 32666 -111 32718 -102
rect 32666 -145 32675 -111
rect 32675 -145 32709 -111
rect 32709 -145 32718 -111
rect 32666 -154 32718 -145
rect 32870 -111 32922 -102
rect 32870 -145 32879 -111
rect 32879 -145 32913 -111
rect 32913 -145 32922 -111
rect 32870 -154 32922 -145
rect 33074 -111 33126 -102
rect 33074 -145 33083 -111
rect 33083 -145 33117 -111
rect 33117 -145 33126 -111
rect 33074 -154 33126 -145
rect 33278 -111 33330 -102
rect 33278 -145 33287 -111
rect 33287 -145 33321 -111
rect 33321 -145 33330 -111
rect 33278 -154 33330 -145
rect 33482 -111 33534 -102
rect 33482 -145 33491 -111
rect 33491 -145 33525 -111
rect 33525 -145 33534 -111
rect 33482 -154 33534 -145
rect 33686 -111 33738 -102
rect 33686 -145 33695 -111
rect 33695 -145 33729 -111
rect 33729 -145 33738 -111
rect 33686 -154 33738 -145
rect 33890 -111 33942 -102
rect 33890 -145 33899 -111
rect 33899 -145 33933 -111
rect 33933 -145 33942 -111
rect 33890 -154 33942 -145
rect 34094 -111 34146 -102
rect 34094 -145 34103 -111
rect 34103 -145 34137 -111
rect 34137 -145 34146 -111
rect 34094 -154 34146 -145
rect 34298 -111 34350 -102
rect 34298 -145 34307 -111
rect 34307 -145 34341 -111
rect 34341 -145 34350 -111
rect 34298 -154 34350 -145
rect 34502 -111 34554 -102
rect 34502 -145 34511 -111
rect 34511 -145 34545 -111
rect 34545 -145 34554 -111
rect 34502 -154 34554 -145
rect 34706 -111 34758 -102
rect 34706 -145 34715 -111
rect 34715 -145 34749 -111
rect 34749 -145 34758 -111
rect 34706 -154 34758 -145
rect 34910 -111 34962 -102
rect 34910 -145 34919 -111
rect 34919 -145 34953 -111
rect 34953 -145 34962 -111
rect 34910 -154 34962 -145
rect 35114 -111 35166 -102
rect 35114 -145 35123 -111
rect 35123 -145 35157 -111
rect 35157 -145 35166 -111
rect 35114 -154 35166 -145
rect 35318 -111 35370 -102
rect 35318 -145 35327 -111
rect 35327 -145 35361 -111
rect 35361 -145 35370 -111
rect 35318 -154 35370 -145
rect 35522 -111 35574 -102
rect 35522 -145 35531 -111
rect 35531 -145 35565 -111
rect 35565 -145 35574 -111
rect 35522 -154 35574 -145
rect 35726 -111 35778 -102
rect 35726 -145 35735 -111
rect 35735 -145 35769 -111
rect 35769 -145 35778 -111
rect 35726 -154 35778 -145
rect 35930 -111 35982 -102
rect 35930 -145 35939 -111
rect 35939 -145 35973 -111
rect 35973 -145 35982 -111
rect 35930 -154 35982 -145
rect 36134 -111 36186 -102
rect 36134 -145 36143 -111
rect 36143 -145 36177 -111
rect 36177 -145 36186 -111
rect 36134 -154 36186 -145
rect 36338 -111 36390 -102
rect 36338 -145 36347 -111
rect 36347 -145 36381 -111
rect 36381 -145 36390 -111
rect 36338 -154 36390 -145
rect 36542 -111 36594 -102
rect 36542 -145 36551 -111
rect 36551 -145 36585 -111
rect 36585 -145 36594 -111
rect 36542 -154 36594 -145
rect 36746 -111 36798 -102
rect 36746 -145 36755 -111
rect 36755 -145 36789 -111
rect 36789 -145 36798 -111
rect 36746 -154 36798 -145
rect 36950 -111 37002 -102
rect 36950 -145 36959 -111
rect 36959 -145 36993 -111
rect 36993 -145 37002 -111
rect 36950 -154 37002 -145
rect 37154 -111 37206 -102
rect 37154 -145 37163 -111
rect 37163 -145 37197 -111
rect 37197 -145 37206 -111
rect 37154 -154 37206 -145
rect 37358 -111 37410 -102
rect 37358 -145 37367 -111
rect 37367 -145 37401 -111
rect 37401 -145 37410 -111
rect 37358 -154 37410 -145
rect 37562 -111 37614 -102
rect 37562 -145 37571 -111
rect 37571 -145 37605 -111
rect 37605 -145 37614 -111
rect 37562 -154 37614 -145
rect 37766 -111 37818 -102
rect 37766 -145 37775 -111
rect 37775 -145 37809 -111
rect 37809 -145 37818 -111
rect 37766 -154 37818 -145
rect 37970 -111 38022 -102
rect 37970 -145 37979 -111
rect 37979 -145 38013 -111
rect 38013 -145 38022 -111
rect 37970 -154 38022 -145
rect 38174 -111 38226 -102
rect 38174 -145 38183 -111
rect 38183 -145 38217 -111
rect 38217 -145 38226 -111
rect 38174 -154 38226 -145
rect 38378 -111 38430 -102
rect 38378 -145 38387 -111
rect 38387 -145 38421 -111
rect 38421 -145 38430 -111
rect 38378 -154 38430 -145
rect 38582 -111 38634 -102
rect 38582 -145 38591 -111
rect 38591 -145 38625 -111
rect 38625 -145 38634 -111
rect 38582 -154 38634 -145
rect 38786 -111 38838 -102
rect 38786 -145 38795 -111
rect 38795 -145 38829 -111
rect 38829 -145 38838 -111
rect 38786 -154 38838 -145
rect 38990 -111 39042 -102
rect 38990 -145 38999 -111
rect 38999 -145 39033 -111
rect 39033 -145 39042 -111
rect 38990 -154 39042 -145
rect 39194 -111 39246 -102
rect 39194 -145 39203 -111
rect 39203 -145 39237 -111
rect 39237 -145 39246 -111
rect 39194 -154 39246 -145
rect 39398 -111 39450 -102
rect 39398 -145 39407 -111
rect 39407 -145 39441 -111
rect 39441 -145 39450 -111
rect 39398 -154 39450 -145
rect 39602 -111 39654 -102
rect 39602 -145 39611 -111
rect 39611 -145 39645 -111
rect 39645 -145 39654 -111
rect 39602 -154 39654 -145
rect 39806 -111 39858 -102
rect 39806 -145 39815 -111
rect 39815 -145 39849 -111
rect 39849 -145 39858 -111
rect 39806 -154 39858 -145
rect 40010 -111 40062 -102
rect 40010 -145 40019 -111
rect 40019 -145 40053 -111
rect 40053 -145 40062 -111
rect 40010 -154 40062 -145
rect 40214 -111 40266 -102
rect 40214 -145 40223 -111
rect 40223 -145 40257 -111
rect 40257 -145 40266 -111
rect 40214 -154 40266 -145
rect 40418 -111 40470 -102
rect 40418 -145 40427 -111
rect 40427 -145 40461 -111
rect 40461 -145 40470 -111
rect 40418 -154 40470 -145
rect 40622 -111 40674 -102
rect 40622 -145 40631 -111
rect 40631 -145 40665 -111
rect 40665 -145 40674 -111
rect 40622 -154 40674 -145
rect 40826 -111 40878 -102
rect 40826 -145 40835 -111
rect 40835 -145 40869 -111
rect 40869 -145 40878 -111
rect 40826 -154 40878 -145
rect 41030 -111 41082 -102
rect 41030 -145 41039 -111
rect 41039 -145 41073 -111
rect 41073 -145 41082 -111
rect 41030 -154 41082 -145
rect 41234 -111 41286 -102
rect 41234 -145 41243 -111
rect 41243 -145 41277 -111
rect 41277 -145 41286 -111
rect 41234 -154 41286 -145
rect 41438 -111 41490 -102
rect 41438 -145 41447 -111
rect 41447 -145 41481 -111
rect 41481 -145 41490 -111
rect 41438 -154 41490 -145
rect 41642 -111 41694 -102
rect 41642 -145 41651 -111
rect 41651 -145 41685 -111
rect 41685 -145 41694 -111
rect 41642 -154 41694 -145
rect 41846 -111 41898 -102
rect 41846 -145 41855 -111
rect 41855 -145 41889 -111
rect 41889 -145 41898 -111
rect 41846 -154 41898 -145
rect 42050 -111 42102 -102
rect 42050 -145 42059 -111
rect 42059 -145 42093 -111
rect 42093 -145 42102 -111
rect 42050 -154 42102 -145
rect 42254 -111 42306 -102
rect 42254 -145 42263 -111
rect 42263 -145 42297 -111
rect 42297 -145 42306 -111
rect 42254 -154 42306 -145
rect 42458 -111 42510 -102
rect 42458 -145 42467 -111
rect 42467 -145 42501 -111
rect 42501 -145 42510 -111
rect 42458 -154 42510 -145
rect 42662 -111 42714 -102
rect 42662 -145 42671 -111
rect 42671 -145 42705 -111
rect 42705 -145 42714 -111
rect 42662 -154 42714 -145
rect 42866 -111 42918 -102
rect 42866 -145 42875 -111
rect 42875 -145 42909 -111
rect 42909 -145 42918 -111
rect 42866 -154 42918 -145
rect 43070 -111 43122 -102
rect 43070 -145 43079 -111
rect 43079 -145 43113 -111
rect 43113 -145 43122 -111
rect 43070 -154 43122 -145
rect 43274 -111 43326 -102
rect 43274 -145 43283 -111
rect 43283 -145 43317 -111
rect 43317 -145 43326 -111
rect 43274 -154 43326 -145
rect 43478 -111 43530 -102
rect 43478 -145 43487 -111
rect 43487 -145 43521 -111
rect 43521 -145 43530 -111
rect 43478 -154 43530 -145
rect 43682 -111 43734 -102
rect 43682 -145 43691 -111
rect 43691 -145 43725 -111
rect 43725 -145 43734 -111
rect 43682 -154 43734 -145
rect 43886 -111 43938 -102
rect 43886 -145 43895 -111
rect 43895 -145 43929 -111
rect 43929 -145 43938 -111
rect 43886 -154 43938 -145
rect 44090 -111 44142 -102
rect 44090 -145 44099 -111
rect 44099 -145 44133 -111
rect 44133 -145 44142 -111
rect 44090 -154 44142 -145
rect 44294 -111 44346 -102
rect 44294 -145 44303 -111
rect 44303 -145 44337 -111
rect 44337 -145 44346 -111
rect 44294 -154 44346 -145
rect 44498 -111 44550 -102
rect 44498 -145 44507 -111
rect 44507 -145 44541 -111
rect 44541 -145 44550 -111
rect 44498 -154 44550 -145
rect 44702 -111 44754 -102
rect 44702 -145 44711 -111
rect 44711 -145 44745 -111
rect 44745 -145 44754 -111
rect 44702 -154 44754 -145
rect 44906 -111 44958 -102
rect 44906 -145 44915 -111
rect 44915 -145 44949 -111
rect 44949 -145 44958 -111
rect 44906 -154 44958 -145
rect 45110 -111 45162 -102
rect 45110 -145 45119 -111
rect 45119 -145 45153 -111
rect 45153 -145 45162 -111
rect 45110 -154 45162 -145
rect 45314 -111 45366 -102
rect 45314 -145 45323 -111
rect 45323 -145 45357 -111
rect 45357 -145 45366 -111
rect 45314 -154 45366 -145
rect 45518 -111 45570 -102
rect 45518 -145 45527 -111
rect 45527 -145 45561 -111
rect 45561 -145 45570 -111
rect 45518 -154 45570 -145
rect 45722 -111 45774 -102
rect 45722 -145 45731 -111
rect 45731 -145 45765 -111
rect 45765 -145 45774 -111
rect 45722 -154 45774 -145
rect 45926 -111 45978 -102
rect 45926 -145 45935 -111
rect 45935 -145 45969 -111
rect 45969 -145 45978 -111
rect 45926 -154 45978 -145
rect 46130 -111 46182 -102
rect 46130 -145 46139 -111
rect 46139 -145 46173 -111
rect 46173 -145 46182 -111
rect 46130 -154 46182 -145
rect 46334 -111 46386 -102
rect 46334 -145 46343 -111
rect 46343 -145 46377 -111
rect 46377 -145 46386 -111
rect 46334 -154 46386 -145
rect 46538 -111 46590 -102
rect 46538 -145 46547 -111
rect 46547 -145 46581 -111
rect 46581 -145 46590 -111
rect 46538 -154 46590 -145
rect 46742 -111 46794 -102
rect 46742 -145 46751 -111
rect 46751 -145 46785 -111
rect 46785 -145 46794 -111
rect 46742 -154 46794 -145
rect 46946 -111 46998 -102
rect 46946 -145 46955 -111
rect 46955 -145 46989 -111
rect 46989 -145 46998 -111
rect 46946 -154 46998 -145
rect 47150 -111 47202 -102
rect 47150 -145 47159 -111
rect 47159 -145 47193 -111
rect 47193 -145 47202 -111
rect 47150 -154 47202 -145
rect 47354 -111 47406 -102
rect 47354 -145 47363 -111
rect 47363 -145 47397 -111
rect 47397 -145 47406 -111
rect 47354 -154 47406 -145
rect 47558 -111 47610 -102
rect 47558 -145 47567 -111
rect 47567 -145 47601 -111
rect 47601 -145 47610 -111
rect 47558 -154 47610 -145
rect 47762 -111 47814 -102
rect 47762 -145 47771 -111
rect 47771 -145 47805 -111
rect 47805 -145 47814 -111
rect 47762 -154 47814 -145
rect 47966 -111 48018 -102
rect 47966 -145 47975 -111
rect 47975 -145 48009 -111
rect 48009 -145 48018 -111
rect 47966 -154 48018 -145
rect 48170 -111 48222 -102
rect 48170 -145 48179 -111
rect 48179 -145 48213 -111
rect 48213 -145 48222 -111
rect 48170 -154 48222 -145
rect 48374 -111 48426 -102
rect 48374 -145 48383 -111
rect 48383 -145 48417 -111
rect 48417 -145 48426 -111
rect 48374 -154 48426 -145
rect 48578 -111 48630 -102
rect 48578 -145 48587 -111
rect 48587 -145 48621 -111
rect 48621 -145 48630 -111
rect 48578 -154 48630 -145
rect 48782 -111 48834 -102
rect 48782 -145 48791 -111
rect 48791 -145 48825 -111
rect 48825 -145 48834 -111
rect 48782 -154 48834 -145
rect 48986 -111 49038 -102
rect 48986 -145 48995 -111
rect 48995 -145 49029 -111
rect 49029 -145 49038 -111
rect 48986 -154 49038 -145
rect 49190 -111 49242 -102
rect 49190 -145 49199 -111
rect 49199 -145 49233 -111
rect 49233 -145 49242 -111
rect 49190 -154 49242 -145
rect 49394 -111 49446 -102
rect 49394 -145 49403 -111
rect 49403 -145 49437 -111
rect 49437 -145 49446 -111
rect 49394 -154 49446 -145
rect 49598 -111 49650 -102
rect 49598 -145 49607 -111
rect 49607 -145 49641 -111
rect 49641 -145 49650 -111
rect 49598 -154 49650 -145
rect 49802 -111 49854 -102
rect 49802 -145 49811 -111
rect 49811 -145 49845 -111
rect 49845 -145 49854 -111
rect 49802 -154 49854 -145
rect 50006 -111 50058 -102
rect 50006 -145 50015 -111
rect 50015 -145 50049 -111
rect 50049 -145 50058 -111
rect 50006 -154 50058 -145
rect 50210 -111 50262 -102
rect 50210 -145 50219 -111
rect 50219 -145 50253 -111
rect 50253 -145 50262 -111
rect 50210 -154 50262 -145
rect 50414 -111 50466 -102
rect 50414 -145 50423 -111
rect 50423 -145 50457 -111
rect 50457 -145 50466 -111
rect 50414 -154 50466 -145
rect 50618 -111 50670 -102
rect 50618 -145 50627 -111
rect 50627 -145 50661 -111
rect 50661 -145 50670 -111
rect 50618 -154 50670 -145
rect 50822 -111 50874 -102
rect 50822 -145 50831 -111
rect 50831 -145 50865 -111
rect 50865 -145 50874 -111
rect 50822 -154 50874 -145
rect 51026 -111 51078 -102
rect 51026 -145 51035 -111
rect 51035 -145 51069 -111
rect 51069 -145 51078 -111
rect 51026 -154 51078 -145
rect 51230 -111 51282 -102
rect 51230 -145 51239 -111
rect 51239 -145 51273 -111
rect 51273 -145 51282 -111
rect 51230 -154 51282 -145
rect 51434 -111 51486 -102
rect 51434 -145 51443 -111
rect 51443 -145 51477 -111
rect 51477 -145 51486 -111
rect 51434 -154 51486 -145
rect 51638 -111 51690 -102
rect 51638 -145 51647 -111
rect 51647 -145 51681 -111
rect 51681 -145 51690 -111
rect 51638 -154 51690 -145
rect 51842 -111 51894 -102
rect 51842 -145 51851 -111
rect 51851 -145 51885 -111
rect 51885 -145 51894 -111
rect 51842 -154 51894 -145
rect 52046 -111 52098 -102
rect 52046 -145 52055 -111
rect 52055 -145 52089 -111
rect 52089 -145 52098 -111
rect 52046 -154 52098 -145
<< metal2 >>
rect 61 240 52313 268
rect 12 -102 52250 -96
rect 12 -154 26 -102
rect 78 -154 230 -102
rect 282 -154 434 -102
rect 486 -154 638 -102
rect 690 -154 842 -102
rect 894 -154 1046 -102
rect 1098 -154 1250 -102
rect 1302 -154 1454 -102
rect 1506 -154 1658 -102
rect 1710 -154 1862 -102
rect 1914 -154 2066 -102
rect 2118 -154 2270 -102
rect 2322 -154 2474 -102
rect 2526 -154 2678 -102
rect 2730 -154 2882 -102
rect 2934 -154 3086 -102
rect 3138 -154 3290 -102
rect 3342 -154 3494 -102
rect 3546 -154 3698 -102
rect 3750 -154 3902 -102
rect 3954 -154 4106 -102
rect 4158 -154 4310 -102
rect 4362 -154 4514 -102
rect 4566 -154 4718 -102
rect 4770 -154 4922 -102
rect 4974 -154 5126 -102
rect 5178 -154 5330 -102
rect 5382 -154 5534 -102
rect 5586 -154 5738 -102
rect 5790 -154 5942 -102
rect 5994 -154 6146 -102
rect 6198 -154 6350 -102
rect 6402 -154 6554 -102
rect 6606 -154 6758 -102
rect 6810 -154 6962 -102
rect 7014 -154 7166 -102
rect 7218 -154 7370 -102
rect 7422 -154 7574 -102
rect 7626 -154 7778 -102
rect 7830 -154 7982 -102
rect 8034 -154 8186 -102
rect 8238 -154 8390 -102
rect 8442 -154 8594 -102
rect 8646 -154 8798 -102
rect 8850 -154 9002 -102
rect 9054 -154 9206 -102
rect 9258 -154 9410 -102
rect 9462 -154 9614 -102
rect 9666 -154 9818 -102
rect 9870 -154 10022 -102
rect 10074 -154 10226 -102
rect 10278 -154 10430 -102
rect 10482 -154 10634 -102
rect 10686 -154 10838 -102
rect 10890 -154 11042 -102
rect 11094 -154 11246 -102
rect 11298 -154 11450 -102
rect 11502 -154 11654 -102
rect 11706 -154 11858 -102
rect 11910 -154 12062 -102
rect 12114 -154 12266 -102
rect 12318 -154 12470 -102
rect 12522 -154 12674 -102
rect 12726 -154 12878 -102
rect 12930 -154 13082 -102
rect 13134 -154 13286 -102
rect 13338 -154 13490 -102
rect 13542 -154 13694 -102
rect 13746 -154 13898 -102
rect 13950 -154 14102 -102
rect 14154 -154 14306 -102
rect 14358 -154 14510 -102
rect 14562 -154 14714 -102
rect 14766 -154 14918 -102
rect 14970 -154 15122 -102
rect 15174 -154 15326 -102
rect 15378 -154 15530 -102
rect 15582 -154 15734 -102
rect 15786 -154 15938 -102
rect 15990 -154 16142 -102
rect 16194 -154 16346 -102
rect 16398 -154 16550 -102
rect 16602 -154 16754 -102
rect 16806 -154 16958 -102
rect 17010 -154 17162 -102
rect 17214 -154 17366 -102
rect 17418 -154 17570 -102
rect 17622 -154 17774 -102
rect 17826 -154 17978 -102
rect 18030 -154 18182 -102
rect 18234 -154 18386 -102
rect 18438 -154 18590 -102
rect 18642 -154 18794 -102
rect 18846 -154 18998 -102
rect 19050 -154 19202 -102
rect 19254 -154 19406 -102
rect 19458 -154 19610 -102
rect 19662 -154 19814 -102
rect 19866 -154 20018 -102
rect 20070 -154 20222 -102
rect 20274 -154 20426 -102
rect 20478 -154 20630 -102
rect 20682 -154 20834 -102
rect 20886 -154 21038 -102
rect 21090 -154 21242 -102
rect 21294 -154 21446 -102
rect 21498 -154 21650 -102
rect 21702 -154 21854 -102
rect 21906 -154 22058 -102
rect 22110 -154 22262 -102
rect 22314 -154 22466 -102
rect 22518 -154 22670 -102
rect 22722 -154 22874 -102
rect 22926 -154 23078 -102
rect 23130 -154 23282 -102
rect 23334 -154 23486 -102
rect 23538 -154 23690 -102
rect 23742 -154 23894 -102
rect 23946 -154 24098 -102
rect 24150 -154 24302 -102
rect 24354 -154 24506 -102
rect 24558 -154 24710 -102
rect 24762 -154 24914 -102
rect 24966 -154 25118 -102
rect 25170 -154 25322 -102
rect 25374 -154 25526 -102
rect 25578 -154 25730 -102
rect 25782 -154 25934 -102
rect 25986 -154 26138 -102
rect 26190 -154 26342 -102
rect 26394 -154 26546 -102
rect 26598 -154 26750 -102
rect 26802 -154 26954 -102
rect 27006 -154 27158 -102
rect 27210 -154 27362 -102
rect 27414 -154 27566 -102
rect 27618 -154 27770 -102
rect 27822 -154 27974 -102
rect 28026 -154 28178 -102
rect 28230 -154 28382 -102
rect 28434 -154 28586 -102
rect 28638 -154 28790 -102
rect 28842 -154 28994 -102
rect 29046 -154 29198 -102
rect 29250 -154 29402 -102
rect 29454 -154 29606 -102
rect 29658 -154 29810 -102
rect 29862 -154 30014 -102
rect 30066 -154 30218 -102
rect 30270 -154 30422 -102
rect 30474 -154 30626 -102
rect 30678 -154 30830 -102
rect 30882 -154 31034 -102
rect 31086 -154 31238 -102
rect 31290 -154 31442 -102
rect 31494 -154 31646 -102
rect 31698 -154 31850 -102
rect 31902 -154 32054 -102
rect 32106 -154 32258 -102
rect 32310 -154 32462 -102
rect 32514 -154 32666 -102
rect 32718 -154 32870 -102
rect 32922 -154 33074 -102
rect 33126 -154 33278 -102
rect 33330 -154 33482 -102
rect 33534 -154 33686 -102
rect 33738 -154 33890 -102
rect 33942 -154 34094 -102
rect 34146 -154 34298 -102
rect 34350 -154 34502 -102
rect 34554 -154 34706 -102
rect 34758 -154 34910 -102
rect 34962 -154 35114 -102
rect 35166 -154 35318 -102
rect 35370 -154 35522 -102
rect 35574 -154 35726 -102
rect 35778 -154 35930 -102
rect 35982 -154 36134 -102
rect 36186 -154 36338 -102
rect 36390 -154 36542 -102
rect 36594 -154 36746 -102
rect 36798 -154 36950 -102
rect 37002 -154 37154 -102
rect 37206 -154 37358 -102
rect 37410 -154 37562 -102
rect 37614 -154 37766 -102
rect 37818 -154 37970 -102
rect 38022 -154 38174 -102
rect 38226 -154 38378 -102
rect 38430 -154 38582 -102
rect 38634 -154 38786 -102
rect 38838 -154 38990 -102
rect 39042 -154 39194 -102
rect 39246 -154 39398 -102
rect 39450 -154 39602 -102
rect 39654 -154 39806 -102
rect 39858 -154 40010 -102
rect 40062 -154 40214 -102
rect 40266 -154 40418 -102
rect 40470 -154 40622 -102
rect 40674 -154 40826 -102
rect 40878 -154 41030 -102
rect 41082 -154 41234 -102
rect 41286 -154 41438 -102
rect 41490 -154 41642 -102
rect 41694 -154 41846 -102
rect 41898 -154 42050 -102
rect 42102 -154 42254 -102
rect 42306 -154 42458 -102
rect 42510 -154 42662 -102
rect 42714 -154 42866 -102
rect 42918 -154 43070 -102
rect 43122 -154 43274 -102
rect 43326 -154 43478 -102
rect 43530 -154 43682 -102
rect 43734 -154 43886 -102
rect 43938 -154 44090 -102
rect 44142 -154 44294 -102
rect 44346 -154 44498 -102
rect 44550 -154 44702 -102
rect 44754 -154 44906 -102
rect 44958 -154 45110 -102
rect 45162 -154 45314 -102
rect 45366 -154 45518 -102
rect 45570 -154 45722 -102
rect 45774 -154 45926 -102
rect 45978 -154 46130 -102
rect 46182 -154 46334 -102
rect 46386 -154 46538 -102
rect 46590 -154 46742 -102
rect 46794 -154 46946 -102
rect 46998 -154 47150 -102
rect 47202 -154 47354 -102
rect 47406 -154 47558 -102
rect 47610 -154 47762 -102
rect 47814 -154 47966 -102
rect 48018 -154 48170 -102
rect 48222 -154 48374 -102
rect 48426 -154 48578 -102
rect 48630 -154 48782 -102
rect 48834 -154 48986 -102
rect 49038 -154 49190 -102
rect 49242 -154 49394 -102
rect 49446 -154 49598 -102
rect 49650 -154 49802 -102
rect 49854 -154 50006 -102
rect 50058 -154 50210 -102
rect 50262 -154 50414 -102
rect 50466 -154 50618 -102
rect 50670 -154 50822 -102
rect 50874 -154 51026 -102
rect 51078 -154 51230 -102
rect 51282 -154 51434 -102
rect 51486 -154 51638 -102
rect 51690 -154 51842 -102
rect 51894 -154 52046 -102
rect 52098 -154 52250 -102
rect 12 -160 52250 -154
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_0
timestamp 1581449086
transform 1 0 52020 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_1
timestamp 1581449086
transform 1 0 51816 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_2
timestamp 1581449086
transform 1 0 51612 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_3
timestamp 1581449086
transform 1 0 51408 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_4
timestamp 1581449086
transform 1 0 51204 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_5
timestamp 1581449086
transform 1 0 51000 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_6
timestamp 1581449086
transform 1 0 50796 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_7
timestamp 1581449086
transform 1 0 50592 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_8
timestamp 1581449086
transform 1 0 50388 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_9
timestamp 1581449086
transform 1 0 50184 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_10
timestamp 1581449086
transform 1 0 49980 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_11
timestamp 1581449086
transform 1 0 49776 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_12
timestamp 1581449086
transform 1 0 49572 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_13
timestamp 1581449086
transform 1 0 49368 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_14
timestamp 1581449086
transform 1 0 49164 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_15
timestamp 1581449086
transform 1 0 48960 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_16
timestamp 1581449086
transform 1 0 48756 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_17
timestamp 1581449086
transform 1 0 48552 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_18
timestamp 1581449086
transform 1 0 48348 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_19
timestamp 1581449086
transform 1 0 48144 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_20
timestamp 1581449086
transform 1 0 47940 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_21
timestamp 1581449086
transform 1 0 47736 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_22
timestamp 1581449086
transform 1 0 47532 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_23
timestamp 1581449086
transform 1 0 47328 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_24
timestamp 1581449086
transform 1 0 47124 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_25
timestamp 1581449086
transform 1 0 46920 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_26
timestamp 1581449086
transform 1 0 46716 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_27
timestamp 1581449086
transform 1 0 46512 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_28
timestamp 1581449086
transform 1 0 46308 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_29
timestamp 1581449086
transform 1 0 46104 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_30
timestamp 1581449086
transform 1 0 45900 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_31
timestamp 1581449086
transform 1 0 45696 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_32
timestamp 1581449086
transform 1 0 45492 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_33
timestamp 1581449086
transform 1 0 45288 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_34
timestamp 1581449086
transform 1 0 45084 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_35
timestamp 1581449086
transform 1 0 44880 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_36
timestamp 1581449086
transform 1 0 44676 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_37
timestamp 1581449086
transform 1 0 44472 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_38
timestamp 1581449086
transform 1 0 44268 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_39
timestamp 1581449086
transform 1 0 44064 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_40
timestamp 1581449086
transform 1 0 43860 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_41
timestamp 1581449086
transform 1 0 43656 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_42
timestamp 1581449086
transform 1 0 43452 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_43
timestamp 1581449086
transform 1 0 43248 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_44
timestamp 1581449086
transform 1 0 43044 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_45
timestamp 1581449086
transform 1 0 42840 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_46
timestamp 1581449086
transform 1 0 42636 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_47
timestamp 1581449086
transform 1 0 42432 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_48
timestamp 1581449086
transform 1 0 42228 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_49
timestamp 1581449086
transform 1 0 42024 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_50
timestamp 1581449086
transform 1 0 41820 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_51
timestamp 1581449086
transform 1 0 41616 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_52
timestamp 1581449086
transform 1 0 41412 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_53
timestamp 1581449086
transform 1 0 41208 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_54
timestamp 1581449086
transform 1 0 41004 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_55
timestamp 1581449086
transform 1 0 40800 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_56
timestamp 1581449086
transform 1 0 40596 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_57
timestamp 1581449086
transform 1 0 40392 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_58
timestamp 1581449086
transform 1 0 40188 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_59
timestamp 1581449086
transform 1 0 39984 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_60
timestamp 1581449086
transform 1 0 39780 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_61
timestamp 1581449086
transform 1 0 39576 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_62
timestamp 1581449086
transform 1 0 39372 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_63
timestamp 1581449086
transform 1 0 39168 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_64
timestamp 1581449086
transform 1 0 38964 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_65
timestamp 1581449086
transform 1 0 38760 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_66
timestamp 1581449086
transform 1 0 38556 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_67
timestamp 1581449086
transform 1 0 38352 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_68
timestamp 1581449086
transform 1 0 38148 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_69
timestamp 1581449086
transform 1 0 37944 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_70
timestamp 1581449086
transform 1 0 37740 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_71
timestamp 1581449086
transform 1 0 37536 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_72
timestamp 1581449086
transform 1 0 37332 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_73
timestamp 1581449086
transform 1 0 37128 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_74
timestamp 1581449086
transform 1 0 36924 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_75
timestamp 1581449086
transform 1 0 36720 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_76
timestamp 1581449086
transform 1 0 36516 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_77
timestamp 1581449086
transform 1 0 36312 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_78
timestamp 1581449086
transform 1 0 36108 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_79
timestamp 1581449086
transform 1 0 35904 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_80
timestamp 1581449086
transform 1 0 35700 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_81
timestamp 1581449086
transform 1 0 35496 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_82
timestamp 1581449086
transform 1 0 35292 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_83
timestamp 1581449086
transform 1 0 35088 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_84
timestamp 1581449086
transform 1 0 34884 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_85
timestamp 1581449086
transform 1 0 34680 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_86
timestamp 1581449086
transform 1 0 34476 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_87
timestamp 1581449086
transform 1 0 34272 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_88
timestamp 1581449086
transform 1 0 34068 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_89
timestamp 1581449086
transform 1 0 33864 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_90
timestamp 1581449086
transform 1 0 33660 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_91
timestamp 1581449086
transform 1 0 33456 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_92
timestamp 1581449086
transform 1 0 33252 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_93
timestamp 1581449086
transform 1 0 33048 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_94
timestamp 1581449086
transform 1 0 32844 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_95
timestamp 1581449086
transform 1 0 32640 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_96
timestamp 1581449086
transform 1 0 32436 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_97
timestamp 1581449086
transform 1 0 32232 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_98
timestamp 1581449086
transform 1 0 32028 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_99
timestamp 1581449086
transform 1 0 31824 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_100
timestamp 1581449086
transform 1 0 31620 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_101
timestamp 1581449086
transform 1 0 31416 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_102
timestamp 1581449086
transform 1 0 31212 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_103
timestamp 1581449086
transform 1 0 31008 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_104
timestamp 1581449086
transform 1 0 30804 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_105
timestamp 1581449086
transform 1 0 30600 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_106
timestamp 1581449086
transform 1 0 30396 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_107
timestamp 1581449086
transform 1 0 30192 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_108
timestamp 1581449086
transform 1 0 29988 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_109
timestamp 1581449086
transform 1 0 29784 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_110
timestamp 1581449086
transform 1 0 29580 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_111
timestamp 1581449086
transform 1 0 29376 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_112
timestamp 1581449086
transform 1 0 29172 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_113
timestamp 1581449086
transform 1 0 28968 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_114
timestamp 1581449086
transform 1 0 28764 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_115
timestamp 1581449086
transform 1 0 28560 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_116
timestamp 1581449086
transform 1 0 28356 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_117
timestamp 1581449086
transform 1 0 28152 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_118
timestamp 1581449086
transform 1 0 27948 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_119
timestamp 1581449086
transform 1 0 27744 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_120
timestamp 1581449086
transform 1 0 27540 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_121
timestamp 1581449086
transform 1 0 27336 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_122
timestamp 1581449086
transform 1 0 27132 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_123
timestamp 1581449086
transform 1 0 26928 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_124
timestamp 1581449086
transform 1 0 26724 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_125
timestamp 1581449086
transform 1 0 26520 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_126
timestamp 1581449086
transform 1 0 26316 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_127
timestamp 1581449086
transform 1 0 26112 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_128
timestamp 1581449086
transform 1 0 25908 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_129
timestamp 1581449086
transform 1 0 25704 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_130
timestamp 1581449086
transform 1 0 25500 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_131
timestamp 1581449086
transform 1 0 25296 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_132
timestamp 1581449086
transform 1 0 25092 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_133
timestamp 1581449086
transform 1 0 24888 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_134
timestamp 1581449086
transform 1 0 24684 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_135
timestamp 1581449086
transform 1 0 24480 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_136
timestamp 1581449086
transform 1 0 24276 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_137
timestamp 1581449086
transform 1 0 24072 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_138
timestamp 1581449086
transform 1 0 23868 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_139
timestamp 1581449086
transform 1 0 23664 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_140
timestamp 1581449086
transform 1 0 23460 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_141
timestamp 1581449086
transform 1 0 23256 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_142
timestamp 1581449086
transform 1 0 23052 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_143
timestamp 1581449086
transform 1 0 22848 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_144
timestamp 1581449086
transform 1 0 22644 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_145
timestamp 1581449086
transform 1 0 22440 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_146
timestamp 1581449086
transform 1 0 22236 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_147
timestamp 1581449086
transform 1 0 22032 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_148
timestamp 1581449086
transform 1 0 21828 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_149
timestamp 1581449086
transform 1 0 21624 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_150
timestamp 1581449086
transform 1 0 21420 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_151
timestamp 1581449086
transform 1 0 21216 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_152
timestamp 1581449086
transform 1 0 21012 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_153
timestamp 1581449086
transform 1 0 20808 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_154
timestamp 1581449086
transform 1 0 20604 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_155
timestamp 1581449086
transform 1 0 20400 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_156
timestamp 1581449086
transform 1 0 20196 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_157
timestamp 1581449086
transform 1 0 19992 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_158
timestamp 1581449086
transform 1 0 19788 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_159
timestamp 1581449086
transform 1 0 19584 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_160
timestamp 1581449086
transform 1 0 19380 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_161
timestamp 1581449086
transform 1 0 19176 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_162
timestamp 1581449086
transform 1 0 18972 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_163
timestamp 1581449086
transform 1 0 18768 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_164
timestamp 1581449086
transform 1 0 18564 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_165
timestamp 1581449086
transform 1 0 18360 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_166
timestamp 1581449086
transform 1 0 18156 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_167
timestamp 1581449086
transform 1 0 17952 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_168
timestamp 1581449086
transform 1 0 17748 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_169
timestamp 1581449086
transform 1 0 17544 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_170
timestamp 1581449086
transform 1 0 17340 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_171
timestamp 1581449086
transform 1 0 17136 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_172
timestamp 1581449086
transform 1 0 16932 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_173
timestamp 1581449086
transform 1 0 16728 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_174
timestamp 1581449086
transform 1 0 16524 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_175
timestamp 1581449086
transform 1 0 16320 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_176
timestamp 1581449086
transform 1 0 16116 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_177
timestamp 1581449086
transform 1 0 15912 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_178
timestamp 1581449086
transform 1 0 15708 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_179
timestamp 1581449086
transform 1 0 15504 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_180
timestamp 1581449086
transform 1 0 15300 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_181
timestamp 1581449086
transform 1 0 15096 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_182
timestamp 1581449086
transform 1 0 14892 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_183
timestamp 1581449086
transform 1 0 14688 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_184
timestamp 1581449086
transform 1 0 14484 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_185
timestamp 1581449086
transform 1 0 14280 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_186
timestamp 1581449086
transform 1 0 14076 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_187
timestamp 1581449086
transform 1 0 13872 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_188
timestamp 1581449086
transform 1 0 13668 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_189
timestamp 1581449086
transform 1 0 13464 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_190
timestamp 1581449086
transform 1 0 13260 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_191
timestamp 1581449086
transform 1 0 13056 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_192
timestamp 1581449086
transform 1 0 12852 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_193
timestamp 1581449086
transform 1 0 12648 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_194
timestamp 1581449086
transform 1 0 12444 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_195
timestamp 1581449086
transform 1 0 12240 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_196
timestamp 1581449086
transform 1 0 12036 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_197
timestamp 1581449086
transform 1 0 11832 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_198
timestamp 1581449086
transform 1 0 11628 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_199
timestamp 1581449086
transform 1 0 11424 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_200
timestamp 1581449086
transform 1 0 11220 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_201
timestamp 1581449086
transform 1 0 11016 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_202
timestamp 1581449086
transform 1 0 10812 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_203
timestamp 1581449086
transform 1 0 10608 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_204
timestamp 1581449086
transform 1 0 10404 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_205
timestamp 1581449086
transform 1 0 10200 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_206
timestamp 1581449086
transform 1 0 9996 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_207
timestamp 1581449086
transform 1 0 9792 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_208
timestamp 1581449086
transform 1 0 9588 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_209
timestamp 1581449086
transform 1 0 9384 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_210
timestamp 1581449086
transform 1 0 9180 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_211
timestamp 1581449086
transform 1 0 8976 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_212
timestamp 1581449086
transform 1 0 8772 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_213
timestamp 1581449086
transform 1 0 8568 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_214
timestamp 1581449086
transform 1 0 8364 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_215
timestamp 1581449086
transform 1 0 8160 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_216
timestamp 1581449086
transform 1 0 7956 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_217
timestamp 1581449086
transform 1 0 7752 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_218
timestamp 1581449086
transform 1 0 7548 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_219
timestamp 1581449086
transform 1 0 7344 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_220
timestamp 1581449086
transform 1 0 7140 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_221
timestamp 1581449086
transform 1 0 6936 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_222
timestamp 1581449086
transform 1 0 6732 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_223
timestamp 1581449086
transform 1 0 6528 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_224
timestamp 1581449086
transform 1 0 6324 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_225
timestamp 1581449086
transform 1 0 6120 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_226
timestamp 1581449086
transform 1 0 5916 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_227
timestamp 1581449086
transform 1 0 5712 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_228
timestamp 1581449086
transform 1 0 5508 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_229
timestamp 1581449086
transform 1 0 5304 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_230
timestamp 1581449086
transform 1 0 5100 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_231
timestamp 1581449086
transform 1 0 4896 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_232
timestamp 1581449086
transform 1 0 4692 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_233
timestamp 1581449086
transform 1 0 4488 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_234
timestamp 1581449086
transform 1 0 4284 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_235
timestamp 1581449086
transform 1 0 4080 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_236
timestamp 1581449086
transform 1 0 3876 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_237
timestamp 1581449086
transform 1 0 3672 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_238
timestamp 1581449086
transform 1 0 3468 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_239
timestamp 1581449086
transform 1 0 3264 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_240
timestamp 1581449086
transform 1 0 3060 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_241
timestamp 1581449086
transform 1 0 2856 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_242
timestamp 1581449086
transform 1 0 2652 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_243
timestamp 1581449086
transform 1 0 2448 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_244
timestamp 1581449086
transform 1 0 2244 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_245
timestamp 1581449086
transform 1 0 2040 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_246
timestamp 1581449086
transform 1 0 1836 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_247
timestamp 1581449086
transform 1 0 1632 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_248
timestamp 1581449086
transform 1 0 1428 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_249
timestamp 1581449086
transform 1 0 1224 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_250
timestamp 1581449086
transform 1 0 1020 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_251
timestamp 1581449086
transform 1 0 816 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_252
timestamp 1581449086
transform 1 0 612 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_253
timestamp 1581449086
transform 1 0 408 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_254
timestamp 1581449086
transform 1 0 204 0 1 0
box 0 -212 232 184
use sky130_rom_krom_precharge_cell  sky130_rom_krom_precharge_cell_255
timestamp 1581449086
transform 1 0 0 0 1 0
box 0 -212 232 184
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_0
timestamp 1581449086
transform 1 0 52266 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_1
timestamp 1581449086
transform 1 0 50634 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_2
timestamp 1581449086
transform 1 0 49002 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_3
timestamp 1581449086
transform 1 0 47370 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_4
timestamp 1581449086
transform 1 0 45738 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_5
timestamp 1581449086
transform 1 0 44106 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_6
timestamp 1581449086
transform 1 0 42474 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_7
timestamp 1581449086
transform 1 0 40842 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_8
timestamp 1581449086
transform 1 0 39210 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_9
timestamp 1581449086
transform 1 0 37578 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_10
timestamp 1581449086
transform 1 0 35946 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_11
timestamp 1581449086
transform 1 0 34314 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_12
timestamp 1581449086
transform 1 0 32682 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_13
timestamp 1581449086
transform 1 0 31050 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_14
timestamp 1581449086
transform 1 0 29418 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_15
timestamp 1581449086
transform 1 0 27786 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_16
timestamp 1581449086
transform 1 0 26154 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_17
timestamp 1581449086
transform 1 0 24522 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_18
timestamp 1581449086
transform 1 0 22890 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_19
timestamp 1581449086
transform 1 0 21258 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_20
timestamp 1581449086
transform 1 0 19626 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_21
timestamp 1581449086
transform 1 0 17994 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_22
timestamp 1581449086
transform 1 0 16362 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_23
timestamp 1581449086
transform 1 0 14730 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_24
timestamp 1581449086
transform 1 0 13098 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_25
timestamp 1581449086
transform 1 0 11466 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_26
timestamp 1581449086
transform 1 0 9834 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_27
timestamp 1581449086
transform 1 0 8202 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_28
timestamp 1581449086
transform 1 0 6570 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_29
timestamp 1581449086
transform 1 0 4938 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_30
timestamp 1581449086
transform 1 0 3306 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_31
timestamp 1581449086
transform 1 0 1674 0 1 204
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_0  sky130_rom_krom_rom_poly_tap_0_32
timestamp 1581449086
transform 1 0 42 0 1 204
box 0 17 66 83
<< labels >>
rlabel nwell s 52332 408 52332 408 4 upper right
rlabel metal2 s 61 240 89 268 4 gate
port 3 nsew
rlabel metal2 s 52285 240 52313 268 4 precharge_r
port 5 nsew
rlabel metal1 s 122 86 150 114 4 pre_bl0_out
port 7 nsew
rlabel metal1 s 326 86 354 114 4 pre_bl1_out
port 9 nsew
rlabel metal1 s 530 86 558 114 4 pre_bl2_out
port 11 nsew
rlabel metal1 s 734 86 762 114 4 pre_bl3_out
port 13 nsew
rlabel metal1 s 938 86 966 114 4 pre_bl4_out
port 15 nsew
rlabel metal1 s 1142 86 1170 114 4 pre_bl5_out
port 17 nsew
rlabel metal1 s 1346 86 1374 114 4 pre_bl6_out
port 19 nsew
rlabel metal1 s 1550 86 1578 114 4 pre_bl7_out
port 21 nsew
rlabel metal1 s 1754 86 1782 114 4 pre_bl8_out
port 23 nsew
rlabel metal1 s 1958 86 1986 114 4 pre_bl9_out
port 25 nsew
rlabel metal1 s 2162 86 2190 114 4 pre_bl10_out
port 27 nsew
rlabel metal1 s 2366 86 2394 114 4 pre_bl11_out
port 29 nsew
rlabel metal1 s 2570 86 2598 114 4 pre_bl12_out
port 31 nsew
rlabel metal1 s 2774 86 2802 114 4 pre_bl13_out
port 33 nsew
rlabel metal1 s 2978 86 3006 114 4 pre_bl14_out
port 35 nsew
rlabel metal1 s 3182 86 3210 114 4 pre_bl15_out
port 37 nsew
rlabel metal1 s 3386 86 3414 114 4 pre_bl16_out
port 39 nsew
rlabel metal1 s 3590 86 3618 114 4 pre_bl17_out
port 41 nsew
rlabel metal1 s 3794 86 3822 114 4 pre_bl18_out
port 43 nsew
rlabel metal1 s 3998 86 4026 114 4 pre_bl19_out
port 45 nsew
rlabel metal1 s 4202 86 4230 114 4 pre_bl20_out
port 47 nsew
rlabel metal1 s 4406 86 4434 114 4 pre_bl21_out
port 49 nsew
rlabel metal1 s 4610 86 4638 114 4 pre_bl22_out
port 51 nsew
rlabel metal1 s 4814 86 4842 114 4 pre_bl23_out
port 53 nsew
rlabel metal1 s 5018 86 5046 114 4 pre_bl24_out
port 55 nsew
rlabel metal1 s 5222 86 5250 114 4 pre_bl25_out
port 57 nsew
rlabel metal1 s 5426 86 5454 114 4 pre_bl26_out
port 59 nsew
rlabel metal1 s 5630 86 5658 114 4 pre_bl27_out
port 61 nsew
rlabel metal1 s 5834 86 5862 114 4 pre_bl28_out
port 63 nsew
rlabel metal1 s 6038 86 6066 114 4 pre_bl29_out
port 65 nsew
rlabel metal1 s 6242 86 6270 114 4 pre_bl30_out
port 67 nsew
rlabel metal1 s 6446 86 6474 114 4 pre_bl31_out
port 69 nsew
rlabel metal1 s 6650 86 6678 114 4 pre_bl32_out
port 71 nsew
rlabel metal1 s 6854 86 6882 114 4 pre_bl33_out
port 73 nsew
rlabel metal1 s 7058 86 7086 114 4 pre_bl34_out
port 75 nsew
rlabel metal1 s 7262 86 7290 114 4 pre_bl35_out
port 77 nsew
rlabel metal1 s 7466 86 7494 114 4 pre_bl36_out
port 79 nsew
rlabel metal1 s 7670 86 7698 114 4 pre_bl37_out
port 81 nsew
rlabel metal1 s 7874 86 7902 114 4 pre_bl38_out
port 83 nsew
rlabel metal1 s 8078 86 8106 114 4 pre_bl39_out
port 85 nsew
rlabel metal1 s 8282 86 8310 114 4 pre_bl40_out
port 87 nsew
rlabel metal1 s 8486 86 8514 114 4 pre_bl41_out
port 89 nsew
rlabel metal1 s 8690 86 8718 114 4 pre_bl42_out
port 91 nsew
rlabel metal1 s 8894 86 8922 114 4 pre_bl43_out
port 93 nsew
rlabel metal1 s 9098 86 9126 114 4 pre_bl44_out
port 95 nsew
rlabel metal1 s 9302 86 9330 114 4 pre_bl45_out
port 97 nsew
rlabel metal1 s 9506 86 9534 114 4 pre_bl46_out
port 99 nsew
rlabel metal1 s 9710 86 9738 114 4 pre_bl47_out
port 101 nsew
rlabel metal1 s 9914 86 9942 114 4 pre_bl48_out
port 103 nsew
rlabel metal1 s 10118 86 10146 114 4 pre_bl49_out
port 105 nsew
rlabel metal1 s 10322 86 10350 114 4 pre_bl50_out
port 107 nsew
rlabel metal1 s 10526 86 10554 114 4 pre_bl51_out
port 109 nsew
rlabel metal1 s 10730 86 10758 114 4 pre_bl52_out
port 111 nsew
rlabel metal1 s 10934 86 10962 114 4 pre_bl53_out
port 113 nsew
rlabel metal1 s 11138 86 11166 114 4 pre_bl54_out
port 115 nsew
rlabel metal1 s 11342 86 11370 114 4 pre_bl55_out
port 117 nsew
rlabel metal1 s 11546 86 11574 114 4 pre_bl56_out
port 119 nsew
rlabel metal1 s 11750 86 11778 114 4 pre_bl57_out
port 121 nsew
rlabel metal1 s 11954 86 11982 114 4 pre_bl58_out
port 123 nsew
rlabel metal1 s 12158 86 12186 114 4 pre_bl59_out
port 125 nsew
rlabel metal1 s 12362 86 12390 114 4 pre_bl60_out
port 127 nsew
rlabel metal1 s 12566 86 12594 114 4 pre_bl61_out
port 129 nsew
rlabel metal1 s 12770 86 12798 114 4 pre_bl62_out
port 131 nsew
rlabel metal1 s 12974 86 13002 114 4 pre_bl63_out
port 133 nsew
rlabel metal1 s 13178 86 13206 114 4 pre_bl64_out
port 135 nsew
rlabel metal1 s 13382 86 13410 114 4 pre_bl65_out
port 137 nsew
rlabel metal1 s 13586 86 13614 114 4 pre_bl66_out
port 139 nsew
rlabel metal1 s 13790 86 13818 114 4 pre_bl67_out
port 141 nsew
rlabel metal1 s 13994 86 14022 114 4 pre_bl68_out
port 143 nsew
rlabel metal1 s 14198 86 14226 114 4 pre_bl69_out
port 145 nsew
rlabel metal1 s 14402 86 14430 114 4 pre_bl70_out
port 147 nsew
rlabel metal1 s 14606 86 14634 114 4 pre_bl71_out
port 149 nsew
rlabel metal1 s 14810 86 14838 114 4 pre_bl72_out
port 151 nsew
rlabel metal1 s 15014 86 15042 114 4 pre_bl73_out
port 153 nsew
rlabel metal1 s 15218 86 15246 114 4 pre_bl74_out
port 155 nsew
rlabel metal1 s 15422 86 15450 114 4 pre_bl75_out
port 157 nsew
rlabel metal1 s 15626 86 15654 114 4 pre_bl76_out
port 159 nsew
rlabel metal1 s 15830 86 15858 114 4 pre_bl77_out
port 161 nsew
rlabel metal1 s 16034 86 16062 114 4 pre_bl78_out
port 163 nsew
rlabel metal1 s 16238 86 16266 114 4 pre_bl79_out
port 165 nsew
rlabel metal1 s 16442 86 16470 114 4 pre_bl80_out
port 167 nsew
rlabel metal1 s 16646 86 16674 114 4 pre_bl81_out
port 169 nsew
rlabel metal1 s 16850 86 16878 114 4 pre_bl82_out
port 171 nsew
rlabel metal1 s 17054 86 17082 114 4 pre_bl83_out
port 173 nsew
rlabel metal1 s 17258 86 17286 114 4 pre_bl84_out
port 175 nsew
rlabel metal1 s 17462 86 17490 114 4 pre_bl85_out
port 177 nsew
rlabel metal1 s 17666 86 17694 114 4 pre_bl86_out
port 179 nsew
rlabel metal1 s 17870 86 17898 114 4 pre_bl87_out
port 181 nsew
rlabel metal1 s 18074 86 18102 114 4 pre_bl88_out
port 183 nsew
rlabel metal1 s 18278 86 18306 114 4 pre_bl89_out
port 185 nsew
rlabel metal1 s 18482 86 18510 114 4 pre_bl90_out
port 187 nsew
rlabel metal1 s 18686 86 18714 114 4 pre_bl91_out
port 189 nsew
rlabel metal1 s 18890 86 18918 114 4 pre_bl92_out
port 191 nsew
rlabel metal1 s 19094 86 19122 114 4 pre_bl93_out
port 193 nsew
rlabel metal1 s 19298 86 19326 114 4 pre_bl94_out
port 195 nsew
rlabel metal1 s 19502 86 19530 114 4 pre_bl95_out
port 197 nsew
rlabel metal1 s 19706 86 19734 114 4 pre_bl96_out
port 199 nsew
rlabel metal1 s 19910 86 19938 114 4 pre_bl97_out
port 201 nsew
rlabel metal1 s 20114 86 20142 114 4 pre_bl98_out
port 203 nsew
rlabel metal1 s 20318 86 20346 114 4 pre_bl99_out
port 205 nsew
rlabel metal1 s 20522 86 20550 114 4 pre_bl100_out
port 207 nsew
rlabel metal1 s 20726 86 20754 114 4 pre_bl101_out
port 209 nsew
rlabel metal1 s 20930 86 20958 114 4 pre_bl102_out
port 211 nsew
rlabel metal1 s 21134 86 21162 114 4 pre_bl103_out
port 213 nsew
rlabel metal1 s 21338 86 21366 114 4 pre_bl104_out
port 215 nsew
rlabel metal1 s 21542 86 21570 114 4 pre_bl105_out
port 217 nsew
rlabel metal1 s 21746 86 21774 114 4 pre_bl106_out
port 219 nsew
rlabel metal1 s 21950 86 21978 114 4 pre_bl107_out
port 221 nsew
rlabel metal1 s 22154 86 22182 114 4 pre_bl108_out
port 223 nsew
rlabel metal1 s 22358 86 22386 114 4 pre_bl109_out
port 225 nsew
rlabel metal1 s 22562 86 22590 114 4 pre_bl110_out
port 227 nsew
rlabel metal1 s 22766 86 22794 114 4 pre_bl111_out
port 229 nsew
rlabel metal1 s 22970 86 22998 114 4 pre_bl112_out
port 231 nsew
rlabel metal1 s 23174 86 23202 114 4 pre_bl113_out
port 233 nsew
rlabel metal1 s 23378 86 23406 114 4 pre_bl114_out
port 235 nsew
rlabel metal1 s 23582 86 23610 114 4 pre_bl115_out
port 237 nsew
rlabel metal1 s 23786 86 23814 114 4 pre_bl116_out
port 239 nsew
rlabel metal1 s 23990 86 24018 114 4 pre_bl117_out
port 241 nsew
rlabel metal1 s 24194 86 24222 114 4 pre_bl118_out
port 243 nsew
rlabel metal1 s 24398 86 24426 114 4 pre_bl119_out
port 245 nsew
rlabel metal1 s 24602 86 24630 114 4 pre_bl120_out
port 247 nsew
rlabel metal1 s 24806 86 24834 114 4 pre_bl121_out
port 249 nsew
rlabel metal1 s 25010 86 25038 114 4 pre_bl122_out
port 251 nsew
rlabel metal1 s 25214 86 25242 114 4 pre_bl123_out
port 253 nsew
rlabel metal1 s 25418 86 25446 114 4 pre_bl124_out
port 255 nsew
rlabel metal1 s 25622 86 25650 114 4 pre_bl125_out
port 257 nsew
rlabel metal1 s 25826 86 25854 114 4 pre_bl126_out
port 259 nsew
rlabel metal1 s 26030 86 26058 114 4 pre_bl127_out
port 261 nsew
rlabel metal1 s 26234 86 26262 114 4 pre_bl128_out
port 263 nsew
rlabel metal1 s 26438 86 26466 114 4 pre_bl129_out
port 265 nsew
rlabel metal1 s 26642 86 26670 114 4 pre_bl130_out
port 267 nsew
rlabel metal1 s 26846 86 26874 114 4 pre_bl131_out
port 269 nsew
rlabel metal1 s 27050 86 27078 114 4 pre_bl132_out
port 271 nsew
rlabel metal1 s 27254 86 27282 114 4 pre_bl133_out
port 273 nsew
rlabel metal1 s 27458 86 27486 114 4 pre_bl134_out
port 275 nsew
rlabel metal1 s 27662 86 27690 114 4 pre_bl135_out
port 277 nsew
rlabel metal1 s 27866 86 27894 114 4 pre_bl136_out
port 279 nsew
rlabel metal1 s 28070 86 28098 114 4 pre_bl137_out
port 281 nsew
rlabel metal1 s 28274 86 28302 114 4 pre_bl138_out
port 283 nsew
rlabel metal1 s 28478 86 28506 114 4 pre_bl139_out
port 285 nsew
rlabel metal1 s 28682 86 28710 114 4 pre_bl140_out
port 287 nsew
rlabel metal1 s 28886 86 28914 114 4 pre_bl141_out
port 289 nsew
rlabel metal1 s 29090 86 29118 114 4 pre_bl142_out
port 291 nsew
rlabel metal1 s 29294 86 29322 114 4 pre_bl143_out
port 293 nsew
rlabel metal1 s 29498 86 29526 114 4 pre_bl144_out
port 295 nsew
rlabel metal1 s 29702 86 29730 114 4 pre_bl145_out
port 297 nsew
rlabel metal1 s 29906 86 29934 114 4 pre_bl146_out
port 299 nsew
rlabel metal1 s 30110 86 30138 114 4 pre_bl147_out
port 301 nsew
rlabel metal1 s 30314 86 30342 114 4 pre_bl148_out
port 303 nsew
rlabel metal1 s 30518 86 30546 114 4 pre_bl149_out
port 305 nsew
rlabel metal1 s 30722 86 30750 114 4 pre_bl150_out
port 307 nsew
rlabel metal1 s 30926 86 30954 114 4 pre_bl151_out
port 309 nsew
rlabel metal1 s 31130 86 31158 114 4 pre_bl152_out
port 311 nsew
rlabel metal1 s 31334 86 31362 114 4 pre_bl153_out
port 313 nsew
rlabel metal1 s 31538 86 31566 114 4 pre_bl154_out
port 315 nsew
rlabel metal1 s 31742 86 31770 114 4 pre_bl155_out
port 317 nsew
rlabel metal1 s 31946 86 31974 114 4 pre_bl156_out
port 319 nsew
rlabel metal1 s 32150 86 32178 114 4 pre_bl157_out
port 321 nsew
rlabel metal1 s 32354 86 32382 114 4 pre_bl158_out
port 323 nsew
rlabel metal1 s 32558 86 32586 114 4 pre_bl159_out
port 325 nsew
rlabel metal1 s 32762 86 32790 114 4 pre_bl160_out
port 327 nsew
rlabel metal1 s 32966 86 32994 114 4 pre_bl161_out
port 329 nsew
rlabel metal1 s 33170 86 33198 114 4 pre_bl162_out
port 331 nsew
rlabel metal1 s 33374 86 33402 114 4 pre_bl163_out
port 333 nsew
rlabel metal1 s 33578 86 33606 114 4 pre_bl164_out
port 335 nsew
rlabel metal1 s 33782 86 33810 114 4 pre_bl165_out
port 337 nsew
rlabel metal1 s 33986 86 34014 114 4 pre_bl166_out
port 339 nsew
rlabel metal1 s 34190 86 34218 114 4 pre_bl167_out
port 341 nsew
rlabel metal1 s 34394 86 34422 114 4 pre_bl168_out
port 343 nsew
rlabel metal1 s 34598 86 34626 114 4 pre_bl169_out
port 345 nsew
rlabel metal1 s 34802 86 34830 114 4 pre_bl170_out
port 347 nsew
rlabel metal1 s 35006 86 35034 114 4 pre_bl171_out
port 349 nsew
rlabel metal1 s 35210 86 35238 114 4 pre_bl172_out
port 351 nsew
rlabel metal1 s 35414 86 35442 114 4 pre_bl173_out
port 353 nsew
rlabel metal1 s 35618 86 35646 114 4 pre_bl174_out
port 355 nsew
rlabel metal1 s 35822 86 35850 114 4 pre_bl175_out
port 357 nsew
rlabel metal1 s 36026 86 36054 114 4 pre_bl176_out
port 359 nsew
rlabel metal1 s 36230 86 36258 114 4 pre_bl177_out
port 361 nsew
rlabel metal1 s 36434 86 36462 114 4 pre_bl178_out
port 363 nsew
rlabel metal1 s 36638 86 36666 114 4 pre_bl179_out
port 365 nsew
rlabel metal1 s 36842 86 36870 114 4 pre_bl180_out
port 367 nsew
rlabel metal1 s 37046 86 37074 114 4 pre_bl181_out
port 369 nsew
rlabel metal1 s 37250 86 37278 114 4 pre_bl182_out
port 371 nsew
rlabel metal1 s 37454 86 37482 114 4 pre_bl183_out
port 373 nsew
rlabel metal1 s 37658 86 37686 114 4 pre_bl184_out
port 375 nsew
rlabel metal1 s 37862 86 37890 114 4 pre_bl185_out
port 377 nsew
rlabel metal1 s 38066 86 38094 114 4 pre_bl186_out
port 379 nsew
rlabel metal1 s 38270 86 38298 114 4 pre_bl187_out
port 381 nsew
rlabel metal1 s 38474 86 38502 114 4 pre_bl188_out
port 383 nsew
rlabel metal1 s 38678 86 38706 114 4 pre_bl189_out
port 385 nsew
rlabel metal1 s 38882 86 38910 114 4 pre_bl190_out
port 387 nsew
rlabel metal1 s 39086 86 39114 114 4 pre_bl191_out
port 389 nsew
rlabel metal1 s 39290 86 39318 114 4 pre_bl192_out
port 391 nsew
rlabel metal1 s 39494 86 39522 114 4 pre_bl193_out
port 393 nsew
rlabel metal1 s 39698 86 39726 114 4 pre_bl194_out
port 395 nsew
rlabel metal1 s 39902 86 39930 114 4 pre_bl195_out
port 397 nsew
rlabel metal1 s 40106 86 40134 114 4 pre_bl196_out
port 399 nsew
rlabel metal1 s 40310 86 40338 114 4 pre_bl197_out
port 401 nsew
rlabel metal1 s 40514 86 40542 114 4 pre_bl198_out
port 403 nsew
rlabel metal1 s 40718 86 40746 114 4 pre_bl199_out
port 405 nsew
rlabel metal1 s 40922 86 40950 114 4 pre_bl200_out
port 407 nsew
rlabel metal1 s 41126 86 41154 114 4 pre_bl201_out
port 409 nsew
rlabel metal1 s 41330 86 41358 114 4 pre_bl202_out
port 411 nsew
rlabel metal1 s 41534 86 41562 114 4 pre_bl203_out
port 413 nsew
rlabel metal1 s 41738 86 41766 114 4 pre_bl204_out
port 415 nsew
rlabel metal1 s 41942 86 41970 114 4 pre_bl205_out
port 417 nsew
rlabel metal1 s 42146 86 42174 114 4 pre_bl206_out
port 419 nsew
rlabel metal1 s 42350 86 42378 114 4 pre_bl207_out
port 421 nsew
rlabel metal1 s 42554 86 42582 114 4 pre_bl208_out
port 423 nsew
rlabel metal1 s 42758 86 42786 114 4 pre_bl209_out
port 425 nsew
rlabel metal1 s 42962 86 42990 114 4 pre_bl210_out
port 427 nsew
rlabel metal1 s 43166 86 43194 114 4 pre_bl211_out
port 429 nsew
rlabel metal1 s 43370 86 43398 114 4 pre_bl212_out
port 431 nsew
rlabel metal1 s 43574 86 43602 114 4 pre_bl213_out
port 433 nsew
rlabel metal1 s 43778 86 43806 114 4 pre_bl214_out
port 435 nsew
rlabel metal1 s 43982 86 44010 114 4 pre_bl215_out
port 437 nsew
rlabel metal1 s 44186 86 44214 114 4 pre_bl216_out
port 439 nsew
rlabel metal1 s 44390 86 44418 114 4 pre_bl217_out
port 441 nsew
rlabel metal1 s 44594 86 44622 114 4 pre_bl218_out
port 443 nsew
rlabel metal1 s 44798 86 44826 114 4 pre_bl219_out
port 445 nsew
rlabel metal1 s 45002 86 45030 114 4 pre_bl220_out
port 447 nsew
rlabel metal1 s 45206 86 45234 114 4 pre_bl221_out
port 449 nsew
rlabel metal1 s 45410 86 45438 114 4 pre_bl222_out
port 451 nsew
rlabel metal1 s 45614 86 45642 114 4 pre_bl223_out
port 453 nsew
rlabel metal1 s 45818 86 45846 114 4 pre_bl224_out
port 455 nsew
rlabel metal1 s 46022 86 46050 114 4 pre_bl225_out
port 457 nsew
rlabel metal1 s 46226 86 46254 114 4 pre_bl226_out
port 459 nsew
rlabel metal1 s 46430 86 46458 114 4 pre_bl227_out
port 461 nsew
rlabel metal1 s 46634 86 46662 114 4 pre_bl228_out
port 463 nsew
rlabel metal1 s 46838 86 46866 114 4 pre_bl229_out
port 465 nsew
rlabel metal1 s 47042 86 47070 114 4 pre_bl230_out
port 467 nsew
rlabel metal1 s 47246 86 47274 114 4 pre_bl231_out
port 469 nsew
rlabel metal1 s 47450 86 47478 114 4 pre_bl232_out
port 471 nsew
rlabel metal1 s 47654 86 47682 114 4 pre_bl233_out
port 473 nsew
rlabel metal1 s 47858 86 47886 114 4 pre_bl234_out
port 475 nsew
rlabel metal1 s 48062 86 48090 114 4 pre_bl235_out
port 477 nsew
rlabel metal1 s 48266 86 48294 114 4 pre_bl236_out
port 479 nsew
rlabel metal1 s 48470 86 48498 114 4 pre_bl237_out
port 481 nsew
rlabel metal1 s 48674 86 48702 114 4 pre_bl238_out
port 483 nsew
rlabel metal1 s 48878 86 48906 114 4 pre_bl239_out
port 485 nsew
rlabel metal1 s 49082 86 49110 114 4 pre_bl240_out
port 487 nsew
rlabel metal1 s 49286 86 49314 114 4 pre_bl241_out
port 489 nsew
rlabel metal1 s 49490 86 49518 114 4 pre_bl242_out
port 491 nsew
rlabel metal1 s 49694 86 49722 114 4 pre_bl243_out
port 493 nsew
rlabel metal1 s 49898 86 49926 114 4 pre_bl244_out
port 495 nsew
rlabel metal1 s 50102 86 50130 114 4 pre_bl245_out
port 497 nsew
rlabel metal1 s 50306 86 50334 114 4 pre_bl246_out
port 499 nsew
rlabel metal1 s 50510 86 50538 114 4 pre_bl247_out
port 501 nsew
rlabel metal1 s 50714 86 50742 114 4 pre_bl248_out
port 503 nsew
rlabel metal1 s 50918 86 50946 114 4 pre_bl249_out
port 505 nsew
rlabel metal1 s 51122 86 51150 114 4 pre_bl250_out
port 507 nsew
rlabel metal1 s 51326 86 51354 114 4 pre_bl251_out
port 509 nsew
rlabel metal1 s 51530 86 51558 114 4 pre_bl252_out
port 511 nsew
rlabel metal1 s 51734 86 51762 114 4 pre_bl253_out
port 513 nsew
rlabel metal1 s 51938 86 51966 114 4 pre_bl254_out
port 515 nsew
rlabel metal1 s 52142 86 52170 114 4 pre_bl255_out
port 517 nsew
rlabel metal2 s 12 -160 40 -96 4 vdd
port 519 nsew
<< properties >>
string FIXED_BBOX 52043 -161 52101 -160
<< end >>
