magic
tech sky130A
magscale 1 2
timestamp 1581320205
<< checkpaint >>
rect -1260 -1344 14565 9281
<< pwell >>
rect 177 6030 13177 6132
rect 177 4294 13177 4396
rect 177 2558 13177 2660
rect 177 822 13177 924
<< psubdiff >>
rect 203 6098 285 6106
rect 203 6064 227 6098
rect 261 6064 285 6098
rect 203 6056 285 6064
rect 407 6098 489 6106
rect 407 6064 431 6098
rect 465 6064 489 6098
rect 407 6056 489 6064
rect 611 6098 693 6106
rect 611 6064 635 6098
rect 669 6064 693 6098
rect 611 6056 693 6064
rect 815 6098 897 6106
rect 815 6064 839 6098
rect 873 6064 897 6098
rect 815 6056 897 6064
rect 1019 6098 1101 6106
rect 1019 6064 1043 6098
rect 1077 6064 1101 6098
rect 1019 6056 1101 6064
rect 1223 6098 1305 6106
rect 1223 6064 1247 6098
rect 1281 6064 1305 6098
rect 1223 6056 1305 6064
rect 1427 6098 1509 6106
rect 1427 6064 1451 6098
rect 1485 6064 1509 6098
rect 1427 6056 1509 6064
rect 1631 6098 1713 6106
rect 1631 6064 1655 6098
rect 1689 6064 1713 6098
rect 1631 6056 1713 6064
rect 1835 6098 1917 6106
rect 1835 6064 1859 6098
rect 1893 6064 1917 6098
rect 1835 6056 1917 6064
rect 2039 6098 2121 6106
rect 2039 6064 2063 6098
rect 2097 6064 2121 6098
rect 2039 6056 2121 6064
rect 2243 6098 2325 6106
rect 2243 6064 2267 6098
rect 2301 6064 2325 6098
rect 2243 6056 2325 6064
rect 2447 6098 2529 6106
rect 2447 6064 2471 6098
rect 2505 6064 2529 6098
rect 2447 6056 2529 6064
rect 2651 6098 2733 6106
rect 2651 6064 2675 6098
rect 2709 6064 2733 6098
rect 2651 6056 2733 6064
rect 2855 6098 2937 6106
rect 2855 6064 2879 6098
rect 2913 6064 2937 6098
rect 2855 6056 2937 6064
rect 3059 6098 3141 6106
rect 3059 6064 3083 6098
rect 3117 6064 3141 6098
rect 3059 6056 3141 6064
rect 3263 6098 3345 6106
rect 3263 6064 3287 6098
rect 3321 6064 3345 6098
rect 3263 6056 3345 6064
rect 3467 6098 3549 6106
rect 3467 6064 3491 6098
rect 3525 6064 3549 6098
rect 3467 6056 3549 6064
rect 3671 6098 3753 6106
rect 3671 6064 3695 6098
rect 3729 6064 3753 6098
rect 3671 6056 3753 6064
rect 3875 6098 3957 6106
rect 3875 6064 3899 6098
rect 3933 6064 3957 6098
rect 3875 6056 3957 6064
rect 4079 6098 4161 6106
rect 4079 6064 4103 6098
rect 4137 6064 4161 6098
rect 4079 6056 4161 6064
rect 4283 6098 4365 6106
rect 4283 6064 4307 6098
rect 4341 6064 4365 6098
rect 4283 6056 4365 6064
rect 4487 6098 4569 6106
rect 4487 6064 4511 6098
rect 4545 6064 4569 6098
rect 4487 6056 4569 6064
rect 4691 6098 4773 6106
rect 4691 6064 4715 6098
rect 4749 6064 4773 6098
rect 4691 6056 4773 6064
rect 4895 6098 4977 6106
rect 4895 6064 4919 6098
rect 4953 6064 4977 6098
rect 4895 6056 4977 6064
rect 5099 6098 5181 6106
rect 5099 6064 5123 6098
rect 5157 6064 5181 6098
rect 5099 6056 5181 6064
rect 5303 6098 5385 6106
rect 5303 6064 5327 6098
rect 5361 6064 5385 6098
rect 5303 6056 5385 6064
rect 5507 6098 5589 6106
rect 5507 6064 5531 6098
rect 5565 6064 5589 6098
rect 5507 6056 5589 6064
rect 5711 6098 5793 6106
rect 5711 6064 5735 6098
rect 5769 6064 5793 6098
rect 5711 6056 5793 6064
rect 5915 6098 5997 6106
rect 5915 6064 5939 6098
rect 5973 6064 5997 6098
rect 5915 6056 5997 6064
rect 6119 6098 6201 6106
rect 6119 6064 6143 6098
rect 6177 6064 6201 6098
rect 6119 6056 6201 6064
rect 6323 6098 6405 6106
rect 6323 6064 6347 6098
rect 6381 6064 6405 6098
rect 6323 6056 6405 6064
rect 6527 6098 6609 6106
rect 6527 6064 6551 6098
rect 6585 6064 6609 6098
rect 6527 6056 6609 6064
rect 6731 6098 6813 6106
rect 6731 6064 6755 6098
rect 6789 6064 6813 6098
rect 6731 6056 6813 6064
rect 6935 6098 7017 6106
rect 6935 6064 6959 6098
rect 6993 6064 7017 6098
rect 6935 6056 7017 6064
rect 7139 6098 7221 6106
rect 7139 6064 7163 6098
rect 7197 6064 7221 6098
rect 7139 6056 7221 6064
rect 7343 6098 7425 6106
rect 7343 6064 7367 6098
rect 7401 6064 7425 6098
rect 7343 6056 7425 6064
rect 7547 6098 7629 6106
rect 7547 6064 7571 6098
rect 7605 6064 7629 6098
rect 7547 6056 7629 6064
rect 7751 6098 7833 6106
rect 7751 6064 7775 6098
rect 7809 6064 7833 6098
rect 7751 6056 7833 6064
rect 7955 6098 8037 6106
rect 7955 6064 7979 6098
rect 8013 6064 8037 6098
rect 7955 6056 8037 6064
rect 8159 6098 8241 6106
rect 8159 6064 8183 6098
rect 8217 6064 8241 6098
rect 8159 6056 8241 6064
rect 8363 6098 8445 6106
rect 8363 6064 8387 6098
rect 8421 6064 8445 6098
rect 8363 6056 8445 6064
rect 8567 6098 8649 6106
rect 8567 6064 8591 6098
rect 8625 6064 8649 6098
rect 8567 6056 8649 6064
rect 8771 6098 8853 6106
rect 8771 6064 8795 6098
rect 8829 6064 8853 6098
rect 8771 6056 8853 6064
rect 8975 6098 9057 6106
rect 8975 6064 8999 6098
rect 9033 6064 9057 6098
rect 8975 6056 9057 6064
rect 9179 6098 9261 6106
rect 9179 6064 9203 6098
rect 9237 6064 9261 6098
rect 9179 6056 9261 6064
rect 9383 6098 9465 6106
rect 9383 6064 9407 6098
rect 9441 6064 9465 6098
rect 9383 6056 9465 6064
rect 9587 6098 9669 6106
rect 9587 6064 9611 6098
rect 9645 6064 9669 6098
rect 9587 6056 9669 6064
rect 9791 6098 9873 6106
rect 9791 6064 9815 6098
rect 9849 6064 9873 6098
rect 9791 6056 9873 6064
rect 9995 6098 10077 6106
rect 9995 6064 10019 6098
rect 10053 6064 10077 6098
rect 9995 6056 10077 6064
rect 10199 6098 10281 6106
rect 10199 6064 10223 6098
rect 10257 6064 10281 6098
rect 10199 6056 10281 6064
rect 10403 6098 10485 6106
rect 10403 6064 10427 6098
rect 10461 6064 10485 6098
rect 10403 6056 10485 6064
rect 10607 6098 10689 6106
rect 10607 6064 10631 6098
rect 10665 6064 10689 6098
rect 10607 6056 10689 6064
rect 10811 6098 10893 6106
rect 10811 6064 10835 6098
rect 10869 6064 10893 6098
rect 10811 6056 10893 6064
rect 11015 6098 11097 6106
rect 11015 6064 11039 6098
rect 11073 6064 11097 6098
rect 11015 6056 11097 6064
rect 11219 6098 11301 6106
rect 11219 6064 11243 6098
rect 11277 6064 11301 6098
rect 11219 6056 11301 6064
rect 11423 6098 11505 6106
rect 11423 6064 11447 6098
rect 11481 6064 11505 6098
rect 11423 6056 11505 6064
rect 11627 6098 11709 6106
rect 11627 6064 11651 6098
rect 11685 6064 11709 6098
rect 11627 6056 11709 6064
rect 11831 6098 11913 6106
rect 11831 6064 11855 6098
rect 11889 6064 11913 6098
rect 11831 6056 11913 6064
rect 12035 6098 12117 6106
rect 12035 6064 12059 6098
rect 12093 6064 12117 6098
rect 12035 6056 12117 6064
rect 12239 6098 12321 6106
rect 12239 6064 12263 6098
rect 12297 6064 12321 6098
rect 12239 6056 12321 6064
rect 12443 6098 12525 6106
rect 12443 6064 12467 6098
rect 12501 6064 12525 6098
rect 12443 6056 12525 6064
rect 12647 6098 12729 6106
rect 12647 6064 12671 6098
rect 12705 6064 12729 6098
rect 12647 6056 12729 6064
rect 12851 6098 12933 6106
rect 12851 6064 12875 6098
rect 12909 6064 12933 6098
rect 12851 6056 12933 6064
rect 13069 6098 13151 6106
rect 13069 6064 13093 6098
rect 13127 6064 13151 6098
rect 13069 6056 13151 6064
rect 203 4362 285 4370
rect 203 4328 227 4362
rect 261 4328 285 4362
rect 203 4320 285 4328
rect 407 4362 489 4370
rect 407 4328 431 4362
rect 465 4328 489 4362
rect 407 4320 489 4328
rect 611 4362 693 4370
rect 611 4328 635 4362
rect 669 4328 693 4362
rect 611 4320 693 4328
rect 815 4362 897 4370
rect 815 4328 839 4362
rect 873 4328 897 4362
rect 815 4320 897 4328
rect 1019 4362 1101 4370
rect 1019 4328 1043 4362
rect 1077 4328 1101 4362
rect 1019 4320 1101 4328
rect 1223 4362 1305 4370
rect 1223 4328 1247 4362
rect 1281 4328 1305 4362
rect 1223 4320 1305 4328
rect 1427 4362 1509 4370
rect 1427 4328 1451 4362
rect 1485 4328 1509 4362
rect 1427 4320 1509 4328
rect 1631 4362 1713 4370
rect 1631 4328 1655 4362
rect 1689 4328 1713 4362
rect 1631 4320 1713 4328
rect 1835 4362 1917 4370
rect 1835 4328 1859 4362
rect 1893 4328 1917 4362
rect 1835 4320 1917 4328
rect 2039 4362 2121 4370
rect 2039 4328 2063 4362
rect 2097 4328 2121 4362
rect 2039 4320 2121 4328
rect 2243 4362 2325 4370
rect 2243 4328 2267 4362
rect 2301 4328 2325 4362
rect 2243 4320 2325 4328
rect 2447 4362 2529 4370
rect 2447 4328 2471 4362
rect 2505 4328 2529 4362
rect 2447 4320 2529 4328
rect 2651 4362 2733 4370
rect 2651 4328 2675 4362
rect 2709 4328 2733 4362
rect 2651 4320 2733 4328
rect 2855 4362 2937 4370
rect 2855 4328 2879 4362
rect 2913 4328 2937 4362
rect 2855 4320 2937 4328
rect 3059 4362 3141 4370
rect 3059 4328 3083 4362
rect 3117 4328 3141 4362
rect 3059 4320 3141 4328
rect 3263 4362 3345 4370
rect 3263 4328 3287 4362
rect 3321 4328 3345 4362
rect 3263 4320 3345 4328
rect 3467 4362 3549 4370
rect 3467 4328 3491 4362
rect 3525 4328 3549 4362
rect 3467 4320 3549 4328
rect 3671 4362 3753 4370
rect 3671 4328 3695 4362
rect 3729 4328 3753 4362
rect 3671 4320 3753 4328
rect 3875 4362 3957 4370
rect 3875 4328 3899 4362
rect 3933 4328 3957 4362
rect 3875 4320 3957 4328
rect 4079 4362 4161 4370
rect 4079 4328 4103 4362
rect 4137 4328 4161 4362
rect 4079 4320 4161 4328
rect 4283 4362 4365 4370
rect 4283 4328 4307 4362
rect 4341 4328 4365 4362
rect 4283 4320 4365 4328
rect 4487 4362 4569 4370
rect 4487 4328 4511 4362
rect 4545 4328 4569 4362
rect 4487 4320 4569 4328
rect 4691 4362 4773 4370
rect 4691 4328 4715 4362
rect 4749 4328 4773 4362
rect 4691 4320 4773 4328
rect 4895 4362 4977 4370
rect 4895 4328 4919 4362
rect 4953 4328 4977 4362
rect 4895 4320 4977 4328
rect 5099 4362 5181 4370
rect 5099 4328 5123 4362
rect 5157 4328 5181 4362
rect 5099 4320 5181 4328
rect 5303 4362 5385 4370
rect 5303 4328 5327 4362
rect 5361 4328 5385 4362
rect 5303 4320 5385 4328
rect 5507 4362 5589 4370
rect 5507 4328 5531 4362
rect 5565 4328 5589 4362
rect 5507 4320 5589 4328
rect 5711 4362 5793 4370
rect 5711 4328 5735 4362
rect 5769 4328 5793 4362
rect 5711 4320 5793 4328
rect 5915 4362 5997 4370
rect 5915 4328 5939 4362
rect 5973 4328 5997 4362
rect 5915 4320 5997 4328
rect 6119 4362 6201 4370
rect 6119 4328 6143 4362
rect 6177 4328 6201 4362
rect 6119 4320 6201 4328
rect 6323 4362 6405 4370
rect 6323 4328 6347 4362
rect 6381 4328 6405 4362
rect 6323 4320 6405 4328
rect 6527 4362 6609 4370
rect 6527 4328 6551 4362
rect 6585 4328 6609 4362
rect 6527 4320 6609 4328
rect 6731 4362 6813 4370
rect 6731 4328 6755 4362
rect 6789 4328 6813 4362
rect 6731 4320 6813 4328
rect 6935 4362 7017 4370
rect 6935 4328 6959 4362
rect 6993 4328 7017 4362
rect 6935 4320 7017 4328
rect 7139 4362 7221 4370
rect 7139 4328 7163 4362
rect 7197 4328 7221 4362
rect 7139 4320 7221 4328
rect 7343 4362 7425 4370
rect 7343 4328 7367 4362
rect 7401 4328 7425 4362
rect 7343 4320 7425 4328
rect 7547 4362 7629 4370
rect 7547 4328 7571 4362
rect 7605 4328 7629 4362
rect 7547 4320 7629 4328
rect 7751 4362 7833 4370
rect 7751 4328 7775 4362
rect 7809 4328 7833 4362
rect 7751 4320 7833 4328
rect 7955 4362 8037 4370
rect 7955 4328 7979 4362
rect 8013 4328 8037 4362
rect 7955 4320 8037 4328
rect 8159 4362 8241 4370
rect 8159 4328 8183 4362
rect 8217 4328 8241 4362
rect 8159 4320 8241 4328
rect 8363 4362 8445 4370
rect 8363 4328 8387 4362
rect 8421 4328 8445 4362
rect 8363 4320 8445 4328
rect 8567 4362 8649 4370
rect 8567 4328 8591 4362
rect 8625 4328 8649 4362
rect 8567 4320 8649 4328
rect 8771 4362 8853 4370
rect 8771 4328 8795 4362
rect 8829 4328 8853 4362
rect 8771 4320 8853 4328
rect 8975 4362 9057 4370
rect 8975 4328 8999 4362
rect 9033 4328 9057 4362
rect 8975 4320 9057 4328
rect 9179 4362 9261 4370
rect 9179 4328 9203 4362
rect 9237 4328 9261 4362
rect 9179 4320 9261 4328
rect 9383 4362 9465 4370
rect 9383 4328 9407 4362
rect 9441 4328 9465 4362
rect 9383 4320 9465 4328
rect 9587 4362 9669 4370
rect 9587 4328 9611 4362
rect 9645 4328 9669 4362
rect 9587 4320 9669 4328
rect 9791 4362 9873 4370
rect 9791 4328 9815 4362
rect 9849 4328 9873 4362
rect 9791 4320 9873 4328
rect 9995 4362 10077 4370
rect 9995 4328 10019 4362
rect 10053 4328 10077 4362
rect 9995 4320 10077 4328
rect 10199 4362 10281 4370
rect 10199 4328 10223 4362
rect 10257 4328 10281 4362
rect 10199 4320 10281 4328
rect 10403 4362 10485 4370
rect 10403 4328 10427 4362
rect 10461 4328 10485 4362
rect 10403 4320 10485 4328
rect 10607 4362 10689 4370
rect 10607 4328 10631 4362
rect 10665 4328 10689 4362
rect 10607 4320 10689 4328
rect 10811 4362 10893 4370
rect 10811 4328 10835 4362
rect 10869 4328 10893 4362
rect 10811 4320 10893 4328
rect 11015 4362 11097 4370
rect 11015 4328 11039 4362
rect 11073 4328 11097 4362
rect 11015 4320 11097 4328
rect 11219 4362 11301 4370
rect 11219 4328 11243 4362
rect 11277 4328 11301 4362
rect 11219 4320 11301 4328
rect 11423 4362 11505 4370
rect 11423 4328 11447 4362
rect 11481 4328 11505 4362
rect 11423 4320 11505 4328
rect 11627 4362 11709 4370
rect 11627 4328 11651 4362
rect 11685 4328 11709 4362
rect 11627 4320 11709 4328
rect 11831 4362 11913 4370
rect 11831 4328 11855 4362
rect 11889 4328 11913 4362
rect 11831 4320 11913 4328
rect 12035 4362 12117 4370
rect 12035 4328 12059 4362
rect 12093 4328 12117 4362
rect 12035 4320 12117 4328
rect 12239 4362 12321 4370
rect 12239 4328 12263 4362
rect 12297 4328 12321 4362
rect 12239 4320 12321 4328
rect 12443 4362 12525 4370
rect 12443 4328 12467 4362
rect 12501 4328 12525 4362
rect 12443 4320 12525 4328
rect 12647 4362 12729 4370
rect 12647 4328 12671 4362
rect 12705 4328 12729 4362
rect 12647 4320 12729 4328
rect 12851 4362 12933 4370
rect 12851 4328 12875 4362
rect 12909 4328 12933 4362
rect 12851 4320 12933 4328
rect 13069 4362 13151 4370
rect 13069 4328 13093 4362
rect 13127 4328 13151 4362
rect 13069 4320 13151 4328
rect 203 2626 285 2634
rect 203 2592 227 2626
rect 261 2592 285 2626
rect 203 2584 285 2592
rect 407 2626 489 2634
rect 407 2592 431 2626
rect 465 2592 489 2626
rect 407 2584 489 2592
rect 611 2626 693 2634
rect 611 2592 635 2626
rect 669 2592 693 2626
rect 611 2584 693 2592
rect 815 2626 897 2634
rect 815 2592 839 2626
rect 873 2592 897 2626
rect 815 2584 897 2592
rect 1019 2626 1101 2634
rect 1019 2592 1043 2626
rect 1077 2592 1101 2626
rect 1019 2584 1101 2592
rect 1223 2626 1305 2634
rect 1223 2592 1247 2626
rect 1281 2592 1305 2626
rect 1223 2584 1305 2592
rect 1427 2626 1509 2634
rect 1427 2592 1451 2626
rect 1485 2592 1509 2626
rect 1427 2584 1509 2592
rect 1631 2626 1713 2634
rect 1631 2592 1655 2626
rect 1689 2592 1713 2626
rect 1631 2584 1713 2592
rect 1835 2626 1917 2634
rect 1835 2592 1859 2626
rect 1893 2592 1917 2626
rect 1835 2584 1917 2592
rect 2039 2626 2121 2634
rect 2039 2592 2063 2626
rect 2097 2592 2121 2626
rect 2039 2584 2121 2592
rect 2243 2626 2325 2634
rect 2243 2592 2267 2626
rect 2301 2592 2325 2626
rect 2243 2584 2325 2592
rect 2447 2626 2529 2634
rect 2447 2592 2471 2626
rect 2505 2592 2529 2626
rect 2447 2584 2529 2592
rect 2651 2626 2733 2634
rect 2651 2592 2675 2626
rect 2709 2592 2733 2626
rect 2651 2584 2733 2592
rect 2855 2626 2937 2634
rect 2855 2592 2879 2626
rect 2913 2592 2937 2626
rect 2855 2584 2937 2592
rect 3059 2626 3141 2634
rect 3059 2592 3083 2626
rect 3117 2592 3141 2626
rect 3059 2584 3141 2592
rect 3263 2626 3345 2634
rect 3263 2592 3287 2626
rect 3321 2592 3345 2626
rect 3263 2584 3345 2592
rect 3467 2626 3549 2634
rect 3467 2592 3491 2626
rect 3525 2592 3549 2626
rect 3467 2584 3549 2592
rect 3671 2626 3753 2634
rect 3671 2592 3695 2626
rect 3729 2592 3753 2626
rect 3671 2584 3753 2592
rect 3875 2626 3957 2634
rect 3875 2592 3899 2626
rect 3933 2592 3957 2626
rect 3875 2584 3957 2592
rect 4079 2626 4161 2634
rect 4079 2592 4103 2626
rect 4137 2592 4161 2626
rect 4079 2584 4161 2592
rect 4283 2626 4365 2634
rect 4283 2592 4307 2626
rect 4341 2592 4365 2626
rect 4283 2584 4365 2592
rect 4487 2626 4569 2634
rect 4487 2592 4511 2626
rect 4545 2592 4569 2626
rect 4487 2584 4569 2592
rect 4691 2626 4773 2634
rect 4691 2592 4715 2626
rect 4749 2592 4773 2626
rect 4691 2584 4773 2592
rect 4895 2626 4977 2634
rect 4895 2592 4919 2626
rect 4953 2592 4977 2626
rect 4895 2584 4977 2592
rect 5099 2626 5181 2634
rect 5099 2592 5123 2626
rect 5157 2592 5181 2626
rect 5099 2584 5181 2592
rect 5303 2626 5385 2634
rect 5303 2592 5327 2626
rect 5361 2592 5385 2626
rect 5303 2584 5385 2592
rect 5507 2626 5589 2634
rect 5507 2592 5531 2626
rect 5565 2592 5589 2626
rect 5507 2584 5589 2592
rect 5711 2626 5793 2634
rect 5711 2592 5735 2626
rect 5769 2592 5793 2626
rect 5711 2584 5793 2592
rect 5915 2626 5997 2634
rect 5915 2592 5939 2626
rect 5973 2592 5997 2626
rect 5915 2584 5997 2592
rect 6119 2626 6201 2634
rect 6119 2592 6143 2626
rect 6177 2592 6201 2626
rect 6119 2584 6201 2592
rect 6323 2626 6405 2634
rect 6323 2592 6347 2626
rect 6381 2592 6405 2626
rect 6323 2584 6405 2592
rect 6527 2626 6609 2634
rect 6527 2592 6551 2626
rect 6585 2592 6609 2626
rect 6527 2584 6609 2592
rect 6731 2626 6813 2634
rect 6731 2592 6755 2626
rect 6789 2592 6813 2626
rect 6731 2584 6813 2592
rect 6935 2626 7017 2634
rect 6935 2592 6959 2626
rect 6993 2592 7017 2626
rect 6935 2584 7017 2592
rect 7139 2626 7221 2634
rect 7139 2592 7163 2626
rect 7197 2592 7221 2626
rect 7139 2584 7221 2592
rect 7343 2626 7425 2634
rect 7343 2592 7367 2626
rect 7401 2592 7425 2626
rect 7343 2584 7425 2592
rect 7547 2626 7629 2634
rect 7547 2592 7571 2626
rect 7605 2592 7629 2626
rect 7547 2584 7629 2592
rect 7751 2626 7833 2634
rect 7751 2592 7775 2626
rect 7809 2592 7833 2626
rect 7751 2584 7833 2592
rect 7955 2626 8037 2634
rect 7955 2592 7979 2626
rect 8013 2592 8037 2626
rect 7955 2584 8037 2592
rect 8159 2626 8241 2634
rect 8159 2592 8183 2626
rect 8217 2592 8241 2626
rect 8159 2584 8241 2592
rect 8363 2626 8445 2634
rect 8363 2592 8387 2626
rect 8421 2592 8445 2626
rect 8363 2584 8445 2592
rect 8567 2626 8649 2634
rect 8567 2592 8591 2626
rect 8625 2592 8649 2626
rect 8567 2584 8649 2592
rect 8771 2626 8853 2634
rect 8771 2592 8795 2626
rect 8829 2592 8853 2626
rect 8771 2584 8853 2592
rect 8975 2626 9057 2634
rect 8975 2592 8999 2626
rect 9033 2592 9057 2626
rect 8975 2584 9057 2592
rect 9179 2626 9261 2634
rect 9179 2592 9203 2626
rect 9237 2592 9261 2626
rect 9179 2584 9261 2592
rect 9383 2626 9465 2634
rect 9383 2592 9407 2626
rect 9441 2592 9465 2626
rect 9383 2584 9465 2592
rect 9587 2626 9669 2634
rect 9587 2592 9611 2626
rect 9645 2592 9669 2626
rect 9587 2584 9669 2592
rect 9791 2626 9873 2634
rect 9791 2592 9815 2626
rect 9849 2592 9873 2626
rect 9791 2584 9873 2592
rect 9995 2626 10077 2634
rect 9995 2592 10019 2626
rect 10053 2592 10077 2626
rect 9995 2584 10077 2592
rect 10199 2626 10281 2634
rect 10199 2592 10223 2626
rect 10257 2592 10281 2626
rect 10199 2584 10281 2592
rect 10403 2626 10485 2634
rect 10403 2592 10427 2626
rect 10461 2592 10485 2626
rect 10403 2584 10485 2592
rect 10607 2626 10689 2634
rect 10607 2592 10631 2626
rect 10665 2592 10689 2626
rect 10607 2584 10689 2592
rect 10811 2626 10893 2634
rect 10811 2592 10835 2626
rect 10869 2592 10893 2626
rect 10811 2584 10893 2592
rect 11015 2626 11097 2634
rect 11015 2592 11039 2626
rect 11073 2592 11097 2626
rect 11015 2584 11097 2592
rect 11219 2626 11301 2634
rect 11219 2592 11243 2626
rect 11277 2592 11301 2626
rect 11219 2584 11301 2592
rect 11423 2626 11505 2634
rect 11423 2592 11447 2626
rect 11481 2592 11505 2626
rect 11423 2584 11505 2592
rect 11627 2626 11709 2634
rect 11627 2592 11651 2626
rect 11685 2592 11709 2626
rect 11627 2584 11709 2592
rect 11831 2626 11913 2634
rect 11831 2592 11855 2626
rect 11889 2592 11913 2626
rect 11831 2584 11913 2592
rect 12035 2626 12117 2634
rect 12035 2592 12059 2626
rect 12093 2592 12117 2626
rect 12035 2584 12117 2592
rect 12239 2626 12321 2634
rect 12239 2592 12263 2626
rect 12297 2592 12321 2626
rect 12239 2584 12321 2592
rect 12443 2626 12525 2634
rect 12443 2592 12467 2626
rect 12501 2592 12525 2626
rect 12443 2584 12525 2592
rect 12647 2626 12729 2634
rect 12647 2592 12671 2626
rect 12705 2592 12729 2626
rect 12647 2584 12729 2592
rect 12851 2626 12933 2634
rect 12851 2592 12875 2626
rect 12909 2592 12933 2626
rect 12851 2584 12933 2592
rect 13069 2626 13151 2634
rect 13069 2592 13093 2626
rect 13127 2592 13151 2626
rect 13069 2584 13151 2592
rect 203 890 285 898
rect 203 856 227 890
rect 261 856 285 890
rect 203 848 285 856
rect 407 890 489 898
rect 407 856 431 890
rect 465 856 489 890
rect 407 848 489 856
rect 611 890 693 898
rect 611 856 635 890
rect 669 856 693 890
rect 611 848 693 856
rect 815 890 897 898
rect 815 856 839 890
rect 873 856 897 890
rect 815 848 897 856
rect 1019 890 1101 898
rect 1019 856 1043 890
rect 1077 856 1101 890
rect 1019 848 1101 856
rect 1223 890 1305 898
rect 1223 856 1247 890
rect 1281 856 1305 890
rect 1223 848 1305 856
rect 1427 890 1509 898
rect 1427 856 1451 890
rect 1485 856 1509 890
rect 1427 848 1509 856
rect 1631 890 1713 898
rect 1631 856 1655 890
rect 1689 856 1713 890
rect 1631 848 1713 856
rect 1835 890 1917 898
rect 1835 856 1859 890
rect 1893 856 1917 890
rect 1835 848 1917 856
rect 2039 890 2121 898
rect 2039 856 2063 890
rect 2097 856 2121 890
rect 2039 848 2121 856
rect 2243 890 2325 898
rect 2243 856 2267 890
rect 2301 856 2325 890
rect 2243 848 2325 856
rect 2447 890 2529 898
rect 2447 856 2471 890
rect 2505 856 2529 890
rect 2447 848 2529 856
rect 2651 890 2733 898
rect 2651 856 2675 890
rect 2709 856 2733 890
rect 2651 848 2733 856
rect 2855 890 2937 898
rect 2855 856 2879 890
rect 2913 856 2937 890
rect 2855 848 2937 856
rect 3059 890 3141 898
rect 3059 856 3083 890
rect 3117 856 3141 890
rect 3059 848 3141 856
rect 3263 890 3345 898
rect 3263 856 3287 890
rect 3321 856 3345 890
rect 3263 848 3345 856
rect 3467 890 3549 898
rect 3467 856 3491 890
rect 3525 856 3549 890
rect 3467 848 3549 856
rect 3671 890 3753 898
rect 3671 856 3695 890
rect 3729 856 3753 890
rect 3671 848 3753 856
rect 3875 890 3957 898
rect 3875 856 3899 890
rect 3933 856 3957 890
rect 3875 848 3957 856
rect 4079 890 4161 898
rect 4079 856 4103 890
rect 4137 856 4161 890
rect 4079 848 4161 856
rect 4283 890 4365 898
rect 4283 856 4307 890
rect 4341 856 4365 890
rect 4283 848 4365 856
rect 4487 890 4569 898
rect 4487 856 4511 890
rect 4545 856 4569 890
rect 4487 848 4569 856
rect 4691 890 4773 898
rect 4691 856 4715 890
rect 4749 856 4773 890
rect 4691 848 4773 856
rect 4895 890 4977 898
rect 4895 856 4919 890
rect 4953 856 4977 890
rect 4895 848 4977 856
rect 5099 890 5181 898
rect 5099 856 5123 890
rect 5157 856 5181 890
rect 5099 848 5181 856
rect 5303 890 5385 898
rect 5303 856 5327 890
rect 5361 856 5385 890
rect 5303 848 5385 856
rect 5507 890 5589 898
rect 5507 856 5531 890
rect 5565 856 5589 890
rect 5507 848 5589 856
rect 5711 890 5793 898
rect 5711 856 5735 890
rect 5769 856 5793 890
rect 5711 848 5793 856
rect 5915 890 5997 898
rect 5915 856 5939 890
rect 5973 856 5997 890
rect 5915 848 5997 856
rect 6119 890 6201 898
rect 6119 856 6143 890
rect 6177 856 6201 890
rect 6119 848 6201 856
rect 6323 890 6405 898
rect 6323 856 6347 890
rect 6381 856 6405 890
rect 6323 848 6405 856
rect 6527 890 6609 898
rect 6527 856 6551 890
rect 6585 856 6609 890
rect 6527 848 6609 856
rect 6731 890 6813 898
rect 6731 856 6755 890
rect 6789 856 6813 890
rect 6731 848 6813 856
rect 6935 890 7017 898
rect 6935 856 6959 890
rect 6993 856 7017 890
rect 6935 848 7017 856
rect 7139 890 7221 898
rect 7139 856 7163 890
rect 7197 856 7221 890
rect 7139 848 7221 856
rect 7343 890 7425 898
rect 7343 856 7367 890
rect 7401 856 7425 890
rect 7343 848 7425 856
rect 7547 890 7629 898
rect 7547 856 7571 890
rect 7605 856 7629 890
rect 7547 848 7629 856
rect 7751 890 7833 898
rect 7751 856 7775 890
rect 7809 856 7833 890
rect 7751 848 7833 856
rect 7955 890 8037 898
rect 7955 856 7979 890
rect 8013 856 8037 890
rect 7955 848 8037 856
rect 8159 890 8241 898
rect 8159 856 8183 890
rect 8217 856 8241 890
rect 8159 848 8241 856
rect 8363 890 8445 898
rect 8363 856 8387 890
rect 8421 856 8445 890
rect 8363 848 8445 856
rect 8567 890 8649 898
rect 8567 856 8591 890
rect 8625 856 8649 890
rect 8567 848 8649 856
rect 8771 890 8853 898
rect 8771 856 8795 890
rect 8829 856 8853 890
rect 8771 848 8853 856
rect 8975 890 9057 898
rect 8975 856 8999 890
rect 9033 856 9057 890
rect 8975 848 9057 856
rect 9179 890 9261 898
rect 9179 856 9203 890
rect 9237 856 9261 890
rect 9179 848 9261 856
rect 9383 890 9465 898
rect 9383 856 9407 890
rect 9441 856 9465 890
rect 9383 848 9465 856
rect 9587 890 9669 898
rect 9587 856 9611 890
rect 9645 856 9669 890
rect 9587 848 9669 856
rect 9791 890 9873 898
rect 9791 856 9815 890
rect 9849 856 9873 890
rect 9791 848 9873 856
rect 9995 890 10077 898
rect 9995 856 10019 890
rect 10053 856 10077 890
rect 9995 848 10077 856
rect 10199 890 10281 898
rect 10199 856 10223 890
rect 10257 856 10281 890
rect 10199 848 10281 856
rect 10403 890 10485 898
rect 10403 856 10427 890
rect 10461 856 10485 890
rect 10403 848 10485 856
rect 10607 890 10689 898
rect 10607 856 10631 890
rect 10665 856 10689 890
rect 10607 848 10689 856
rect 10811 890 10893 898
rect 10811 856 10835 890
rect 10869 856 10893 890
rect 10811 848 10893 856
rect 11015 890 11097 898
rect 11015 856 11039 890
rect 11073 856 11097 890
rect 11015 848 11097 856
rect 11219 890 11301 898
rect 11219 856 11243 890
rect 11277 856 11301 890
rect 11219 848 11301 856
rect 11423 890 11505 898
rect 11423 856 11447 890
rect 11481 856 11505 890
rect 11423 848 11505 856
rect 11627 890 11709 898
rect 11627 856 11651 890
rect 11685 856 11709 890
rect 11627 848 11709 856
rect 11831 890 11913 898
rect 11831 856 11855 890
rect 11889 856 11913 890
rect 11831 848 11913 856
rect 12035 890 12117 898
rect 12035 856 12059 890
rect 12093 856 12117 890
rect 12035 848 12117 856
rect 12239 890 12321 898
rect 12239 856 12263 890
rect 12297 856 12321 890
rect 12239 848 12321 856
rect 12443 890 12525 898
rect 12443 856 12467 890
rect 12501 856 12525 890
rect 12443 848 12525 856
rect 12647 890 12729 898
rect 12647 856 12671 890
rect 12705 856 12729 890
rect 12647 848 12729 856
rect 12851 890 12933 898
rect 12851 856 12875 890
rect 12909 856 12933 890
rect 12851 848 12933 856
rect 13069 890 13151 898
rect 13069 856 13093 890
rect 13127 856 13151 890
rect 13069 848 13151 856
<< psubdiffcont >>
rect 227 6064 261 6098
rect 431 6064 465 6098
rect 635 6064 669 6098
rect 839 6064 873 6098
rect 1043 6064 1077 6098
rect 1247 6064 1281 6098
rect 1451 6064 1485 6098
rect 1655 6064 1689 6098
rect 1859 6064 1893 6098
rect 2063 6064 2097 6098
rect 2267 6064 2301 6098
rect 2471 6064 2505 6098
rect 2675 6064 2709 6098
rect 2879 6064 2913 6098
rect 3083 6064 3117 6098
rect 3287 6064 3321 6098
rect 3491 6064 3525 6098
rect 3695 6064 3729 6098
rect 3899 6064 3933 6098
rect 4103 6064 4137 6098
rect 4307 6064 4341 6098
rect 4511 6064 4545 6098
rect 4715 6064 4749 6098
rect 4919 6064 4953 6098
rect 5123 6064 5157 6098
rect 5327 6064 5361 6098
rect 5531 6064 5565 6098
rect 5735 6064 5769 6098
rect 5939 6064 5973 6098
rect 6143 6064 6177 6098
rect 6347 6064 6381 6098
rect 6551 6064 6585 6098
rect 6755 6064 6789 6098
rect 6959 6064 6993 6098
rect 7163 6064 7197 6098
rect 7367 6064 7401 6098
rect 7571 6064 7605 6098
rect 7775 6064 7809 6098
rect 7979 6064 8013 6098
rect 8183 6064 8217 6098
rect 8387 6064 8421 6098
rect 8591 6064 8625 6098
rect 8795 6064 8829 6098
rect 8999 6064 9033 6098
rect 9203 6064 9237 6098
rect 9407 6064 9441 6098
rect 9611 6064 9645 6098
rect 9815 6064 9849 6098
rect 10019 6064 10053 6098
rect 10223 6064 10257 6098
rect 10427 6064 10461 6098
rect 10631 6064 10665 6098
rect 10835 6064 10869 6098
rect 11039 6064 11073 6098
rect 11243 6064 11277 6098
rect 11447 6064 11481 6098
rect 11651 6064 11685 6098
rect 11855 6064 11889 6098
rect 12059 6064 12093 6098
rect 12263 6064 12297 6098
rect 12467 6064 12501 6098
rect 12671 6064 12705 6098
rect 12875 6064 12909 6098
rect 13093 6064 13127 6098
rect 227 4328 261 4362
rect 431 4328 465 4362
rect 635 4328 669 4362
rect 839 4328 873 4362
rect 1043 4328 1077 4362
rect 1247 4328 1281 4362
rect 1451 4328 1485 4362
rect 1655 4328 1689 4362
rect 1859 4328 1893 4362
rect 2063 4328 2097 4362
rect 2267 4328 2301 4362
rect 2471 4328 2505 4362
rect 2675 4328 2709 4362
rect 2879 4328 2913 4362
rect 3083 4328 3117 4362
rect 3287 4328 3321 4362
rect 3491 4328 3525 4362
rect 3695 4328 3729 4362
rect 3899 4328 3933 4362
rect 4103 4328 4137 4362
rect 4307 4328 4341 4362
rect 4511 4328 4545 4362
rect 4715 4328 4749 4362
rect 4919 4328 4953 4362
rect 5123 4328 5157 4362
rect 5327 4328 5361 4362
rect 5531 4328 5565 4362
rect 5735 4328 5769 4362
rect 5939 4328 5973 4362
rect 6143 4328 6177 4362
rect 6347 4328 6381 4362
rect 6551 4328 6585 4362
rect 6755 4328 6789 4362
rect 6959 4328 6993 4362
rect 7163 4328 7197 4362
rect 7367 4328 7401 4362
rect 7571 4328 7605 4362
rect 7775 4328 7809 4362
rect 7979 4328 8013 4362
rect 8183 4328 8217 4362
rect 8387 4328 8421 4362
rect 8591 4328 8625 4362
rect 8795 4328 8829 4362
rect 8999 4328 9033 4362
rect 9203 4328 9237 4362
rect 9407 4328 9441 4362
rect 9611 4328 9645 4362
rect 9815 4328 9849 4362
rect 10019 4328 10053 4362
rect 10223 4328 10257 4362
rect 10427 4328 10461 4362
rect 10631 4328 10665 4362
rect 10835 4328 10869 4362
rect 11039 4328 11073 4362
rect 11243 4328 11277 4362
rect 11447 4328 11481 4362
rect 11651 4328 11685 4362
rect 11855 4328 11889 4362
rect 12059 4328 12093 4362
rect 12263 4328 12297 4362
rect 12467 4328 12501 4362
rect 12671 4328 12705 4362
rect 12875 4328 12909 4362
rect 13093 4328 13127 4362
rect 227 2592 261 2626
rect 431 2592 465 2626
rect 635 2592 669 2626
rect 839 2592 873 2626
rect 1043 2592 1077 2626
rect 1247 2592 1281 2626
rect 1451 2592 1485 2626
rect 1655 2592 1689 2626
rect 1859 2592 1893 2626
rect 2063 2592 2097 2626
rect 2267 2592 2301 2626
rect 2471 2592 2505 2626
rect 2675 2592 2709 2626
rect 2879 2592 2913 2626
rect 3083 2592 3117 2626
rect 3287 2592 3321 2626
rect 3491 2592 3525 2626
rect 3695 2592 3729 2626
rect 3899 2592 3933 2626
rect 4103 2592 4137 2626
rect 4307 2592 4341 2626
rect 4511 2592 4545 2626
rect 4715 2592 4749 2626
rect 4919 2592 4953 2626
rect 5123 2592 5157 2626
rect 5327 2592 5361 2626
rect 5531 2592 5565 2626
rect 5735 2592 5769 2626
rect 5939 2592 5973 2626
rect 6143 2592 6177 2626
rect 6347 2592 6381 2626
rect 6551 2592 6585 2626
rect 6755 2592 6789 2626
rect 6959 2592 6993 2626
rect 7163 2592 7197 2626
rect 7367 2592 7401 2626
rect 7571 2592 7605 2626
rect 7775 2592 7809 2626
rect 7979 2592 8013 2626
rect 8183 2592 8217 2626
rect 8387 2592 8421 2626
rect 8591 2592 8625 2626
rect 8795 2592 8829 2626
rect 8999 2592 9033 2626
rect 9203 2592 9237 2626
rect 9407 2592 9441 2626
rect 9611 2592 9645 2626
rect 9815 2592 9849 2626
rect 10019 2592 10053 2626
rect 10223 2592 10257 2626
rect 10427 2592 10461 2626
rect 10631 2592 10665 2626
rect 10835 2592 10869 2626
rect 11039 2592 11073 2626
rect 11243 2592 11277 2626
rect 11447 2592 11481 2626
rect 11651 2592 11685 2626
rect 11855 2592 11889 2626
rect 12059 2592 12093 2626
rect 12263 2592 12297 2626
rect 12467 2592 12501 2626
rect 12671 2592 12705 2626
rect 12875 2592 12909 2626
rect 13093 2592 13127 2626
rect 227 856 261 890
rect 431 856 465 890
rect 635 856 669 890
rect 839 856 873 890
rect 1043 856 1077 890
rect 1247 856 1281 890
rect 1451 856 1485 890
rect 1655 856 1689 890
rect 1859 856 1893 890
rect 2063 856 2097 890
rect 2267 856 2301 890
rect 2471 856 2505 890
rect 2675 856 2709 890
rect 2879 856 2913 890
rect 3083 856 3117 890
rect 3287 856 3321 890
rect 3491 856 3525 890
rect 3695 856 3729 890
rect 3899 856 3933 890
rect 4103 856 4137 890
rect 4307 856 4341 890
rect 4511 856 4545 890
rect 4715 856 4749 890
rect 4919 856 4953 890
rect 5123 856 5157 890
rect 5327 856 5361 890
rect 5531 856 5565 890
rect 5735 856 5769 890
rect 5939 856 5973 890
rect 6143 856 6177 890
rect 6347 856 6381 890
rect 6551 856 6585 890
rect 6755 856 6789 890
rect 6959 856 6993 890
rect 7163 856 7197 890
rect 7367 856 7401 890
rect 7571 856 7605 890
rect 7775 856 7809 890
rect 7979 856 8013 890
rect 8183 856 8217 890
rect 8387 856 8421 890
rect 8591 856 8625 890
rect 8795 856 8829 890
rect 8999 856 9033 890
rect 9203 856 9237 890
rect 9407 856 9441 890
rect 9611 856 9645 890
rect 9815 856 9849 890
rect 10019 856 10053 890
rect 10223 856 10257 890
rect 10427 856 10461 890
rect 10631 856 10665 890
rect 10835 856 10869 890
rect 11039 856 11073 890
rect 11243 856 11277 890
rect 11447 856 11481 890
rect 11651 856 11685 890
rect 11855 856 11889 890
rect 12059 856 12093 890
rect 12263 856 12297 890
rect 12467 856 12501 890
rect 12671 856 12705 890
rect 12875 856 12909 890
rect 13093 856 13127 890
<< poly >>
rect 0 7884 66 7900
rect 0 7850 16 7884
rect 50 7882 66 7884
rect 1632 7884 1698 7900
rect 1632 7882 1648 7884
rect 50 7852 1648 7882
rect 50 7850 66 7852
rect 0 7834 66 7850
rect 1632 7850 1648 7852
rect 1682 7882 1698 7884
rect 3264 7884 3330 7900
rect 3264 7882 3280 7884
rect 1682 7852 3280 7882
rect 1682 7850 1698 7852
rect 1632 7834 1698 7850
rect 3264 7850 3280 7852
rect 3314 7882 3330 7884
rect 4896 7884 4962 7900
rect 4896 7882 4912 7884
rect 3314 7852 4912 7882
rect 3314 7850 3330 7852
rect 3264 7834 3330 7850
rect 4896 7850 4912 7852
rect 4946 7882 4962 7884
rect 6528 7884 6594 7900
rect 6528 7882 6544 7884
rect 4946 7852 6544 7882
rect 4946 7850 4962 7852
rect 4896 7834 4962 7850
rect 6528 7850 6544 7852
rect 6578 7882 6594 7884
rect 8160 7884 8226 7900
rect 8160 7882 8176 7884
rect 6578 7852 8176 7882
rect 6578 7850 6594 7852
rect 6528 7834 6594 7850
rect 8160 7850 8176 7852
rect 8210 7882 8226 7884
rect 9792 7884 9858 7900
rect 9792 7882 9808 7884
rect 8210 7852 9808 7882
rect 8210 7850 8226 7852
rect 8160 7834 8226 7850
rect 9792 7850 9808 7852
rect 9842 7882 9858 7884
rect 11424 7884 11490 7900
rect 11424 7882 11440 7884
rect 9842 7852 11440 7882
rect 9842 7850 9858 7852
rect 9792 7834 9858 7850
rect 11424 7850 11440 7852
rect 11474 7882 11490 7884
rect 13056 7884 13122 7900
rect 13056 7882 13072 7884
rect 11474 7852 13072 7882
rect 11474 7850 11490 7852
rect 11424 7834 11490 7850
rect 13056 7850 13072 7852
rect 13106 7850 13122 7884
rect 13056 7834 13122 7850
rect 0 7680 66 7696
rect 0 7646 16 7680
rect 50 7678 66 7680
rect 1632 7680 1698 7696
rect 1632 7678 1648 7680
rect 50 7648 1648 7678
rect 50 7646 66 7648
rect 0 7630 66 7646
rect 1632 7646 1648 7648
rect 1682 7678 1698 7680
rect 3264 7680 3330 7696
rect 3264 7678 3280 7680
rect 1682 7648 3280 7678
rect 1682 7646 1698 7648
rect 1632 7630 1698 7646
rect 3264 7646 3280 7648
rect 3314 7678 3330 7680
rect 4896 7680 4962 7696
rect 4896 7678 4912 7680
rect 3314 7648 4912 7678
rect 3314 7646 3330 7648
rect 3264 7630 3330 7646
rect 4896 7646 4912 7648
rect 4946 7678 4962 7680
rect 6528 7680 6594 7696
rect 6528 7678 6544 7680
rect 4946 7648 6544 7678
rect 4946 7646 4962 7648
rect 4896 7630 4962 7646
rect 6528 7646 6544 7648
rect 6578 7678 6594 7680
rect 8160 7680 8226 7696
rect 8160 7678 8176 7680
rect 6578 7648 8176 7678
rect 6578 7646 6594 7648
rect 6528 7630 6594 7646
rect 8160 7646 8176 7648
rect 8210 7678 8226 7680
rect 9792 7680 9858 7696
rect 9792 7678 9808 7680
rect 8210 7648 9808 7678
rect 8210 7646 8226 7648
rect 8160 7630 8226 7646
rect 9792 7646 9808 7648
rect 9842 7678 9858 7680
rect 11424 7680 11490 7696
rect 11424 7678 11440 7680
rect 9842 7648 11440 7678
rect 9842 7646 9858 7648
rect 9792 7630 9858 7646
rect 11424 7646 11440 7648
rect 11474 7678 11490 7680
rect 13056 7680 13122 7696
rect 13056 7678 13072 7680
rect 11474 7648 13072 7678
rect 11474 7646 11490 7648
rect 11424 7630 11490 7646
rect 13056 7646 13072 7648
rect 13106 7646 13122 7680
rect 13056 7630 13122 7646
rect 0 7476 66 7492
rect 0 7442 16 7476
rect 50 7474 66 7476
rect 1632 7476 1698 7492
rect 1632 7474 1648 7476
rect 50 7444 1648 7474
rect 50 7442 66 7444
rect 0 7426 66 7442
rect 1632 7442 1648 7444
rect 1682 7474 1698 7476
rect 3264 7476 3330 7492
rect 3264 7474 3280 7476
rect 1682 7444 3280 7474
rect 1682 7442 1698 7444
rect 1632 7426 1698 7442
rect 3264 7442 3280 7444
rect 3314 7474 3330 7476
rect 4896 7476 4962 7492
rect 4896 7474 4912 7476
rect 3314 7444 4912 7474
rect 3314 7442 3330 7444
rect 3264 7426 3330 7442
rect 4896 7442 4912 7444
rect 4946 7474 4962 7476
rect 6528 7476 6594 7492
rect 6528 7474 6544 7476
rect 4946 7444 6544 7474
rect 4946 7442 4962 7444
rect 4896 7426 4962 7442
rect 6528 7442 6544 7444
rect 6578 7474 6594 7476
rect 8160 7476 8226 7492
rect 8160 7474 8176 7476
rect 6578 7444 8176 7474
rect 6578 7442 6594 7444
rect 6528 7426 6594 7442
rect 8160 7442 8176 7444
rect 8210 7474 8226 7476
rect 9792 7476 9858 7492
rect 9792 7474 9808 7476
rect 8210 7444 9808 7474
rect 8210 7442 8226 7444
rect 8160 7426 8226 7442
rect 9792 7442 9808 7444
rect 9842 7474 9858 7476
rect 11424 7476 11490 7492
rect 11424 7474 11440 7476
rect 9842 7444 11440 7474
rect 9842 7442 9858 7444
rect 9792 7426 9858 7442
rect 11424 7442 11440 7444
rect 11474 7474 11490 7476
rect 13056 7476 13122 7492
rect 13056 7474 13072 7476
rect 11474 7444 13072 7474
rect 11474 7442 11490 7444
rect 11424 7426 11490 7442
rect 13056 7442 13072 7444
rect 13106 7442 13122 7476
rect 13056 7426 13122 7442
rect 0 7272 66 7288
rect 0 7238 16 7272
rect 50 7270 66 7272
rect 1632 7272 1698 7288
rect 1632 7270 1648 7272
rect 50 7240 1648 7270
rect 50 7238 66 7240
rect 0 7222 66 7238
rect 1632 7238 1648 7240
rect 1682 7270 1698 7272
rect 3264 7272 3330 7288
rect 3264 7270 3280 7272
rect 1682 7240 3280 7270
rect 1682 7238 1698 7240
rect 1632 7222 1698 7238
rect 3264 7238 3280 7240
rect 3314 7270 3330 7272
rect 4896 7272 4962 7288
rect 4896 7270 4912 7272
rect 3314 7240 4912 7270
rect 3314 7238 3330 7240
rect 3264 7222 3330 7238
rect 4896 7238 4912 7240
rect 4946 7270 4962 7272
rect 6528 7272 6594 7288
rect 6528 7270 6544 7272
rect 4946 7240 6544 7270
rect 4946 7238 4962 7240
rect 4896 7222 4962 7238
rect 6528 7238 6544 7240
rect 6578 7270 6594 7272
rect 8160 7272 8226 7288
rect 8160 7270 8176 7272
rect 6578 7240 8176 7270
rect 6578 7238 6594 7240
rect 6528 7222 6594 7238
rect 8160 7238 8176 7240
rect 8210 7270 8226 7272
rect 9792 7272 9858 7288
rect 9792 7270 9808 7272
rect 8210 7240 9808 7270
rect 8210 7238 8226 7240
rect 8160 7222 8226 7238
rect 9792 7238 9808 7240
rect 9842 7270 9858 7272
rect 11424 7272 11490 7288
rect 11424 7270 11440 7272
rect 9842 7240 11440 7270
rect 9842 7238 9858 7240
rect 9792 7222 9858 7238
rect 11424 7238 11440 7240
rect 11474 7270 11490 7272
rect 13056 7272 13122 7288
rect 13056 7270 13072 7272
rect 11474 7240 13072 7270
rect 11474 7238 11490 7240
rect 11424 7222 11490 7238
rect 13056 7238 13072 7240
rect 13106 7238 13122 7272
rect 13056 7222 13122 7238
rect 0 7068 66 7084
rect 0 7034 16 7068
rect 50 7066 66 7068
rect 1632 7068 1698 7084
rect 1632 7066 1648 7068
rect 50 7036 1648 7066
rect 50 7034 66 7036
rect 0 7018 66 7034
rect 1632 7034 1648 7036
rect 1682 7066 1698 7068
rect 3264 7068 3330 7084
rect 3264 7066 3280 7068
rect 1682 7036 3280 7066
rect 1682 7034 1698 7036
rect 1632 7018 1698 7034
rect 3264 7034 3280 7036
rect 3314 7066 3330 7068
rect 4896 7068 4962 7084
rect 4896 7066 4912 7068
rect 3314 7036 4912 7066
rect 3314 7034 3330 7036
rect 3264 7018 3330 7034
rect 4896 7034 4912 7036
rect 4946 7066 4962 7068
rect 6528 7068 6594 7084
rect 6528 7066 6544 7068
rect 4946 7036 6544 7066
rect 4946 7034 4962 7036
rect 4896 7018 4962 7034
rect 6528 7034 6544 7036
rect 6578 7066 6594 7068
rect 8160 7068 8226 7084
rect 8160 7066 8176 7068
rect 6578 7036 8176 7066
rect 6578 7034 6594 7036
rect 6528 7018 6594 7034
rect 8160 7034 8176 7036
rect 8210 7066 8226 7068
rect 9792 7068 9858 7084
rect 9792 7066 9808 7068
rect 8210 7036 9808 7066
rect 8210 7034 8226 7036
rect 8160 7018 8226 7034
rect 9792 7034 9808 7036
rect 9842 7066 9858 7068
rect 11424 7068 11490 7084
rect 11424 7066 11440 7068
rect 9842 7036 11440 7066
rect 9842 7034 9858 7036
rect 9792 7018 9858 7034
rect 11424 7034 11440 7036
rect 11474 7066 11490 7068
rect 13056 7068 13122 7084
rect 13056 7066 13072 7068
rect 11474 7036 13072 7066
rect 11474 7034 11490 7036
rect 11424 7018 11490 7034
rect 13056 7034 13072 7036
rect 13106 7034 13122 7068
rect 13056 7018 13122 7034
rect 0 6864 66 6880
rect 0 6830 16 6864
rect 50 6862 66 6864
rect 1632 6864 1698 6880
rect 1632 6862 1648 6864
rect 50 6832 1648 6862
rect 50 6830 66 6832
rect 0 6814 66 6830
rect 1632 6830 1648 6832
rect 1682 6862 1698 6864
rect 3264 6864 3330 6880
rect 3264 6862 3280 6864
rect 1682 6832 3280 6862
rect 1682 6830 1698 6832
rect 1632 6814 1698 6830
rect 3264 6830 3280 6832
rect 3314 6862 3330 6864
rect 4896 6864 4962 6880
rect 4896 6862 4912 6864
rect 3314 6832 4912 6862
rect 3314 6830 3330 6832
rect 3264 6814 3330 6830
rect 4896 6830 4912 6832
rect 4946 6862 4962 6864
rect 6528 6864 6594 6880
rect 6528 6862 6544 6864
rect 4946 6832 6544 6862
rect 4946 6830 4962 6832
rect 4896 6814 4962 6830
rect 6528 6830 6544 6832
rect 6578 6862 6594 6864
rect 8160 6864 8226 6880
rect 8160 6862 8176 6864
rect 6578 6832 8176 6862
rect 6578 6830 6594 6832
rect 6528 6814 6594 6830
rect 8160 6830 8176 6832
rect 8210 6862 8226 6864
rect 9792 6864 9858 6880
rect 9792 6862 9808 6864
rect 8210 6832 9808 6862
rect 8210 6830 8226 6832
rect 8160 6814 8226 6830
rect 9792 6830 9808 6832
rect 9842 6862 9858 6864
rect 11424 6864 11490 6880
rect 11424 6862 11440 6864
rect 9842 6832 11440 6862
rect 9842 6830 9858 6832
rect 9792 6814 9858 6830
rect 11424 6830 11440 6832
rect 11474 6862 11490 6864
rect 13056 6864 13122 6880
rect 13056 6862 13072 6864
rect 11474 6832 13072 6862
rect 11474 6830 11490 6832
rect 11424 6814 11490 6830
rect 13056 6830 13072 6832
rect 13106 6830 13122 6864
rect 13056 6814 13122 6830
rect 0 6660 66 6676
rect 0 6626 16 6660
rect 50 6658 66 6660
rect 1632 6660 1698 6676
rect 1632 6658 1648 6660
rect 50 6628 1648 6658
rect 50 6626 66 6628
rect 0 6610 66 6626
rect 1632 6626 1648 6628
rect 1682 6658 1698 6660
rect 3264 6660 3330 6676
rect 3264 6658 3280 6660
rect 1682 6628 3280 6658
rect 1682 6626 1698 6628
rect 1632 6610 1698 6626
rect 3264 6626 3280 6628
rect 3314 6658 3330 6660
rect 4896 6660 4962 6676
rect 4896 6658 4912 6660
rect 3314 6628 4912 6658
rect 3314 6626 3330 6628
rect 3264 6610 3330 6626
rect 4896 6626 4912 6628
rect 4946 6658 4962 6660
rect 6528 6660 6594 6676
rect 6528 6658 6544 6660
rect 4946 6628 6544 6658
rect 4946 6626 4962 6628
rect 4896 6610 4962 6626
rect 6528 6626 6544 6628
rect 6578 6658 6594 6660
rect 8160 6660 8226 6676
rect 8160 6658 8176 6660
rect 6578 6628 8176 6658
rect 6578 6626 6594 6628
rect 6528 6610 6594 6626
rect 8160 6626 8176 6628
rect 8210 6658 8226 6660
rect 9792 6660 9858 6676
rect 9792 6658 9808 6660
rect 8210 6628 9808 6658
rect 8210 6626 8226 6628
rect 8160 6610 8226 6626
rect 9792 6626 9808 6628
rect 9842 6658 9858 6660
rect 11424 6660 11490 6676
rect 11424 6658 11440 6660
rect 9842 6628 11440 6658
rect 9842 6626 9858 6628
rect 9792 6610 9858 6626
rect 11424 6626 11440 6628
rect 11474 6658 11490 6660
rect 13056 6660 13122 6676
rect 13056 6658 13072 6660
rect 11474 6628 13072 6658
rect 11474 6626 11490 6628
rect 11424 6610 11490 6626
rect 13056 6626 13072 6628
rect 13106 6626 13122 6660
rect 13056 6610 13122 6626
rect 0 6456 66 6472
rect 0 6422 16 6456
rect 50 6454 66 6456
rect 1632 6456 1698 6472
rect 1632 6454 1648 6456
rect 50 6424 1648 6454
rect 50 6422 66 6424
rect 0 6406 66 6422
rect 1632 6422 1648 6424
rect 1682 6454 1698 6456
rect 3264 6456 3330 6472
rect 3264 6454 3280 6456
rect 1682 6424 3280 6454
rect 1682 6422 1698 6424
rect 1632 6406 1698 6422
rect 3264 6422 3280 6424
rect 3314 6454 3330 6456
rect 4896 6456 4962 6472
rect 4896 6454 4912 6456
rect 3314 6424 4912 6454
rect 3314 6422 3330 6424
rect 3264 6406 3330 6422
rect 4896 6422 4912 6424
rect 4946 6454 4962 6456
rect 6528 6456 6594 6472
rect 6528 6454 6544 6456
rect 4946 6424 6544 6454
rect 4946 6422 4962 6424
rect 4896 6406 4962 6422
rect 6528 6422 6544 6424
rect 6578 6454 6594 6456
rect 8160 6456 8226 6472
rect 8160 6454 8176 6456
rect 6578 6424 8176 6454
rect 6578 6422 6594 6424
rect 6528 6406 6594 6422
rect 8160 6422 8176 6424
rect 8210 6454 8226 6456
rect 9792 6456 9858 6472
rect 9792 6454 9808 6456
rect 8210 6424 9808 6454
rect 8210 6422 8226 6424
rect 8160 6406 8226 6422
rect 9792 6422 9808 6424
rect 9842 6454 9858 6456
rect 11424 6456 11490 6472
rect 11424 6454 11440 6456
rect 9842 6424 11440 6454
rect 9842 6422 9858 6424
rect 9792 6406 9858 6422
rect 11424 6422 11440 6424
rect 11474 6454 11490 6456
rect 13056 6456 13122 6472
rect 13056 6454 13072 6456
rect 11474 6424 13072 6454
rect 11474 6422 11490 6424
rect 11424 6406 11490 6422
rect 13056 6422 13072 6424
rect 13106 6422 13122 6456
rect 13056 6406 13122 6422
rect 0 6252 66 6268
rect 0 6218 16 6252
rect 50 6250 66 6252
rect 1632 6252 1698 6268
rect 1632 6250 1648 6252
rect 50 6220 1648 6250
rect 50 6218 66 6220
rect 0 6202 66 6218
rect 1632 6218 1648 6220
rect 1682 6250 1698 6252
rect 3264 6252 3330 6268
rect 3264 6250 3280 6252
rect 1682 6220 3280 6250
rect 1682 6218 1698 6220
rect 1632 6202 1698 6218
rect 3264 6218 3280 6220
rect 3314 6250 3330 6252
rect 4896 6252 4962 6268
rect 4896 6250 4912 6252
rect 3314 6220 4912 6250
rect 3314 6218 3330 6220
rect 3264 6202 3330 6218
rect 4896 6218 4912 6220
rect 4946 6250 4962 6252
rect 6528 6252 6594 6268
rect 6528 6250 6544 6252
rect 4946 6220 6544 6250
rect 4946 6218 4962 6220
rect 4896 6202 4962 6218
rect 6528 6218 6544 6220
rect 6578 6250 6594 6252
rect 8160 6252 8226 6268
rect 8160 6250 8176 6252
rect 6578 6220 8176 6250
rect 6578 6218 6594 6220
rect 6528 6202 6594 6218
rect 8160 6218 8176 6220
rect 8210 6250 8226 6252
rect 9792 6252 9858 6268
rect 9792 6250 9808 6252
rect 8210 6220 9808 6250
rect 8210 6218 8226 6220
rect 8160 6202 8226 6218
rect 9792 6218 9808 6220
rect 9842 6250 9858 6252
rect 11424 6252 11490 6268
rect 11424 6250 11440 6252
rect 9842 6220 11440 6250
rect 9842 6218 9858 6220
rect 9792 6202 9858 6218
rect 11424 6218 11440 6220
rect 11474 6250 11490 6252
rect 13056 6252 13122 6268
rect 13056 6250 13072 6252
rect 11474 6220 13072 6250
rect 11474 6218 11490 6220
rect 11424 6202 11490 6218
rect 13056 6218 13072 6220
rect 13106 6218 13122 6252
rect 13056 6202 13122 6218
rect 0 5944 66 5960
rect 0 5910 16 5944
rect 50 5942 66 5944
rect 1632 5944 1698 5960
rect 1632 5942 1648 5944
rect 50 5912 1648 5942
rect 50 5910 66 5912
rect 0 5894 66 5910
rect 1632 5910 1648 5912
rect 1682 5942 1698 5944
rect 3264 5944 3330 5960
rect 3264 5942 3280 5944
rect 1682 5912 3280 5942
rect 1682 5910 1698 5912
rect 1632 5894 1698 5910
rect 3264 5910 3280 5912
rect 3314 5942 3330 5944
rect 4896 5944 4962 5960
rect 4896 5942 4912 5944
rect 3314 5912 4912 5942
rect 3314 5910 3330 5912
rect 3264 5894 3330 5910
rect 4896 5910 4912 5912
rect 4946 5942 4962 5944
rect 6528 5944 6594 5960
rect 6528 5942 6544 5944
rect 4946 5912 6544 5942
rect 4946 5910 4962 5912
rect 4896 5894 4962 5910
rect 6528 5910 6544 5912
rect 6578 5942 6594 5944
rect 8160 5944 8226 5960
rect 8160 5942 8176 5944
rect 6578 5912 8176 5942
rect 6578 5910 6594 5912
rect 6528 5894 6594 5910
rect 8160 5910 8176 5912
rect 8210 5942 8226 5944
rect 9792 5944 9858 5960
rect 9792 5942 9808 5944
rect 8210 5912 9808 5942
rect 8210 5910 8226 5912
rect 8160 5894 8226 5910
rect 9792 5910 9808 5912
rect 9842 5942 9858 5944
rect 11424 5944 11490 5960
rect 11424 5942 11440 5944
rect 9842 5912 11440 5942
rect 9842 5910 9858 5912
rect 9792 5894 9858 5910
rect 11424 5910 11440 5912
rect 11474 5942 11490 5944
rect 13056 5944 13122 5960
rect 13056 5942 13072 5944
rect 11474 5912 13072 5942
rect 11474 5910 11490 5912
rect 11424 5894 11490 5910
rect 13056 5910 13072 5912
rect 13106 5910 13122 5944
rect 13056 5894 13122 5910
rect 0 5740 66 5756
rect 0 5706 16 5740
rect 50 5738 66 5740
rect 1632 5740 1698 5756
rect 1632 5738 1648 5740
rect 50 5708 1648 5738
rect 50 5706 66 5708
rect 0 5690 66 5706
rect 1632 5706 1648 5708
rect 1682 5738 1698 5740
rect 3264 5740 3330 5756
rect 3264 5738 3280 5740
rect 1682 5708 3280 5738
rect 1682 5706 1698 5708
rect 1632 5690 1698 5706
rect 3264 5706 3280 5708
rect 3314 5738 3330 5740
rect 4896 5740 4962 5756
rect 4896 5738 4912 5740
rect 3314 5708 4912 5738
rect 3314 5706 3330 5708
rect 3264 5690 3330 5706
rect 4896 5706 4912 5708
rect 4946 5738 4962 5740
rect 6528 5740 6594 5756
rect 6528 5738 6544 5740
rect 4946 5708 6544 5738
rect 4946 5706 4962 5708
rect 4896 5690 4962 5706
rect 6528 5706 6544 5708
rect 6578 5738 6594 5740
rect 8160 5740 8226 5756
rect 8160 5738 8176 5740
rect 6578 5708 8176 5738
rect 6578 5706 6594 5708
rect 6528 5690 6594 5706
rect 8160 5706 8176 5708
rect 8210 5738 8226 5740
rect 9792 5740 9858 5756
rect 9792 5738 9808 5740
rect 8210 5708 9808 5738
rect 8210 5706 8226 5708
rect 8160 5690 8226 5706
rect 9792 5706 9808 5708
rect 9842 5738 9858 5740
rect 11424 5740 11490 5756
rect 11424 5738 11440 5740
rect 9842 5708 11440 5738
rect 9842 5706 9858 5708
rect 9792 5690 9858 5706
rect 11424 5706 11440 5708
rect 11474 5738 11490 5740
rect 13056 5740 13122 5756
rect 13056 5738 13072 5740
rect 11474 5708 13072 5738
rect 11474 5706 11490 5708
rect 11424 5690 11490 5706
rect 13056 5706 13072 5708
rect 13106 5706 13122 5740
rect 13056 5690 13122 5706
rect 0 5536 66 5552
rect 0 5502 16 5536
rect 50 5534 66 5536
rect 1632 5536 1698 5552
rect 1632 5534 1648 5536
rect 50 5504 1648 5534
rect 50 5502 66 5504
rect 0 5486 66 5502
rect 1632 5502 1648 5504
rect 1682 5534 1698 5536
rect 3264 5536 3330 5552
rect 3264 5534 3280 5536
rect 1682 5504 3280 5534
rect 1682 5502 1698 5504
rect 1632 5486 1698 5502
rect 3264 5502 3280 5504
rect 3314 5534 3330 5536
rect 4896 5536 4962 5552
rect 4896 5534 4912 5536
rect 3314 5504 4912 5534
rect 3314 5502 3330 5504
rect 3264 5486 3330 5502
rect 4896 5502 4912 5504
rect 4946 5534 4962 5536
rect 6528 5536 6594 5552
rect 6528 5534 6544 5536
rect 4946 5504 6544 5534
rect 4946 5502 4962 5504
rect 4896 5486 4962 5502
rect 6528 5502 6544 5504
rect 6578 5534 6594 5536
rect 8160 5536 8226 5552
rect 8160 5534 8176 5536
rect 6578 5504 8176 5534
rect 6578 5502 6594 5504
rect 6528 5486 6594 5502
rect 8160 5502 8176 5504
rect 8210 5534 8226 5536
rect 9792 5536 9858 5552
rect 9792 5534 9808 5536
rect 8210 5504 9808 5534
rect 8210 5502 8226 5504
rect 8160 5486 8226 5502
rect 9792 5502 9808 5504
rect 9842 5534 9858 5536
rect 11424 5536 11490 5552
rect 11424 5534 11440 5536
rect 9842 5504 11440 5534
rect 9842 5502 9858 5504
rect 9792 5486 9858 5502
rect 11424 5502 11440 5504
rect 11474 5534 11490 5536
rect 13056 5536 13122 5552
rect 13056 5534 13072 5536
rect 11474 5504 13072 5534
rect 11474 5502 11490 5504
rect 11424 5486 11490 5502
rect 13056 5502 13072 5504
rect 13106 5502 13122 5536
rect 13056 5486 13122 5502
rect 0 5332 66 5348
rect 0 5298 16 5332
rect 50 5330 66 5332
rect 1632 5332 1698 5348
rect 1632 5330 1648 5332
rect 50 5300 1648 5330
rect 50 5298 66 5300
rect 0 5282 66 5298
rect 1632 5298 1648 5300
rect 1682 5330 1698 5332
rect 3264 5332 3330 5348
rect 3264 5330 3280 5332
rect 1682 5300 3280 5330
rect 1682 5298 1698 5300
rect 1632 5282 1698 5298
rect 3264 5298 3280 5300
rect 3314 5330 3330 5332
rect 4896 5332 4962 5348
rect 4896 5330 4912 5332
rect 3314 5300 4912 5330
rect 3314 5298 3330 5300
rect 3264 5282 3330 5298
rect 4896 5298 4912 5300
rect 4946 5330 4962 5332
rect 6528 5332 6594 5348
rect 6528 5330 6544 5332
rect 4946 5300 6544 5330
rect 4946 5298 4962 5300
rect 4896 5282 4962 5298
rect 6528 5298 6544 5300
rect 6578 5330 6594 5332
rect 8160 5332 8226 5348
rect 8160 5330 8176 5332
rect 6578 5300 8176 5330
rect 6578 5298 6594 5300
rect 6528 5282 6594 5298
rect 8160 5298 8176 5300
rect 8210 5330 8226 5332
rect 9792 5332 9858 5348
rect 9792 5330 9808 5332
rect 8210 5300 9808 5330
rect 8210 5298 8226 5300
rect 8160 5282 8226 5298
rect 9792 5298 9808 5300
rect 9842 5330 9858 5332
rect 11424 5332 11490 5348
rect 11424 5330 11440 5332
rect 9842 5300 11440 5330
rect 9842 5298 9858 5300
rect 9792 5282 9858 5298
rect 11424 5298 11440 5300
rect 11474 5330 11490 5332
rect 13056 5332 13122 5348
rect 13056 5330 13072 5332
rect 11474 5300 13072 5330
rect 11474 5298 11490 5300
rect 11424 5282 11490 5298
rect 13056 5298 13072 5300
rect 13106 5298 13122 5332
rect 13056 5282 13122 5298
rect 0 5128 66 5144
rect 0 5094 16 5128
rect 50 5126 66 5128
rect 1632 5128 1698 5144
rect 1632 5126 1648 5128
rect 50 5096 1648 5126
rect 50 5094 66 5096
rect 0 5078 66 5094
rect 1632 5094 1648 5096
rect 1682 5126 1698 5128
rect 3264 5128 3330 5144
rect 3264 5126 3280 5128
rect 1682 5096 3280 5126
rect 1682 5094 1698 5096
rect 1632 5078 1698 5094
rect 3264 5094 3280 5096
rect 3314 5126 3330 5128
rect 4896 5128 4962 5144
rect 4896 5126 4912 5128
rect 3314 5096 4912 5126
rect 3314 5094 3330 5096
rect 3264 5078 3330 5094
rect 4896 5094 4912 5096
rect 4946 5126 4962 5128
rect 6528 5128 6594 5144
rect 6528 5126 6544 5128
rect 4946 5096 6544 5126
rect 4946 5094 4962 5096
rect 4896 5078 4962 5094
rect 6528 5094 6544 5096
rect 6578 5126 6594 5128
rect 8160 5128 8226 5144
rect 8160 5126 8176 5128
rect 6578 5096 8176 5126
rect 6578 5094 6594 5096
rect 6528 5078 6594 5094
rect 8160 5094 8176 5096
rect 8210 5126 8226 5128
rect 9792 5128 9858 5144
rect 9792 5126 9808 5128
rect 8210 5096 9808 5126
rect 8210 5094 8226 5096
rect 8160 5078 8226 5094
rect 9792 5094 9808 5096
rect 9842 5126 9858 5128
rect 11424 5128 11490 5144
rect 11424 5126 11440 5128
rect 9842 5096 11440 5126
rect 9842 5094 9858 5096
rect 9792 5078 9858 5094
rect 11424 5094 11440 5096
rect 11474 5126 11490 5128
rect 13056 5128 13122 5144
rect 13056 5126 13072 5128
rect 11474 5096 13072 5126
rect 11474 5094 11490 5096
rect 11424 5078 11490 5094
rect 13056 5094 13072 5096
rect 13106 5094 13122 5128
rect 13056 5078 13122 5094
rect 0 4924 66 4940
rect 0 4890 16 4924
rect 50 4922 66 4924
rect 1632 4924 1698 4940
rect 1632 4922 1648 4924
rect 50 4892 1648 4922
rect 50 4890 66 4892
rect 0 4874 66 4890
rect 1632 4890 1648 4892
rect 1682 4922 1698 4924
rect 3264 4924 3330 4940
rect 3264 4922 3280 4924
rect 1682 4892 3280 4922
rect 1682 4890 1698 4892
rect 1632 4874 1698 4890
rect 3264 4890 3280 4892
rect 3314 4922 3330 4924
rect 4896 4924 4962 4940
rect 4896 4922 4912 4924
rect 3314 4892 4912 4922
rect 3314 4890 3330 4892
rect 3264 4874 3330 4890
rect 4896 4890 4912 4892
rect 4946 4922 4962 4924
rect 6528 4924 6594 4940
rect 6528 4922 6544 4924
rect 4946 4892 6544 4922
rect 4946 4890 4962 4892
rect 4896 4874 4962 4890
rect 6528 4890 6544 4892
rect 6578 4922 6594 4924
rect 8160 4924 8226 4940
rect 8160 4922 8176 4924
rect 6578 4892 8176 4922
rect 6578 4890 6594 4892
rect 6528 4874 6594 4890
rect 8160 4890 8176 4892
rect 8210 4922 8226 4924
rect 9792 4924 9858 4940
rect 9792 4922 9808 4924
rect 8210 4892 9808 4922
rect 8210 4890 8226 4892
rect 8160 4874 8226 4890
rect 9792 4890 9808 4892
rect 9842 4922 9858 4924
rect 11424 4924 11490 4940
rect 11424 4922 11440 4924
rect 9842 4892 11440 4922
rect 9842 4890 9858 4892
rect 9792 4874 9858 4890
rect 11424 4890 11440 4892
rect 11474 4922 11490 4924
rect 13056 4924 13122 4940
rect 13056 4922 13072 4924
rect 11474 4892 13072 4922
rect 11474 4890 11490 4892
rect 11424 4874 11490 4890
rect 13056 4890 13072 4892
rect 13106 4890 13122 4924
rect 13056 4874 13122 4890
rect 0 4720 66 4736
rect 0 4686 16 4720
rect 50 4718 66 4720
rect 1632 4720 1698 4736
rect 1632 4718 1648 4720
rect 50 4688 1648 4718
rect 50 4686 66 4688
rect 0 4670 66 4686
rect 1632 4686 1648 4688
rect 1682 4718 1698 4720
rect 3264 4720 3330 4736
rect 3264 4718 3280 4720
rect 1682 4688 3280 4718
rect 1682 4686 1698 4688
rect 1632 4670 1698 4686
rect 3264 4686 3280 4688
rect 3314 4718 3330 4720
rect 4896 4720 4962 4736
rect 4896 4718 4912 4720
rect 3314 4688 4912 4718
rect 3314 4686 3330 4688
rect 3264 4670 3330 4686
rect 4896 4686 4912 4688
rect 4946 4718 4962 4720
rect 6528 4720 6594 4736
rect 6528 4718 6544 4720
rect 4946 4688 6544 4718
rect 4946 4686 4962 4688
rect 4896 4670 4962 4686
rect 6528 4686 6544 4688
rect 6578 4718 6594 4720
rect 8160 4720 8226 4736
rect 8160 4718 8176 4720
rect 6578 4688 8176 4718
rect 6578 4686 6594 4688
rect 6528 4670 6594 4686
rect 8160 4686 8176 4688
rect 8210 4718 8226 4720
rect 9792 4720 9858 4736
rect 9792 4718 9808 4720
rect 8210 4688 9808 4718
rect 8210 4686 8226 4688
rect 8160 4670 8226 4686
rect 9792 4686 9808 4688
rect 9842 4718 9858 4720
rect 11424 4720 11490 4736
rect 11424 4718 11440 4720
rect 9842 4688 11440 4718
rect 9842 4686 9858 4688
rect 9792 4670 9858 4686
rect 11424 4686 11440 4688
rect 11474 4718 11490 4720
rect 13056 4720 13122 4736
rect 13056 4718 13072 4720
rect 11474 4688 13072 4718
rect 11474 4686 11490 4688
rect 11424 4670 11490 4686
rect 13056 4686 13072 4688
rect 13106 4686 13122 4720
rect 13056 4670 13122 4686
rect 0 4516 66 4532
rect 0 4482 16 4516
rect 50 4514 66 4516
rect 1632 4516 1698 4532
rect 1632 4514 1648 4516
rect 50 4484 1648 4514
rect 50 4482 66 4484
rect 0 4466 66 4482
rect 1632 4482 1648 4484
rect 1682 4514 1698 4516
rect 3264 4516 3330 4532
rect 3264 4514 3280 4516
rect 1682 4484 3280 4514
rect 1682 4482 1698 4484
rect 1632 4466 1698 4482
rect 3264 4482 3280 4484
rect 3314 4514 3330 4516
rect 4896 4516 4962 4532
rect 4896 4514 4912 4516
rect 3314 4484 4912 4514
rect 3314 4482 3330 4484
rect 3264 4466 3330 4482
rect 4896 4482 4912 4484
rect 4946 4514 4962 4516
rect 6528 4516 6594 4532
rect 6528 4514 6544 4516
rect 4946 4484 6544 4514
rect 4946 4482 4962 4484
rect 4896 4466 4962 4482
rect 6528 4482 6544 4484
rect 6578 4514 6594 4516
rect 8160 4516 8226 4532
rect 8160 4514 8176 4516
rect 6578 4484 8176 4514
rect 6578 4482 6594 4484
rect 6528 4466 6594 4482
rect 8160 4482 8176 4484
rect 8210 4514 8226 4516
rect 9792 4516 9858 4532
rect 9792 4514 9808 4516
rect 8210 4484 9808 4514
rect 8210 4482 8226 4484
rect 8160 4466 8226 4482
rect 9792 4482 9808 4484
rect 9842 4514 9858 4516
rect 11424 4516 11490 4532
rect 11424 4514 11440 4516
rect 9842 4484 11440 4514
rect 9842 4482 9858 4484
rect 9792 4466 9858 4482
rect 11424 4482 11440 4484
rect 11474 4514 11490 4516
rect 13056 4516 13122 4532
rect 13056 4514 13072 4516
rect 11474 4484 13072 4514
rect 11474 4482 11490 4484
rect 11424 4466 11490 4482
rect 13056 4482 13072 4484
rect 13106 4482 13122 4516
rect 13056 4466 13122 4482
rect 0 4208 66 4224
rect 0 4174 16 4208
rect 50 4206 66 4208
rect 1632 4208 1698 4224
rect 1632 4206 1648 4208
rect 50 4176 1648 4206
rect 50 4174 66 4176
rect 0 4158 66 4174
rect 1632 4174 1648 4176
rect 1682 4206 1698 4208
rect 3264 4208 3330 4224
rect 3264 4206 3280 4208
rect 1682 4176 3280 4206
rect 1682 4174 1698 4176
rect 1632 4158 1698 4174
rect 3264 4174 3280 4176
rect 3314 4206 3330 4208
rect 4896 4208 4962 4224
rect 4896 4206 4912 4208
rect 3314 4176 4912 4206
rect 3314 4174 3330 4176
rect 3264 4158 3330 4174
rect 4896 4174 4912 4176
rect 4946 4206 4962 4208
rect 6528 4208 6594 4224
rect 6528 4206 6544 4208
rect 4946 4176 6544 4206
rect 4946 4174 4962 4176
rect 4896 4158 4962 4174
rect 6528 4174 6544 4176
rect 6578 4206 6594 4208
rect 8160 4208 8226 4224
rect 8160 4206 8176 4208
rect 6578 4176 8176 4206
rect 6578 4174 6594 4176
rect 6528 4158 6594 4174
rect 8160 4174 8176 4176
rect 8210 4206 8226 4208
rect 9792 4208 9858 4224
rect 9792 4206 9808 4208
rect 8210 4176 9808 4206
rect 8210 4174 8226 4176
rect 8160 4158 8226 4174
rect 9792 4174 9808 4176
rect 9842 4206 9858 4208
rect 11424 4208 11490 4224
rect 11424 4206 11440 4208
rect 9842 4176 11440 4206
rect 9842 4174 9858 4176
rect 9792 4158 9858 4174
rect 11424 4174 11440 4176
rect 11474 4206 11490 4208
rect 13056 4208 13122 4224
rect 13056 4206 13072 4208
rect 11474 4176 13072 4206
rect 11474 4174 11490 4176
rect 11424 4158 11490 4174
rect 13056 4174 13072 4176
rect 13106 4174 13122 4208
rect 13056 4158 13122 4174
rect 0 4004 66 4020
rect 0 3970 16 4004
rect 50 4002 66 4004
rect 1632 4004 1698 4020
rect 1632 4002 1648 4004
rect 50 3972 1648 4002
rect 50 3970 66 3972
rect 0 3954 66 3970
rect 1632 3970 1648 3972
rect 1682 4002 1698 4004
rect 3264 4004 3330 4020
rect 3264 4002 3280 4004
rect 1682 3972 3280 4002
rect 1682 3970 1698 3972
rect 1632 3954 1698 3970
rect 3264 3970 3280 3972
rect 3314 4002 3330 4004
rect 4896 4004 4962 4020
rect 4896 4002 4912 4004
rect 3314 3972 4912 4002
rect 3314 3970 3330 3972
rect 3264 3954 3330 3970
rect 4896 3970 4912 3972
rect 4946 4002 4962 4004
rect 6528 4004 6594 4020
rect 6528 4002 6544 4004
rect 4946 3972 6544 4002
rect 4946 3970 4962 3972
rect 4896 3954 4962 3970
rect 6528 3970 6544 3972
rect 6578 4002 6594 4004
rect 8160 4004 8226 4020
rect 8160 4002 8176 4004
rect 6578 3972 8176 4002
rect 6578 3970 6594 3972
rect 6528 3954 6594 3970
rect 8160 3970 8176 3972
rect 8210 4002 8226 4004
rect 9792 4004 9858 4020
rect 9792 4002 9808 4004
rect 8210 3972 9808 4002
rect 8210 3970 8226 3972
rect 8160 3954 8226 3970
rect 9792 3970 9808 3972
rect 9842 4002 9858 4004
rect 11424 4004 11490 4020
rect 11424 4002 11440 4004
rect 9842 3972 11440 4002
rect 9842 3970 9858 3972
rect 9792 3954 9858 3970
rect 11424 3970 11440 3972
rect 11474 4002 11490 4004
rect 13056 4004 13122 4020
rect 13056 4002 13072 4004
rect 11474 3972 13072 4002
rect 11474 3970 11490 3972
rect 11424 3954 11490 3970
rect 13056 3970 13072 3972
rect 13106 3970 13122 4004
rect 13056 3954 13122 3970
rect 0 3800 66 3816
rect 0 3766 16 3800
rect 50 3798 66 3800
rect 1632 3800 1698 3816
rect 1632 3798 1648 3800
rect 50 3768 1648 3798
rect 50 3766 66 3768
rect 0 3750 66 3766
rect 1632 3766 1648 3768
rect 1682 3798 1698 3800
rect 3264 3800 3330 3816
rect 3264 3798 3280 3800
rect 1682 3768 3280 3798
rect 1682 3766 1698 3768
rect 1632 3750 1698 3766
rect 3264 3766 3280 3768
rect 3314 3798 3330 3800
rect 4896 3800 4962 3816
rect 4896 3798 4912 3800
rect 3314 3768 4912 3798
rect 3314 3766 3330 3768
rect 3264 3750 3330 3766
rect 4896 3766 4912 3768
rect 4946 3798 4962 3800
rect 6528 3800 6594 3816
rect 6528 3798 6544 3800
rect 4946 3768 6544 3798
rect 4946 3766 4962 3768
rect 4896 3750 4962 3766
rect 6528 3766 6544 3768
rect 6578 3798 6594 3800
rect 8160 3800 8226 3816
rect 8160 3798 8176 3800
rect 6578 3768 8176 3798
rect 6578 3766 6594 3768
rect 6528 3750 6594 3766
rect 8160 3766 8176 3768
rect 8210 3798 8226 3800
rect 9792 3800 9858 3816
rect 9792 3798 9808 3800
rect 8210 3768 9808 3798
rect 8210 3766 8226 3768
rect 8160 3750 8226 3766
rect 9792 3766 9808 3768
rect 9842 3798 9858 3800
rect 11424 3800 11490 3816
rect 11424 3798 11440 3800
rect 9842 3768 11440 3798
rect 9842 3766 9858 3768
rect 9792 3750 9858 3766
rect 11424 3766 11440 3768
rect 11474 3798 11490 3800
rect 13056 3800 13122 3816
rect 13056 3798 13072 3800
rect 11474 3768 13072 3798
rect 11474 3766 11490 3768
rect 11424 3750 11490 3766
rect 13056 3766 13072 3768
rect 13106 3766 13122 3800
rect 13056 3750 13122 3766
rect 0 3596 66 3612
rect 0 3562 16 3596
rect 50 3594 66 3596
rect 1632 3596 1698 3612
rect 1632 3594 1648 3596
rect 50 3564 1648 3594
rect 50 3562 66 3564
rect 0 3546 66 3562
rect 1632 3562 1648 3564
rect 1682 3594 1698 3596
rect 3264 3596 3330 3612
rect 3264 3594 3280 3596
rect 1682 3564 3280 3594
rect 1682 3562 1698 3564
rect 1632 3546 1698 3562
rect 3264 3562 3280 3564
rect 3314 3594 3330 3596
rect 4896 3596 4962 3612
rect 4896 3594 4912 3596
rect 3314 3564 4912 3594
rect 3314 3562 3330 3564
rect 3264 3546 3330 3562
rect 4896 3562 4912 3564
rect 4946 3594 4962 3596
rect 6528 3596 6594 3612
rect 6528 3594 6544 3596
rect 4946 3564 6544 3594
rect 4946 3562 4962 3564
rect 4896 3546 4962 3562
rect 6528 3562 6544 3564
rect 6578 3594 6594 3596
rect 8160 3596 8226 3612
rect 8160 3594 8176 3596
rect 6578 3564 8176 3594
rect 6578 3562 6594 3564
rect 6528 3546 6594 3562
rect 8160 3562 8176 3564
rect 8210 3594 8226 3596
rect 9792 3596 9858 3612
rect 9792 3594 9808 3596
rect 8210 3564 9808 3594
rect 8210 3562 8226 3564
rect 8160 3546 8226 3562
rect 9792 3562 9808 3564
rect 9842 3594 9858 3596
rect 11424 3596 11490 3612
rect 11424 3594 11440 3596
rect 9842 3564 11440 3594
rect 9842 3562 9858 3564
rect 9792 3546 9858 3562
rect 11424 3562 11440 3564
rect 11474 3594 11490 3596
rect 13056 3596 13122 3612
rect 13056 3594 13072 3596
rect 11474 3564 13072 3594
rect 11474 3562 11490 3564
rect 11424 3546 11490 3562
rect 13056 3562 13072 3564
rect 13106 3562 13122 3596
rect 13056 3546 13122 3562
rect 0 3392 66 3408
rect 0 3358 16 3392
rect 50 3390 66 3392
rect 1632 3392 1698 3408
rect 1632 3390 1648 3392
rect 50 3360 1648 3390
rect 50 3358 66 3360
rect 0 3342 66 3358
rect 1632 3358 1648 3360
rect 1682 3390 1698 3392
rect 3264 3392 3330 3408
rect 3264 3390 3280 3392
rect 1682 3360 3280 3390
rect 1682 3358 1698 3360
rect 1632 3342 1698 3358
rect 3264 3358 3280 3360
rect 3314 3390 3330 3392
rect 4896 3392 4962 3408
rect 4896 3390 4912 3392
rect 3314 3360 4912 3390
rect 3314 3358 3330 3360
rect 3264 3342 3330 3358
rect 4896 3358 4912 3360
rect 4946 3390 4962 3392
rect 6528 3392 6594 3408
rect 6528 3390 6544 3392
rect 4946 3360 6544 3390
rect 4946 3358 4962 3360
rect 4896 3342 4962 3358
rect 6528 3358 6544 3360
rect 6578 3390 6594 3392
rect 8160 3392 8226 3408
rect 8160 3390 8176 3392
rect 6578 3360 8176 3390
rect 6578 3358 6594 3360
rect 6528 3342 6594 3358
rect 8160 3358 8176 3360
rect 8210 3390 8226 3392
rect 9792 3392 9858 3408
rect 9792 3390 9808 3392
rect 8210 3360 9808 3390
rect 8210 3358 8226 3360
rect 8160 3342 8226 3358
rect 9792 3358 9808 3360
rect 9842 3390 9858 3392
rect 11424 3392 11490 3408
rect 11424 3390 11440 3392
rect 9842 3360 11440 3390
rect 9842 3358 9858 3360
rect 9792 3342 9858 3358
rect 11424 3358 11440 3360
rect 11474 3390 11490 3392
rect 13056 3392 13122 3408
rect 13056 3390 13072 3392
rect 11474 3360 13072 3390
rect 11474 3358 11490 3360
rect 11424 3342 11490 3358
rect 13056 3358 13072 3360
rect 13106 3358 13122 3392
rect 13056 3342 13122 3358
rect 0 3188 66 3204
rect 0 3154 16 3188
rect 50 3186 66 3188
rect 1632 3188 1698 3204
rect 1632 3186 1648 3188
rect 50 3156 1648 3186
rect 50 3154 66 3156
rect 0 3138 66 3154
rect 1632 3154 1648 3156
rect 1682 3186 1698 3188
rect 3264 3188 3330 3204
rect 3264 3186 3280 3188
rect 1682 3156 3280 3186
rect 1682 3154 1698 3156
rect 1632 3138 1698 3154
rect 3264 3154 3280 3156
rect 3314 3186 3330 3188
rect 4896 3188 4962 3204
rect 4896 3186 4912 3188
rect 3314 3156 4912 3186
rect 3314 3154 3330 3156
rect 3264 3138 3330 3154
rect 4896 3154 4912 3156
rect 4946 3186 4962 3188
rect 6528 3188 6594 3204
rect 6528 3186 6544 3188
rect 4946 3156 6544 3186
rect 4946 3154 4962 3156
rect 4896 3138 4962 3154
rect 6528 3154 6544 3156
rect 6578 3186 6594 3188
rect 8160 3188 8226 3204
rect 8160 3186 8176 3188
rect 6578 3156 8176 3186
rect 6578 3154 6594 3156
rect 6528 3138 6594 3154
rect 8160 3154 8176 3156
rect 8210 3186 8226 3188
rect 9792 3188 9858 3204
rect 9792 3186 9808 3188
rect 8210 3156 9808 3186
rect 8210 3154 8226 3156
rect 8160 3138 8226 3154
rect 9792 3154 9808 3156
rect 9842 3186 9858 3188
rect 11424 3188 11490 3204
rect 11424 3186 11440 3188
rect 9842 3156 11440 3186
rect 9842 3154 9858 3156
rect 9792 3138 9858 3154
rect 11424 3154 11440 3156
rect 11474 3186 11490 3188
rect 13056 3188 13122 3204
rect 13056 3186 13072 3188
rect 11474 3156 13072 3186
rect 11474 3154 11490 3156
rect 11424 3138 11490 3154
rect 13056 3154 13072 3156
rect 13106 3154 13122 3188
rect 13056 3138 13122 3154
rect 0 2984 66 3000
rect 0 2950 16 2984
rect 50 2982 66 2984
rect 1632 2984 1698 3000
rect 1632 2982 1648 2984
rect 50 2952 1648 2982
rect 50 2950 66 2952
rect 0 2934 66 2950
rect 1632 2950 1648 2952
rect 1682 2982 1698 2984
rect 3264 2984 3330 3000
rect 3264 2982 3280 2984
rect 1682 2952 3280 2982
rect 1682 2950 1698 2952
rect 1632 2934 1698 2950
rect 3264 2950 3280 2952
rect 3314 2982 3330 2984
rect 4896 2984 4962 3000
rect 4896 2982 4912 2984
rect 3314 2952 4912 2982
rect 3314 2950 3330 2952
rect 3264 2934 3330 2950
rect 4896 2950 4912 2952
rect 4946 2982 4962 2984
rect 6528 2984 6594 3000
rect 6528 2982 6544 2984
rect 4946 2952 6544 2982
rect 4946 2950 4962 2952
rect 4896 2934 4962 2950
rect 6528 2950 6544 2952
rect 6578 2982 6594 2984
rect 8160 2984 8226 3000
rect 8160 2982 8176 2984
rect 6578 2952 8176 2982
rect 6578 2950 6594 2952
rect 6528 2934 6594 2950
rect 8160 2950 8176 2952
rect 8210 2982 8226 2984
rect 9792 2984 9858 3000
rect 9792 2982 9808 2984
rect 8210 2952 9808 2982
rect 8210 2950 8226 2952
rect 8160 2934 8226 2950
rect 9792 2950 9808 2952
rect 9842 2982 9858 2984
rect 11424 2984 11490 3000
rect 11424 2982 11440 2984
rect 9842 2952 11440 2982
rect 9842 2950 9858 2952
rect 9792 2934 9858 2950
rect 11424 2950 11440 2952
rect 11474 2982 11490 2984
rect 13056 2984 13122 3000
rect 13056 2982 13072 2984
rect 11474 2952 13072 2982
rect 11474 2950 11490 2952
rect 11424 2934 11490 2950
rect 13056 2950 13072 2952
rect 13106 2950 13122 2984
rect 13056 2934 13122 2950
rect 0 2780 66 2796
rect 0 2746 16 2780
rect 50 2778 66 2780
rect 1632 2780 1698 2796
rect 1632 2778 1648 2780
rect 50 2748 1648 2778
rect 50 2746 66 2748
rect 0 2730 66 2746
rect 1632 2746 1648 2748
rect 1682 2778 1698 2780
rect 3264 2780 3330 2796
rect 3264 2778 3280 2780
rect 1682 2748 3280 2778
rect 1682 2746 1698 2748
rect 1632 2730 1698 2746
rect 3264 2746 3280 2748
rect 3314 2778 3330 2780
rect 4896 2780 4962 2796
rect 4896 2778 4912 2780
rect 3314 2748 4912 2778
rect 3314 2746 3330 2748
rect 3264 2730 3330 2746
rect 4896 2746 4912 2748
rect 4946 2778 4962 2780
rect 6528 2780 6594 2796
rect 6528 2778 6544 2780
rect 4946 2748 6544 2778
rect 4946 2746 4962 2748
rect 4896 2730 4962 2746
rect 6528 2746 6544 2748
rect 6578 2778 6594 2780
rect 8160 2780 8226 2796
rect 8160 2778 8176 2780
rect 6578 2748 8176 2778
rect 6578 2746 6594 2748
rect 6528 2730 6594 2746
rect 8160 2746 8176 2748
rect 8210 2778 8226 2780
rect 9792 2780 9858 2796
rect 9792 2778 9808 2780
rect 8210 2748 9808 2778
rect 8210 2746 8226 2748
rect 8160 2730 8226 2746
rect 9792 2746 9808 2748
rect 9842 2778 9858 2780
rect 11424 2780 11490 2796
rect 11424 2778 11440 2780
rect 9842 2748 11440 2778
rect 9842 2746 9858 2748
rect 9792 2730 9858 2746
rect 11424 2746 11440 2748
rect 11474 2778 11490 2780
rect 13056 2780 13122 2796
rect 13056 2778 13072 2780
rect 11474 2748 13072 2778
rect 11474 2746 11490 2748
rect 11424 2730 11490 2746
rect 13056 2746 13072 2748
rect 13106 2746 13122 2780
rect 13056 2730 13122 2746
rect 0 2472 66 2488
rect 0 2438 16 2472
rect 50 2470 66 2472
rect 1632 2472 1698 2488
rect 1632 2470 1648 2472
rect 50 2440 1648 2470
rect 50 2438 66 2440
rect 0 2422 66 2438
rect 1632 2438 1648 2440
rect 1682 2470 1698 2472
rect 3264 2472 3330 2488
rect 3264 2470 3280 2472
rect 1682 2440 3280 2470
rect 1682 2438 1698 2440
rect 1632 2422 1698 2438
rect 3264 2438 3280 2440
rect 3314 2470 3330 2472
rect 4896 2472 4962 2488
rect 4896 2470 4912 2472
rect 3314 2440 4912 2470
rect 3314 2438 3330 2440
rect 3264 2422 3330 2438
rect 4896 2438 4912 2440
rect 4946 2470 4962 2472
rect 6528 2472 6594 2488
rect 6528 2470 6544 2472
rect 4946 2440 6544 2470
rect 4946 2438 4962 2440
rect 4896 2422 4962 2438
rect 6528 2438 6544 2440
rect 6578 2470 6594 2472
rect 8160 2472 8226 2488
rect 8160 2470 8176 2472
rect 6578 2440 8176 2470
rect 6578 2438 6594 2440
rect 6528 2422 6594 2438
rect 8160 2438 8176 2440
rect 8210 2470 8226 2472
rect 9792 2472 9858 2488
rect 9792 2470 9808 2472
rect 8210 2440 9808 2470
rect 8210 2438 8226 2440
rect 8160 2422 8226 2438
rect 9792 2438 9808 2440
rect 9842 2470 9858 2472
rect 11424 2472 11490 2488
rect 11424 2470 11440 2472
rect 9842 2440 11440 2470
rect 9842 2438 9858 2440
rect 9792 2422 9858 2438
rect 11424 2438 11440 2440
rect 11474 2470 11490 2472
rect 13056 2472 13122 2488
rect 13056 2470 13072 2472
rect 11474 2440 13072 2470
rect 11474 2438 11490 2440
rect 11424 2422 11490 2438
rect 13056 2438 13072 2440
rect 13106 2438 13122 2472
rect 13056 2422 13122 2438
rect 0 2268 66 2284
rect 0 2234 16 2268
rect 50 2266 66 2268
rect 1632 2268 1698 2284
rect 1632 2266 1648 2268
rect 50 2236 1648 2266
rect 50 2234 66 2236
rect 0 2218 66 2234
rect 1632 2234 1648 2236
rect 1682 2266 1698 2268
rect 3264 2268 3330 2284
rect 3264 2266 3280 2268
rect 1682 2236 3280 2266
rect 1682 2234 1698 2236
rect 1632 2218 1698 2234
rect 3264 2234 3280 2236
rect 3314 2266 3330 2268
rect 4896 2268 4962 2284
rect 4896 2266 4912 2268
rect 3314 2236 4912 2266
rect 3314 2234 3330 2236
rect 3264 2218 3330 2234
rect 4896 2234 4912 2236
rect 4946 2266 4962 2268
rect 6528 2268 6594 2284
rect 6528 2266 6544 2268
rect 4946 2236 6544 2266
rect 4946 2234 4962 2236
rect 4896 2218 4962 2234
rect 6528 2234 6544 2236
rect 6578 2266 6594 2268
rect 8160 2268 8226 2284
rect 8160 2266 8176 2268
rect 6578 2236 8176 2266
rect 6578 2234 6594 2236
rect 6528 2218 6594 2234
rect 8160 2234 8176 2236
rect 8210 2266 8226 2268
rect 9792 2268 9858 2284
rect 9792 2266 9808 2268
rect 8210 2236 9808 2266
rect 8210 2234 8226 2236
rect 8160 2218 8226 2234
rect 9792 2234 9808 2236
rect 9842 2266 9858 2268
rect 11424 2268 11490 2284
rect 11424 2266 11440 2268
rect 9842 2236 11440 2266
rect 9842 2234 9858 2236
rect 9792 2218 9858 2234
rect 11424 2234 11440 2236
rect 11474 2266 11490 2268
rect 13056 2268 13122 2284
rect 13056 2266 13072 2268
rect 11474 2236 13072 2266
rect 11474 2234 11490 2236
rect 11424 2218 11490 2234
rect 13056 2234 13072 2236
rect 13106 2234 13122 2268
rect 13056 2218 13122 2234
rect 0 2064 66 2080
rect 0 2030 16 2064
rect 50 2062 66 2064
rect 1632 2064 1698 2080
rect 1632 2062 1648 2064
rect 50 2032 1648 2062
rect 50 2030 66 2032
rect 0 2014 66 2030
rect 1632 2030 1648 2032
rect 1682 2062 1698 2064
rect 3264 2064 3330 2080
rect 3264 2062 3280 2064
rect 1682 2032 3280 2062
rect 1682 2030 1698 2032
rect 1632 2014 1698 2030
rect 3264 2030 3280 2032
rect 3314 2062 3330 2064
rect 4896 2064 4962 2080
rect 4896 2062 4912 2064
rect 3314 2032 4912 2062
rect 3314 2030 3330 2032
rect 3264 2014 3330 2030
rect 4896 2030 4912 2032
rect 4946 2062 4962 2064
rect 6528 2064 6594 2080
rect 6528 2062 6544 2064
rect 4946 2032 6544 2062
rect 4946 2030 4962 2032
rect 4896 2014 4962 2030
rect 6528 2030 6544 2032
rect 6578 2062 6594 2064
rect 8160 2064 8226 2080
rect 8160 2062 8176 2064
rect 6578 2032 8176 2062
rect 6578 2030 6594 2032
rect 6528 2014 6594 2030
rect 8160 2030 8176 2032
rect 8210 2062 8226 2064
rect 9792 2064 9858 2080
rect 9792 2062 9808 2064
rect 8210 2032 9808 2062
rect 8210 2030 8226 2032
rect 8160 2014 8226 2030
rect 9792 2030 9808 2032
rect 9842 2062 9858 2064
rect 11424 2064 11490 2080
rect 11424 2062 11440 2064
rect 9842 2032 11440 2062
rect 9842 2030 9858 2032
rect 9792 2014 9858 2030
rect 11424 2030 11440 2032
rect 11474 2062 11490 2064
rect 13056 2064 13122 2080
rect 13056 2062 13072 2064
rect 11474 2032 13072 2062
rect 11474 2030 11490 2032
rect 11424 2014 11490 2030
rect 13056 2030 13072 2032
rect 13106 2030 13122 2064
rect 13056 2014 13122 2030
rect 0 1860 66 1876
rect 0 1826 16 1860
rect 50 1858 66 1860
rect 1632 1860 1698 1876
rect 1632 1858 1648 1860
rect 50 1828 1648 1858
rect 50 1826 66 1828
rect 0 1810 66 1826
rect 1632 1826 1648 1828
rect 1682 1858 1698 1860
rect 3264 1860 3330 1876
rect 3264 1858 3280 1860
rect 1682 1828 3280 1858
rect 1682 1826 1698 1828
rect 1632 1810 1698 1826
rect 3264 1826 3280 1828
rect 3314 1858 3330 1860
rect 4896 1860 4962 1876
rect 4896 1858 4912 1860
rect 3314 1828 4912 1858
rect 3314 1826 3330 1828
rect 3264 1810 3330 1826
rect 4896 1826 4912 1828
rect 4946 1858 4962 1860
rect 6528 1860 6594 1876
rect 6528 1858 6544 1860
rect 4946 1828 6544 1858
rect 4946 1826 4962 1828
rect 4896 1810 4962 1826
rect 6528 1826 6544 1828
rect 6578 1858 6594 1860
rect 8160 1860 8226 1876
rect 8160 1858 8176 1860
rect 6578 1828 8176 1858
rect 6578 1826 6594 1828
rect 6528 1810 6594 1826
rect 8160 1826 8176 1828
rect 8210 1858 8226 1860
rect 9792 1860 9858 1876
rect 9792 1858 9808 1860
rect 8210 1828 9808 1858
rect 8210 1826 8226 1828
rect 8160 1810 8226 1826
rect 9792 1826 9808 1828
rect 9842 1858 9858 1860
rect 11424 1860 11490 1876
rect 11424 1858 11440 1860
rect 9842 1828 11440 1858
rect 9842 1826 9858 1828
rect 9792 1810 9858 1826
rect 11424 1826 11440 1828
rect 11474 1858 11490 1860
rect 13056 1860 13122 1876
rect 13056 1858 13072 1860
rect 11474 1828 13072 1858
rect 11474 1826 11490 1828
rect 11424 1810 11490 1826
rect 13056 1826 13072 1828
rect 13106 1826 13122 1860
rect 13056 1810 13122 1826
rect 0 1656 66 1672
rect 0 1622 16 1656
rect 50 1654 66 1656
rect 1632 1656 1698 1672
rect 1632 1654 1648 1656
rect 50 1624 1648 1654
rect 50 1622 66 1624
rect 0 1606 66 1622
rect 1632 1622 1648 1624
rect 1682 1654 1698 1656
rect 3264 1656 3330 1672
rect 3264 1654 3280 1656
rect 1682 1624 3280 1654
rect 1682 1622 1698 1624
rect 1632 1606 1698 1622
rect 3264 1622 3280 1624
rect 3314 1654 3330 1656
rect 4896 1656 4962 1672
rect 4896 1654 4912 1656
rect 3314 1624 4912 1654
rect 3314 1622 3330 1624
rect 3264 1606 3330 1622
rect 4896 1622 4912 1624
rect 4946 1654 4962 1656
rect 6528 1656 6594 1672
rect 6528 1654 6544 1656
rect 4946 1624 6544 1654
rect 4946 1622 4962 1624
rect 4896 1606 4962 1622
rect 6528 1622 6544 1624
rect 6578 1654 6594 1656
rect 8160 1656 8226 1672
rect 8160 1654 8176 1656
rect 6578 1624 8176 1654
rect 6578 1622 6594 1624
rect 6528 1606 6594 1622
rect 8160 1622 8176 1624
rect 8210 1654 8226 1656
rect 9792 1656 9858 1672
rect 9792 1654 9808 1656
rect 8210 1624 9808 1654
rect 8210 1622 8226 1624
rect 8160 1606 8226 1622
rect 9792 1622 9808 1624
rect 9842 1654 9858 1656
rect 11424 1656 11490 1672
rect 11424 1654 11440 1656
rect 9842 1624 11440 1654
rect 9842 1622 9858 1624
rect 9792 1606 9858 1622
rect 11424 1622 11440 1624
rect 11474 1654 11490 1656
rect 13056 1656 13122 1672
rect 13056 1654 13072 1656
rect 11474 1624 13072 1654
rect 11474 1622 11490 1624
rect 11424 1606 11490 1622
rect 13056 1622 13072 1624
rect 13106 1622 13122 1656
rect 13056 1606 13122 1622
rect 0 1452 66 1468
rect 0 1418 16 1452
rect 50 1450 66 1452
rect 1632 1452 1698 1468
rect 1632 1450 1648 1452
rect 50 1420 1648 1450
rect 50 1418 66 1420
rect 0 1402 66 1418
rect 1632 1418 1648 1420
rect 1682 1450 1698 1452
rect 3264 1452 3330 1468
rect 3264 1450 3280 1452
rect 1682 1420 3280 1450
rect 1682 1418 1698 1420
rect 1632 1402 1698 1418
rect 3264 1418 3280 1420
rect 3314 1450 3330 1452
rect 4896 1452 4962 1468
rect 4896 1450 4912 1452
rect 3314 1420 4912 1450
rect 3314 1418 3330 1420
rect 3264 1402 3330 1418
rect 4896 1418 4912 1420
rect 4946 1450 4962 1452
rect 6528 1452 6594 1468
rect 6528 1450 6544 1452
rect 4946 1420 6544 1450
rect 4946 1418 4962 1420
rect 4896 1402 4962 1418
rect 6528 1418 6544 1420
rect 6578 1450 6594 1452
rect 8160 1452 8226 1468
rect 8160 1450 8176 1452
rect 6578 1420 8176 1450
rect 6578 1418 6594 1420
rect 6528 1402 6594 1418
rect 8160 1418 8176 1420
rect 8210 1450 8226 1452
rect 9792 1452 9858 1468
rect 9792 1450 9808 1452
rect 8210 1420 9808 1450
rect 8210 1418 8226 1420
rect 8160 1402 8226 1418
rect 9792 1418 9808 1420
rect 9842 1450 9858 1452
rect 11424 1452 11490 1468
rect 11424 1450 11440 1452
rect 9842 1420 11440 1450
rect 9842 1418 9858 1420
rect 9792 1402 9858 1418
rect 11424 1418 11440 1420
rect 11474 1450 11490 1452
rect 13056 1452 13122 1468
rect 13056 1450 13072 1452
rect 11474 1420 13072 1450
rect 11474 1418 11490 1420
rect 11424 1402 11490 1418
rect 13056 1418 13072 1420
rect 13106 1418 13122 1452
rect 13056 1402 13122 1418
rect 0 1248 66 1264
rect 0 1214 16 1248
rect 50 1246 66 1248
rect 1632 1248 1698 1264
rect 1632 1246 1648 1248
rect 50 1216 1648 1246
rect 50 1214 66 1216
rect 0 1198 66 1214
rect 1632 1214 1648 1216
rect 1682 1246 1698 1248
rect 3264 1248 3330 1264
rect 3264 1246 3280 1248
rect 1682 1216 3280 1246
rect 1682 1214 1698 1216
rect 1632 1198 1698 1214
rect 3264 1214 3280 1216
rect 3314 1246 3330 1248
rect 4896 1248 4962 1264
rect 4896 1246 4912 1248
rect 3314 1216 4912 1246
rect 3314 1214 3330 1216
rect 3264 1198 3330 1214
rect 4896 1214 4912 1216
rect 4946 1246 4962 1248
rect 6528 1248 6594 1264
rect 6528 1246 6544 1248
rect 4946 1216 6544 1246
rect 4946 1214 4962 1216
rect 4896 1198 4962 1214
rect 6528 1214 6544 1216
rect 6578 1246 6594 1248
rect 8160 1248 8226 1264
rect 8160 1246 8176 1248
rect 6578 1216 8176 1246
rect 6578 1214 6594 1216
rect 6528 1198 6594 1214
rect 8160 1214 8176 1216
rect 8210 1246 8226 1248
rect 9792 1248 9858 1264
rect 9792 1246 9808 1248
rect 8210 1216 9808 1246
rect 8210 1214 8226 1216
rect 8160 1198 8226 1214
rect 9792 1214 9808 1216
rect 9842 1246 9858 1248
rect 11424 1248 11490 1264
rect 11424 1246 11440 1248
rect 9842 1216 11440 1246
rect 9842 1214 9858 1216
rect 9792 1198 9858 1214
rect 11424 1214 11440 1216
rect 11474 1246 11490 1248
rect 13056 1248 13122 1264
rect 13056 1246 13072 1248
rect 11474 1216 13072 1246
rect 11474 1214 11490 1216
rect 11424 1198 11490 1214
rect 13056 1214 13072 1216
rect 13106 1214 13122 1248
rect 13056 1198 13122 1214
rect 0 1044 66 1060
rect 0 1010 16 1044
rect 50 1042 66 1044
rect 1632 1044 1698 1060
rect 1632 1042 1648 1044
rect 50 1012 1648 1042
rect 50 1010 66 1012
rect 0 994 66 1010
rect 1632 1010 1648 1012
rect 1682 1042 1698 1044
rect 3264 1044 3330 1060
rect 3264 1042 3280 1044
rect 1682 1012 3280 1042
rect 1682 1010 1698 1012
rect 1632 994 1698 1010
rect 3264 1010 3280 1012
rect 3314 1042 3330 1044
rect 4896 1044 4962 1060
rect 4896 1042 4912 1044
rect 3314 1012 4912 1042
rect 3314 1010 3330 1012
rect 3264 994 3330 1010
rect 4896 1010 4912 1012
rect 4946 1042 4962 1044
rect 6528 1044 6594 1060
rect 6528 1042 6544 1044
rect 4946 1012 6544 1042
rect 4946 1010 4962 1012
rect 4896 994 4962 1010
rect 6528 1010 6544 1012
rect 6578 1042 6594 1044
rect 8160 1044 8226 1060
rect 8160 1042 8176 1044
rect 6578 1012 8176 1042
rect 6578 1010 6594 1012
rect 6528 994 6594 1010
rect 8160 1010 8176 1012
rect 8210 1042 8226 1044
rect 9792 1044 9858 1060
rect 9792 1042 9808 1044
rect 8210 1012 9808 1042
rect 8210 1010 8226 1012
rect 8160 994 8226 1010
rect 9792 1010 9808 1012
rect 9842 1042 9858 1044
rect 11424 1044 11490 1060
rect 11424 1042 11440 1044
rect 9842 1012 11440 1042
rect 9842 1010 9858 1012
rect 9792 994 9858 1010
rect 11424 1010 11440 1012
rect 11474 1042 11490 1044
rect 13056 1044 13122 1060
rect 13056 1042 13072 1044
rect 11474 1012 13072 1042
rect 11474 1010 11490 1012
rect 11424 994 11490 1010
rect 13056 1010 13072 1012
rect 13106 1010 13122 1044
rect 13056 994 13122 1010
<< polycont >>
rect 16 7850 50 7884
rect 1648 7850 1682 7884
rect 3280 7850 3314 7884
rect 4912 7850 4946 7884
rect 6544 7850 6578 7884
rect 8176 7850 8210 7884
rect 9808 7850 9842 7884
rect 11440 7850 11474 7884
rect 13072 7850 13106 7884
rect 16 7646 50 7680
rect 1648 7646 1682 7680
rect 3280 7646 3314 7680
rect 4912 7646 4946 7680
rect 6544 7646 6578 7680
rect 8176 7646 8210 7680
rect 9808 7646 9842 7680
rect 11440 7646 11474 7680
rect 13072 7646 13106 7680
rect 16 7442 50 7476
rect 1648 7442 1682 7476
rect 3280 7442 3314 7476
rect 4912 7442 4946 7476
rect 6544 7442 6578 7476
rect 8176 7442 8210 7476
rect 9808 7442 9842 7476
rect 11440 7442 11474 7476
rect 13072 7442 13106 7476
rect 16 7238 50 7272
rect 1648 7238 1682 7272
rect 3280 7238 3314 7272
rect 4912 7238 4946 7272
rect 6544 7238 6578 7272
rect 8176 7238 8210 7272
rect 9808 7238 9842 7272
rect 11440 7238 11474 7272
rect 13072 7238 13106 7272
rect 16 7034 50 7068
rect 1648 7034 1682 7068
rect 3280 7034 3314 7068
rect 4912 7034 4946 7068
rect 6544 7034 6578 7068
rect 8176 7034 8210 7068
rect 9808 7034 9842 7068
rect 11440 7034 11474 7068
rect 13072 7034 13106 7068
rect 16 6830 50 6864
rect 1648 6830 1682 6864
rect 3280 6830 3314 6864
rect 4912 6830 4946 6864
rect 6544 6830 6578 6864
rect 8176 6830 8210 6864
rect 9808 6830 9842 6864
rect 11440 6830 11474 6864
rect 13072 6830 13106 6864
rect 16 6626 50 6660
rect 1648 6626 1682 6660
rect 3280 6626 3314 6660
rect 4912 6626 4946 6660
rect 6544 6626 6578 6660
rect 8176 6626 8210 6660
rect 9808 6626 9842 6660
rect 11440 6626 11474 6660
rect 13072 6626 13106 6660
rect 16 6422 50 6456
rect 1648 6422 1682 6456
rect 3280 6422 3314 6456
rect 4912 6422 4946 6456
rect 6544 6422 6578 6456
rect 8176 6422 8210 6456
rect 9808 6422 9842 6456
rect 11440 6422 11474 6456
rect 13072 6422 13106 6456
rect 16 6218 50 6252
rect 1648 6218 1682 6252
rect 3280 6218 3314 6252
rect 4912 6218 4946 6252
rect 6544 6218 6578 6252
rect 8176 6218 8210 6252
rect 9808 6218 9842 6252
rect 11440 6218 11474 6252
rect 13072 6218 13106 6252
rect 16 5910 50 5944
rect 1648 5910 1682 5944
rect 3280 5910 3314 5944
rect 4912 5910 4946 5944
rect 6544 5910 6578 5944
rect 8176 5910 8210 5944
rect 9808 5910 9842 5944
rect 11440 5910 11474 5944
rect 13072 5910 13106 5944
rect 16 5706 50 5740
rect 1648 5706 1682 5740
rect 3280 5706 3314 5740
rect 4912 5706 4946 5740
rect 6544 5706 6578 5740
rect 8176 5706 8210 5740
rect 9808 5706 9842 5740
rect 11440 5706 11474 5740
rect 13072 5706 13106 5740
rect 16 5502 50 5536
rect 1648 5502 1682 5536
rect 3280 5502 3314 5536
rect 4912 5502 4946 5536
rect 6544 5502 6578 5536
rect 8176 5502 8210 5536
rect 9808 5502 9842 5536
rect 11440 5502 11474 5536
rect 13072 5502 13106 5536
rect 16 5298 50 5332
rect 1648 5298 1682 5332
rect 3280 5298 3314 5332
rect 4912 5298 4946 5332
rect 6544 5298 6578 5332
rect 8176 5298 8210 5332
rect 9808 5298 9842 5332
rect 11440 5298 11474 5332
rect 13072 5298 13106 5332
rect 16 5094 50 5128
rect 1648 5094 1682 5128
rect 3280 5094 3314 5128
rect 4912 5094 4946 5128
rect 6544 5094 6578 5128
rect 8176 5094 8210 5128
rect 9808 5094 9842 5128
rect 11440 5094 11474 5128
rect 13072 5094 13106 5128
rect 16 4890 50 4924
rect 1648 4890 1682 4924
rect 3280 4890 3314 4924
rect 4912 4890 4946 4924
rect 6544 4890 6578 4924
rect 8176 4890 8210 4924
rect 9808 4890 9842 4924
rect 11440 4890 11474 4924
rect 13072 4890 13106 4924
rect 16 4686 50 4720
rect 1648 4686 1682 4720
rect 3280 4686 3314 4720
rect 4912 4686 4946 4720
rect 6544 4686 6578 4720
rect 8176 4686 8210 4720
rect 9808 4686 9842 4720
rect 11440 4686 11474 4720
rect 13072 4686 13106 4720
rect 16 4482 50 4516
rect 1648 4482 1682 4516
rect 3280 4482 3314 4516
rect 4912 4482 4946 4516
rect 6544 4482 6578 4516
rect 8176 4482 8210 4516
rect 9808 4482 9842 4516
rect 11440 4482 11474 4516
rect 13072 4482 13106 4516
rect 16 4174 50 4208
rect 1648 4174 1682 4208
rect 3280 4174 3314 4208
rect 4912 4174 4946 4208
rect 6544 4174 6578 4208
rect 8176 4174 8210 4208
rect 9808 4174 9842 4208
rect 11440 4174 11474 4208
rect 13072 4174 13106 4208
rect 16 3970 50 4004
rect 1648 3970 1682 4004
rect 3280 3970 3314 4004
rect 4912 3970 4946 4004
rect 6544 3970 6578 4004
rect 8176 3970 8210 4004
rect 9808 3970 9842 4004
rect 11440 3970 11474 4004
rect 13072 3970 13106 4004
rect 16 3766 50 3800
rect 1648 3766 1682 3800
rect 3280 3766 3314 3800
rect 4912 3766 4946 3800
rect 6544 3766 6578 3800
rect 8176 3766 8210 3800
rect 9808 3766 9842 3800
rect 11440 3766 11474 3800
rect 13072 3766 13106 3800
rect 16 3562 50 3596
rect 1648 3562 1682 3596
rect 3280 3562 3314 3596
rect 4912 3562 4946 3596
rect 6544 3562 6578 3596
rect 8176 3562 8210 3596
rect 9808 3562 9842 3596
rect 11440 3562 11474 3596
rect 13072 3562 13106 3596
rect 16 3358 50 3392
rect 1648 3358 1682 3392
rect 3280 3358 3314 3392
rect 4912 3358 4946 3392
rect 6544 3358 6578 3392
rect 8176 3358 8210 3392
rect 9808 3358 9842 3392
rect 11440 3358 11474 3392
rect 13072 3358 13106 3392
rect 16 3154 50 3188
rect 1648 3154 1682 3188
rect 3280 3154 3314 3188
rect 4912 3154 4946 3188
rect 6544 3154 6578 3188
rect 8176 3154 8210 3188
rect 9808 3154 9842 3188
rect 11440 3154 11474 3188
rect 13072 3154 13106 3188
rect 16 2950 50 2984
rect 1648 2950 1682 2984
rect 3280 2950 3314 2984
rect 4912 2950 4946 2984
rect 6544 2950 6578 2984
rect 8176 2950 8210 2984
rect 9808 2950 9842 2984
rect 11440 2950 11474 2984
rect 13072 2950 13106 2984
rect 16 2746 50 2780
rect 1648 2746 1682 2780
rect 3280 2746 3314 2780
rect 4912 2746 4946 2780
rect 6544 2746 6578 2780
rect 8176 2746 8210 2780
rect 9808 2746 9842 2780
rect 11440 2746 11474 2780
rect 13072 2746 13106 2780
rect 16 2438 50 2472
rect 1648 2438 1682 2472
rect 3280 2438 3314 2472
rect 4912 2438 4946 2472
rect 6544 2438 6578 2472
rect 8176 2438 8210 2472
rect 9808 2438 9842 2472
rect 11440 2438 11474 2472
rect 13072 2438 13106 2472
rect 16 2234 50 2268
rect 1648 2234 1682 2268
rect 3280 2234 3314 2268
rect 4912 2234 4946 2268
rect 6544 2234 6578 2268
rect 8176 2234 8210 2268
rect 9808 2234 9842 2268
rect 11440 2234 11474 2268
rect 13072 2234 13106 2268
rect 16 2030 50 2064
rect 1648 2030 1682 2064
rect 3280 2030 3314 2064
rect 4912 2030 4946 2064
rect 6544 2030 6578 2064
rect 8176 2030 8210 2064
rect 9808 2030 9842 2064
rect 11440 2030 11474 2064
rect 13072 2030 13106 2064
rect 16 1826 50 1860
rect 1648 1826 1682 1860
rect 3280 1826 3314 1860
rect 4912 1826 4946 1860
rect 6544 1826 6578 1860
rect 8176 1826 8210 1860
rect 9808 1826 9842 1860
rect 11440 1826 11474 1860
rect 13072 1826 13106 1860
rect 16 1622 50 1656
rect 1648 1622 1682 1656
rect 3280 1622 3314 1656
rect 4912 1622 4946 1656
rect 6544 1622 6578 1656
rect 8176 1622 8210 1656
rect 9808 1622 9842 1656
rect 11440 1622 11474 1656
rect 13072 1622 13106 1656
rect 16 1418 50 1452
rect 1648 1418 1682 1452
rect 3280 1418 3314 1452
rect 4912 1418 4946 1452
rect 6544 1418 6578 1452
rect 8176 1418 8210 1452
rect 9808 1418 9842 1452
rect 11440 1418 11474 1452
rect 13072 1418 13106 1452
rect 16 1214 50 1248
rect 1648 1214 1682 1248
rect 3280 1214 3314 1248
rect 4912 1214 4946 1248
rect 6544 1214 6578 1248
rect 8176 1214 8210 1248
rect 9808 1214 9842 1248
rect 11440 1214 11474 1248
rect 13072 1214 13106 1248
rect 16 1010 50 1044
rect 1648 1010 1682 1044
rect 3280 1010 3314 1044
rect 4912 1010 4946 1044
rect 6544 1010 6578 1044
rect 8176 1010 8210 1044
rect 9808 1010 9842 1044
rect 11440 1010 11474 1044
rect 13072 1010 13106 1044
<< locali >>
rect 16 7884 50 7900
rect 16 7834 50 7850
rect 1648 7884 1682 7900
rect 1648 7834 1682 7850
rect 3280 7884 3314 7900
rect 3280 7834 3314 7850
rect 4912 7884 4946 7900
rect 4912 7834 4946 7850
rect 6544 7884 6578 7900
rect 6544 7834 6578 7850
rect 8176 7884 8210 7900
rect 8176 7834 8210 7850
rect 9808 7884 9842 7900
rect 9808 7834 9842 7850
rect 11440 7884 11474 7900
rect 11440 7834 11474 7850
rect 13072 7884 13106 7900
rect 13072 7834 13106 7850
rect 16 7680 50 7696
rect 16 7630 50 7646
rect 1648 7680 1682 7696
rect 1648 7630 1682 7646
rect 3280 7680 3314 7696
rect 3280 7630 3314 7646
rect 4912 7680 4946 7696
rect 4912 7630 4946 7646
rect 6544 7680 6578 7696
rect 6544 7630 6578 7646
rect 8176 7680 8210 7696
rect 8176 7630 8210 7646
rect 9808 7680 9842 7696
rect 9808 7630 9842 7646
rect 11440 7680 11474 7696
rect 11440 7630 11474 7646
rect 13072 7680 13106 7696
rect 13072 7630 13106 7646
rect 16 7476 50 7492
rect 16 7426 50 7442
rect 1648 7476 1682 7492
rect 1648 7426 1682 7442
rect 3280 7476 3314 7492
rect 3280 7426 3314 7442
rect 4912 7476 4946 7492
rect 4912 7426 4946 7442
rect 6544 7476 6578 7492
rect 6544 7426 6578 7442
rect 8176 7476 8210 7492
rect 8176 7426 8210 7442
rect 9808 7476 9842 7492
rect 9808 7426 9842 7442
rect 11440 7476 11474 7492
rect 11440 7426 11474 7442
rect 13072 7476 13106 7492
rect 13072 7426 13106 7442
rect 16 7272 50 7288
rect 16 7222 50 7238
rect 1648 7272 1682 7288
rect 1648 7222 1682 7238
rect 3280 7272 3314 7288
rect 3280 7222 3314 7238
rect 4912 7272 4946 7288
rect 4912 7222 4946 7238
rect 6544 7272 6578 7288
rect 6544 7222 6578 7238
rect 8176 7272 8210 7288
rect 8176 7222 8210 7238
rect 9808 7272 9842 7288
rect 9808 7222 9842 7238
rect 11440 7272 11474 7288
rect 11440 7222 11474 7238
rect 13072 7272 13106 7288
rect 13072 7222 13106 7238
rect 16 7068 50 7084
rect 16 7018 50 7034
rect 1648 7068 1682 7084
rect 1648 7018 1682 7034
rect 3280 7068 3314 7084
rect 3280 7018 3314 7034
rect 4912 7068 4946 7084
rect 4912 7018 4946 7034
rect 6544 7068 6578 7084
rect 6544 7018 6578 7034
rect 8176 7068 8210 7084
rect 8176 7018 8210 7034
rect 9808 7068 9842 7084
rect 9808 7018 9842 7034
rect 11440 7068 11474 7084
rect 11440 7018 11474 7034
rect 13072 7068 13106 7084
rect 13072 7018 13106 7034
rect 16 6864 50 6880
rect 16 6814 50 6830
rect 1648 6864 1682 6880
rect 1648 6814 1682 6830
rect 3280 6864 3314 6880
rect 3280 6814 3314 6830
rect 4912 6864 4946 6880
rect 4912 6814 4946 6830
rect 6544 6864 6578 6880
rect 6544 6814 6578 6830
rect 8176 6864 8210 6880
rect 8176 6814 8210 6830
rect 9808 6864 9842 6880
rect 9808 6814 9842 6830
rect 11440 6864 11474 6880
rect 11440 6814 11474 6830
rect 13072 6864 13106 6880
rect 13072 6814 13106 6830
rect 16 6660 50 6676
rect 16 6610 50 6626
rect 1648 6660 1682 6676
rect 1648 6610 1682 6626
rect 3280 6660 3314 6676
rect 3280 6610 3314 6626
rect 4912 6660 4946 6676
rect 4912 6610 4946 6626
rect 6544 6660 6578 6676
rect 6544 6610 6578 6626
rect 8176 6660 8210 6676
rect 8176 6610 8210 6626
rect 9808 6660 9842 6676
rect 9808 6610 9842 6626
rect 11440 6660 11474 6676
rect 11440 6610 11474 6626
rect 13072 6660 13106 6676
rect 13072 6610 13106 6626
rect 16 6456 50 6472
rect 16 6406 50 6422
rect 1648 6456 1682 6472
rect 1648 6406 1682 6422
rect 3280 6456 3314 6472
rect 3280 6406 3314 6422
rect 4912 6456 4946 6472
rect 4912 6406 4946 6422
rect 6544 6456 6578 6472
rect 6544 6406 6578 6422
rect 8176 6456 8210 6472
rect 8176 6406 8210 6422
rect 9808 6456 9842 6472
rect 9808 6406 9842 6422
rect 11440 6456 11474 6472
rect 11440 6406 11474 6422
rect 13072 6456 13106 6472
rect 13072 6406 13106 6422
rect 16 6252 50 6268
rect 16 6202 50 6218
rect 1648 6252 1682 6268
rect 1648 6202 1682 6218
rect 3280 6252 3314 6268
rect 3280 6202 3314 6218
rect 4912 6252 4946 6268
rect 4912 6202 4946 6218
rect 6544 6252 6578 6268
rect 6544 6202 6578 6218
rect 8176 6252 8210 6268
rect 8176 6202 8210 6218
rect 9808 6252 9842 6268
rect 9808 6202 9842 6218
rect 11440 6252 11474 6268
rect 11440 6202 11474 6218
rect 13072 6252 13106 6268
rect 13072 6202 13106 6218
rect 211 6064 227 6098
rect 261 6064 277 6098
rect 415 6064 431 6098
rect 465 6064 481 6098
rect 619 6064 635 6098
rect 669 6064 685 6098
rect 823 6064 839 6098
rect 873 6064 889 6098
rect 1027 6064 1043 6098
rect 1077 6064 1093 6098
rect 1231 6064 1247 6098
rect 1281 6064 1297 6098
rect 1435 6064 1451 6098
rect 1485 6064 1501 6098
rect 1639 6064 1655 6098
rect 1689 6064 1705 6098
rect 1843 6064 1859 6098
rect 1893 6064 1909 6098
rect 2047 6064 2063 6098
rect 2097 6064 2113 6098
rect 2251 6064 2267 6098
rect 2301 6064 2317 6098
rect 2455 6064 2471 6098
rect 2505 6064 2521 6098
rect 2659 6064 2675 6098
rect 2709 6064 2725 6098
rect 2863 6064 2879 6098
rect 2913 6064 2929 6098
rect 3067 6064 3083 6098
rect 3117 6064 3133 6098
rect 3271 6064 3287 6098
rect 3321 6064 3337 6098
rect 3475 6064 3491 6098
rect 3525 6064 3541 6098
rect 3679 6064 3695 6098
rect 3729 6064 3745 6098
rect 3883 6064 3899 6098
rect 3933 6064 3949 6098
rect 4087 6064 4103 6098
rect 4137 6064 4153 6098
rect 4291 6064 4307 6098
rect 4341 6064 4357 6098
rect 4495 6064 4511 6098
rect 4545 6064 4561 6098
rect 4699 6064 4715 6098
rect 4749 6064 4765 6098
rect 4903 6064 4919 6098
rect 4953 6064 4969 6098
rect 5107 6064 5123 6098
rect 5157 6064 5173 6098
rect 5311 6064 5327 6098
rect 5361 6064 5377 6098
rect 5515 6064 5531 6098
rect 5565 6064 5581 6098
rect 5719 6064 5735 6098
rect 5769 6064 5785 6098
rect 5923 6064 5939 6098
rect 5973 6064 5989 6098
rect 6127 6064 6143 6098
rect 6177 6064 6193 6098
rect 6331 6064 6347 6098
rect 6381 6064 6397 6098
rect 6535 6064 6551 6098
rect 6585 6064 6601 6098
rect 6739 6064 6755 6098
rect 6789 6064 6805 6098
rect 6943 6064 6959 6098
rect 6993 6064 7009 6098
rect 7147 6064 7163 6098
rect 7197 6064 7213 6098
rect 7351 6064 7367 6098
rect 7401 6064 7417 6098
rect 7555 6064 7571 6098
rect 7605 6064 7621 6098
rect 7759 6064 7775 6098
rect 7809 6064 7825 6098
rect 7963 6064 7979 6098
rect 8013 6064 8029 6098
rect 8167 6064 8183 6098
rect 8217 6064 8233 6098
rect 8371 6064 8387 6098
rect 8421 6064 8437 6098
rect 8575 6064 8591 6098
rect 8625 6064 8641 6098
rect 8779 6064 8795 6098
rect 8829 6064 8845 6098
rect 8983 6064 8999 6098
rect 9033 6064 9049 6098
rect 9187 6064 9203 6098
rect 9237 6064 9253 6098
rect 9391 6064 9407 6098
rect 9441 6064 9457 6098
rect 9595 6064 9611 6098
rect 9645 6064 9661 6098
rect 9799 6064 9815 6098
rect 9849 6064 9865 6098
rect 10003 6064 10019 6098
rect 10053 6064 10069 6098
rect 10207 6064 10223 6098
rect 10257 6064 10273 6098
rect 10411 6064 10427 6098
rect 10461 6064 10477 6098
rect 10615 6064 10631 6098
rect 10665 6064 10681 6098
rect 10819 6064 10835 6098
rect 10869 6064 10885 6098
rect 11023 6064 11039 6098
rect 11073 6064 11089 6098
rect 11227 6064 11243 6098
rect 11277 6064 11293 6098
rect 11431 6064 11447 6098
rect 11481 6064 11497 6098
rect 11635 6064 11651 6098
rect 11685 6064 11701 6098
rect 11839 6064 11855 6098
rect 11889 6064 11905 6098
rect 12043 6064 12059 6098
rect 12093 6064 12109 6098
rect 12247 6064 12263 6098
rect 12297 6064 12313 6098
rect 12451 6064 12467 6098
rect 12501 6064 12517 6098
rect 12655 6064 12671 6098
rect 12705 6064 12721 6098
rect 12859 6064 12875 6098
rect 12909 6064 12925 6098
rect 13077 6064 13093 6098
rect 13127 6064 13143 6098
rect 16 5944 50 5960
rect 16 5894 50 5910
rect 1648 5944 1682 5960
rect 1648 5894 1682 5910
rect 3280 5944 3314 5960
rect 3280 5894 3314 5910
rect 4912 5944 4946 5960
rect 4912 5894 4946 5910
rect 6544 5944 6578 5960
rect 6544 5894 6578 5910
rect 8176 5944 8210 5960
rect 8176 5894 8210 5910
rect 9808 5944 9842 5960
rect 9808 5894 9842 5910
rect 11440 5944 11474 5960
rect 11440 5894 11474 5910
rect 13072 5944 13106 5960
rect 13072 5894 13106 5910
rect 16 5740 50 5756
rect 16 5690 50 5706
rect 1648 5740 1682 5756
rect 1648 5690 1682 5706
rect 3280 5740 3314 5756
rect 3280 5690 3314 5706
rect 4912 5740 4946 5756
rect 4912 5690 4946 5706
rect 6544 5740 6578 5756
rect 6544 5690 6578 5706
rect 8176 5740 8210 5756
rect 8176 5690 8210 5706
rect 9808 5740 9842 5756
rect 9808 5690 9842 5706
rect 11440 5740 11474 5756
rect 11440 5690 11474 5706
rect 13072 5740 13106 5756
rect 13072 5690 13106 5706
rect 16 5536 50 5552
rect 16 5486 50 5502
rect 1648 5536 1682 5552
rect 1648 5486 1682 5502
rect 3280 5536 3314 5552
rect 3280 5486 3314 5502
rect 4912 5536 4946 5552
rect 4912 5486 4946 5502
rect 6544 5536 6578 5552
rect 6544 5486 6578 5502
rect 8176 5536 8210 5552
rect 8176 5486 8210 5502
rect 9808 5536 9842 5552
rect 9808 5486 9842 5502
rect 11440 5536 11474 5552
rect 11440 5486 11474 5502
rect 13072 5536 13106 5552
rect 13072 5486 13106 5502
rect 16 5332 50 5348
rect 16 5282 50 5298
rect 1648 5332 1682 5348
rect 1648 5282 1682 5298
rect 3280 5332 3314 5348
rect 3280 5282 3314 5298
rect 4912 5332 4946 5348
rect 4912 5282 4946 5298
rect 6544 5332 6578 5348
rect 6544 5282 6578 5298
rect 8176 5332 8210 5348
rect 8176 5282 8210 5298
rect 9808 5332 9842 5348
rect 9808 5282 9842 5298
rect 11440 5332 11474 5348
rect 11440 5282 11474 5298
rect 13072 5332 13106 5348
rect 13072 5282 13106 5298
rect 16 5128 50 5144
rect 16 5078 50 5094
rect 1648 5128 1682 5144
rect 1648 5078 1682 5094
rect 3280 5128 3314 5144
rect 3280 5078 3314 5094
rect 4912 5128 4946 5144
rect 4912 5078 4946 5094
rect 6544 5128 6578 5144
rect 6544 5078 6578 5094
rect 8176 5128 8210 5144
rect 8176 5078 8210 5094
rect 9808 5128 9842 5144
rect 9808 5078 9842 5094
rect 11440 5128 11474 5144
rect 11440 5078 11474 5094
rect 13072 5128 13106 5144
rect 13072 5078 13106 5094
rect 16 4924 50 4940
rect 16 4874 50 4890
rect 1648 4924 1682 4940
rect 1648 4874 1682 4890
rect 3280 4924 3314 4940
rect 3280 4874 3314 4890
rect 4912 4924 4946 4940
rect 4912 4874 4946 4890
rect 6544 4924 6578 4940
rect 6544 4874 6578 4890
rect 8176 4924 8210 4940
rect 8176 4874 8210 4890
rect 9808 4924 9842 4940
rect 9808 4874 9842 4890
rect 11440 4924 11474 4940
rect 11440 4874 11474 4890
rect 13072 4924 13106 4940
rect 13072 4874 13106 4890
rect 16 4720 50 4736
rect 16 4670 50 4686
rect 1648 4720 1682 4736
rect 1648 4670 1682 4686
rect 3280 4720 3314 4736
rect 3280 4670 3314 4686
rect 4912 4720 4946 4736
rect 4912 4670 4946 4686
rect 6544 4720 6578 4736
rect 6544 4670 6578 4686
rect 8176 4720 8210 4736
rect 8176 4670 8210 4686
rect 9808 4720 9842 4736
rect 9808 4670 9842 4686
rect 11440 4720 11474 4736
rect 11440 4670 11474 4686
rect 13072 4720 13106 4736
rect 13072 4670 13106 4686
rect 16 4516 50 4532
rect 16 4466 50 4482
rect 1648 4516 1682 4532
rect 1648 4466 1682 4482
rect 3280 4516 3314 4532
rect 3280 4466 3314 4482
rect 4912 4516 4946 4532
rect 4912 4466 4946 4482
rect 6544 4516 6578 4532
rect 6544 4466 6578 4482
rect 8176 4516 8210 4532
rect 8176 4466 8210 4482
rect 9808 4516 9842 4532
rect 9808 4466 9842 4482
rect 11440 4516 11474 4532
rect 11440 4466 11474 4482
rect 13072 4516 13106 4532
rect 13072 4466 13106 4482
rect 211 4328 227 4362
rect 261 4328 277 4362
rect 415 4328 431 4362
rect 465 4328 481 4362
rect 619 4328 635 4362
rect 669 4328 685 4362
rect 823 4328 839 4362
rect 873 4328 889 4362
rect 1027 4328 1043 4362
rect 1077 4328 1093 4362
rect 1231 4328 1247 4362
rect 1281 4328 1297 4362
rect 1435 4328 1451 4362
rect 1485 4328 1501 4362
rect 1639 4328 1655 4362
rect 1689 4328 1705 4362
rect 1843 4328 1859 4362
rect 1893 4328 1909 4362
rect 2047 4328 2063 4362
rect 2097 4328 2113 4362
rect 2251 4328 2267 4362
rect 2301 4328 2317 4362
rect 2455 4328 2471 4362
rect 2505 4328 2521 4362
rect 2659 4328 2675 4362
rect 2709 4328 2725 4362
rect 2863 4328 2879 4362
rect 2913 4328 2929 4362
rect 3067 4328 3083 4362
rect 3117 4328 3133 4362
rect 3271 4328 3287 4362
rect 3321 4328 3337 4362
rect 3475 4328 3491 4362
rect 3525 4328 3541 4362
rect 3679 4328 3695 4362
rect 3729 4328 3745 4362
rect 3883 4328 3899 4362
rect 3933 4328 3949 4362
rect 4087 4328 4103 4362
rect 4137 4328 4153 4362
rect 4291 4328 4307 4362
rect 4341 4328 4357 4362
rect 4495 4328 4511 4362
rect 4545 4328 4561 4362
rect 4699 4328 4715 4362
rect 4749 4328 4765 4362
rect 4903 4328 4919 4362
rect 4953 4328 4969 4362
rect 5107 4328 5123 4362
rect 5157 4328 5173 4362
rect 5311 4328 5327 4362
rect 5361 4328 5377 4362
rect 5515 4328 5531 4362
rect 5565 4328 5581 4362
rect 5719 4328 5735 4362
rect 5769 4328 5785 4362
rect 5923 4328 5939 4362
rect 5973 4328 5989 4362
rect 6127 4328 6143 4362
rect 6177 4328 6193 4362
rect 6331 4328 6347 4362
rect 6381 4328 6397 4362
rect 6535 4328 6551 4362
rect 6585 4328 6601 4362
rect 6739 4328 6755 4362
rect 6789 4328 6805 4362
rect 6943 4328 6959 4362
rect 6993 4328 7009 4362
rect 7147 4328 7163 4362
rect 7197 4328 7213 4362
rect 7351 4328 7367 4362
rect 7401 4328 7417 4362
rect 7555 4328 7571 4362
rect 7605 4328 7621 4362
rect 7759 4328 7775 4362
rect 7809 4328 7825 4362
rect 7963 4328 7979 4362
rect 8013 4328 8029 4362
rect 8167 4328 8183 4362
rect 8217 4328 8233 4362
rect 8371 4328 8387 4362
rect 8421 4328 8437 4362
rect 8575 4328 8591 4362
rect 8625 4328 8641 4362
rect 8779 4328 8795 4362
rect 8829 4328 8845 4362
rect 8983 4328 8999 4362
rect 9033 4328 9049 4362
rect 9187 4328 9203 4362
rect 9237 4328 9253 4362
rect 9391 4328 9407 4362
rect 9441 4328 9457 4362
rect 9595 4328 9611 4362
rect 9645 4328 9661 4362
rect 9799 4328 9815 4362
rect 9849 4328 9865 4362
rect 10003 4328 10019 4362
rect 10053 4328 10069 4362
rect 10207 4328 10223 4362
rect 10257 4328 10273 4362
rect 10411 4328 10427 4362
rect 10461 4328 10477 4362
rect 10615 4328 10631 4362
rect 10665 4328 10681 4362
rect 10819 4328 10835 4362
rect 10869 4328 10885 4362
rect 11023 4328 11039 4362
rect 11073 4328 11089 4362
rect 11227 4328 11243 4362
rect 11277 4328 11293 4362
rect 11431 4328 11447 4362
rect 11481 4328 11497 4362
rect 11635 4328 11651 4362
rect 11685 4328 11701 4362
rect 11839 4328 11855 4362
rect 11889 4328 11905 4362
rect 12043 4328 12059 4362
rect 12093 4328 12109 4362
rect 12247 4328 12263 4362
rect 12297 4328 12313 4362
rect 12451 4328 12467 4362
rect 12501 4328 12517 4362
rect 12655 4328 12671 4362
rect 12705 4328 12721 4362
rect 12859 4328 12875 4362
rect 12909 4328 12925 4362
rect 13077 4328 13093 4362
rect 13127 4328 13143 4362
rect 16 4208 50 4224
rect 16 4158 50 4174
rect 1648 4208 1682 4224
rect 1648 4158 1682 4174
rect 3280 4208 3314 4224
rect 3280 4158 3314 4174
rect 4912 4208 4946 4224
rect 4912 4158 4946 4174
rect 6544 4208 6578 4224
rect 6544 4158 6578 4174
rect 8176 4208 8210 4224
rect 8176 4158 8210 4174
rect 9808 4208 9842 4224
rect 9808 4158 9842 4174
rect 11440 4208 11474 4224
rect 11440 4158 11474 4174
rect 13072 4208 13106 4224
rect 13072 4158 13106 4174
rect 16 4004 50 4020
rect 16 3954 50 3970
rect 1648 4004 1682 4020
rect 1648 3954 1682 3970
rect 3280 4004 3314 4020
rect 3280 3954 3314 3970
rect 4912 4004 4946 4020
rect 4912 3954 4946 3970
rect 6544 4004 6578 4020
rect 6544 3954 6578 3970
rect 8176 4004 8210 4020
rect 8176 3954 8210 3970
rect 9808 4004 9842 4020
rect 9808 3954 9842 3970
rect 11440 4004 11474 4020
rect 11440 3954 11474 3970
rect 13072 4004 13106 4020
rect 13072 3954 13106 3970
rect 16 3800 50 3816
rect 16 3750 50 3766
rect 1648 3800 1682 3816
rect 1648 3750 1682 3766
rect 3280 3800 3314 3816
rect 3280 3750 3314 3766
rect 4912 3800 4946 3816
rect 4912 3750 4946 3766
rect 6544 3800 6578 3816
rect 6544 3750 6578 3766
rect 8176 3800 8210 3816
rect 8176 3750 8210 3766
rect 9808 3800 9842 3816
rect 9808 3750 9842 3766
rect 11440 3800 11474 3816
rect 11440 3750 11474 3766
rect 13072 3800 13106 3816
rect 13072 3750 13106 3766
rect 16 3596 50 3612
rect 16 3546 50 3562
rect 1648 3596 1682 3612
rect 1648 3546 1682 3562
rect 3280 3596 3314 3612
rect 3280 3546 3314 3562
rect 4912 3596 4946 3612
rect 4912 3546 4946 3562
rect 6544 3596 6578 3612
rect 6544 3546 6578 3562
rect 8176 3596 8210 3612
rect 8176 3546 8210 3562
rect 9808 3596 9842 3612
rect 9808 3546 9842 3562
rect 11440 3596 11474 3612
rect 11440 3546 11474 3562
rect 13072 3596 13106 3612
rect 13072 3546 13106 3562
rect 16 3392 50 3408
rect 16 3342 50 3358
rect 1648 3392 1682 3408
rect 1648 3342 1682 3358
rect 3280 3392 3314 3408
rect 3280 3342 3314 3358
rect 4912 3392 4946 3408
rect 4912 3342 4946 3358
rect 6544 3392 6578 3408
rect 6544 3342 6578 3358
rect 8176 3392 8210 3408
rect 8176 3342 8210 3358
rect 9808 3392 9842 3408
rect 9808 3342 9842 3358
rect 11440 3392 11474 3408
rect 11440 3342 11474 3358
rect 13072 3392 13106 3408
rect 13072 3342 13106 3358
rect 16 3188 50 3204
rect 16 3138 50 3154
rect 1648 3188 1682 3204
rect 1648 3138 1682 3154
rect 3280 3188 3314 3204
rect 3280 3138 3314 3154
rect 4912 3188 4946 3204
rect 4912 3138 4946 3154
rect 6544 3188 6578 3204
rect 6544 3138 6578 3154
rect 8176 3188 8210 3204
rect 8176 3138 8210 3154
rect 9808 3188 9842 3204
rect 9808 3138 9842 3154
rect 11440 3188 11474 3204
rect 11440 3138 11474 3154
rect 13072 3188 13106 3204
rect 13072 3138 13106 3154
rect 16 2984 50 3000
rect 16 2934 50 2950
rect 1648 2984 1682 3000
rect 1648 2934 1682 2950
rect 3280 2984 3314 3000
rect 3280 2934 3314 2950
rect 4912 2984 4946 3000
rect 4912 2934 4946 2950
rect 6544 2984 6578 3000
rect 6544 2934 6578 2950
rect 8176 2984 8210 3000
rect 8176 2934 8210 2950
rect 9808 2984 9842 3000
rect 9808 2934 9842 2950
rect 11440 2984 11474 3000
rect 11440 2934 11474 2950
rect 13072 2984 13106 3000
rect 13072 2934 13106 2950
rect 16 2780 50 2796
rect 16 2730 50 2746
rect 1648 2780 1682 2796
rect 1648 2730 1682 2746
rect 3280 2780 3314 2796
rect 3280 2730 3314 2746
rect 4912 2780 4946 2796
rect 4912 2730 4946 2746
rect 6544 2780 6578 2796
rect 6544 2730 6578 2746
rect 8176 2780 8210 2796
rect 8176 2730 8210 2746
rect 9808 2780 9842 2796
rect 9808 2730 9842 2746
rect 11440 2780 11474 2796
rect 11440 2730 11474 2746
rect 13072 2780 13106 2796
rect 13072 2730 13106 2746
rect 211 2592 227 2626
rect 261 2592 277 2626
rect 415 2592 431 2626
rect 465 2592 481 2626
rect 619 2592 635 2626
rect 669 2592 685 2626
rect 823 2592 839 2626
rect 873 2592 889 2626
rect 1027 2592 1043 2626
rect 1077 2592 1093 2626
rect 1231 2592 1247 2626
rect 1281 2592 1297 2626
rect 1435 2592 1451 2626
rect 1485 2592 1501 2626
rect 1639 2592 1655 2626
rect 1689 2592 1705 2626
rect 1843 2592 1859 2626
rect 1893 2592 1909 2626
rect 2047 2592 2063 2626
rect 2097 2592 2113 2626
rect 2251 2592 2267 2626
rect 2301 2592 2317 2626
rect 2455 2592 2471 2626
rect 2505 2592 2521 2626
rect 2659 2592 2675 2626
rect 2709 2592 2725 2626
rect 2863 2592 2879 2626
rect 2913 2592 2929 2626
rect 3067 2592 3083 2626
rect 3117 2592 3133 2626
rect 3271 2592 3287 2626
rect 3321 2592 3337 2626
rect 3475 2592 3491 2626
rect 3525 2592 3541 2626
rect 3679 2592 3695 2626
rect 3729 2592 3745 2626
rect 3883 2592 3899 2626
rect 3933 2592 3949 2626
rect 4087 2592 4103 2626
rect 4137 2592 4153 2626
rect 4291 2592 4307 2626
rect 4341 2592 4357 2626
rect 4495 2592 4511 2626
rect 4545 2592 4561 2626
rect 4699 2592 4715 2626
rect 4749 2592 4765 2626
rect 4903 2592 4919 2626
rect 4953 2592 4969 2626
rect 5107 2592 5123 2626
rect 5157 2592 5173 2626
rect 5311 2592 5327 2626
rect 5361 2592 5377 2626
rect 5515 2592 5531 2626
rect 5565 2592 5581 2626
rect 5719 2592 5735 2626
rect 5769 2592 5785 2626
rect 5923 2592 5939 2626
rect 5973 2592 5989 2626
rect 6127 2592 6143 2626
rect 6177 2592 6193 2626
rect 6331 2592 6347 2626
rect 6381 2592 6397 2626
rect 6535 2592 6551 2626
rect 6585 2592 6601 2626
rect 6739 2592 6755 2626
rect 6789 2592 6805 2626
rect 6943 2592 6959 2626
rect 6993 2592 7009 2626
rect 7147 2592 7163 2626
rect 7197 2592 7213 2626
rect 7351 2592 7367 2626
rect 7401 2592 7417 2626
rect 7555 2592 7571 2626
rect 7605 2592 7621 2626
rect 7759 2592 7775 2626
rect 7809 2592 7825 2626
rect 7963 2592 7979 2626
rect 8013 2592 8029 2626
rect 8167 2592 8183 2626
rect 8217 2592 8233 2626
rect 8371 2592 8387 2626
rect 8421 2592 8437 2626
rect 8575 2592 8591 2626
rect 8625 2592 8641 2626
rect 8779 2592 8795 2626
rect 8829 2592 8845 2626
rect 8983 2592 8999 2626
rect 9033 2592 9049 2626
rect 9187 2592 9203 2626
rect 9237 2592 9253 2626
rect 9391 2592 9407 2626
rect 9441 2592 9457 2626
rect 9595 2592 9611 2626
rect 9645 2592 9661 2626
rect 9799 2592 9815 2626
rect 9849 2592 9865 2626
rect 10003 2592 10019 2626
rect 10053 2592 10069 2626
rect 10207 2592 10223 2626
rect 10257 2592 10273 2626
rect 10411 2592 10427 2626
rect 10461 2592 10477 2626
rect 10615 2592 10631 2626
rect 10665 2592 10681 2626
rect 10819 2592 10835 2626
rect 10869 2592 10885 2626
rect 11023 2592 11039 2626
rect 11073 2592 11089 2626
rect 11227 2592 11243 2626
rect 11277 2592 11293 2626
rect 11431 2592 11447 2626
rect 11481 2592 11497 2626
rect 11635 2592 11651 2626
rect 11685 2592 11701 2626
rect 11839 2592 11855 2626
rect 11889 2592 11905 2626
rect 12043 2592 12059 2626
rect 12093 2592 12109 2626
rect 12247 2592 12263 2626
rect 12297 2592 12313 2626
rect 12451 2592 12467 2626
rect 12501 2592 12517 2626
rect 12655 2592 12671 2626
rect 12705 2592 12721 2626
rect 12859 2592 12875 2626
rect 12909 2592 12925 2626
rect 13077 2592 13093 2626
rect 13127 2592 13143 2626
rect 16 2472 50 2488
rect 16 2422 50 2438
rect 1648 2472 1682 2488
rect 1648 2422 1682 2438
rect 3280 2472 3314 2488
rect 3280 2422 3314 2438
rect 4912 2472 4946 2488
rect 4912 2422 4946 2438
rect 6544 2472 6578 2488
rect 6544 2422 6578 2438
rect 8176 2472 8210 2488
rect 8176 2422 8210 2438
rect 9808 2472 9842 2488
rect 9808 2422 9842 2438
rect 11440 2472 11474 2488
rect 11440 2422 11474 2438
rect 13072 2472 13106 2488
rect 13072 2422 13106 2438
rect 16 2268 50 2284
rect 16 2218 50 2234
rect 1648 2268 1682 2284
rect 1648 2218 1682 2234
rect 3280 2268 3314 2284
rect 3280 2218 3314 2234
rect 4912 2268 4946 2284
rect 4912 2218 4946 2234
rect 6544 2268 6578 2284
rect 6544 2218 6578 2234
rect 8176 2268 8210 2284
rect 8176 2218 8210 2234
rect 9808 2268 9842 2284
rect 9808 2218 9842 2234
rect 11440 2268 11474 2284
rect 11440 2218 11474 2234
rect 13072 2268 13106 2284
rect 13072 2218 13106 2234
rect 16 2064 50 2080
rect 16 2014 50 2030
rect 1648 2064 1682 2080
rect 1648 2014 1682 2030
rect 3280 2064 3314 2080
rect 3280 2014 3314 2030
rect 4912 2064 4946 2080
rect 4912 2014 4946 2030
rect 6544 2064 6578 2080
rect 6544 2014 6578 2030
rect 8176 2064 8210 2080
rect 8176 2014 8210 2030
rect 9808 2064 9842 2080
rect 9808 2014 9842 2030
rect 11440 2064 11474 2080
rect 11440 2014 11474 2030
rect 13072 2064 13106 2080
rect 13072 2014 13106 2030
rect 16 1860 50 1876
rect 16 1810 50 1826
rect 1648 1860 1682 1876
rect 1648 1810 1682 1826
rect 3280 1860 3314 1876
rect 3280 1810 3314 1826
rect 4912 1860 4946 1876
rect 4912 1810 4946 1826
rect 6544 1860 6578 1876
rect 6544 1810 6578 1826
rect 8176 1860 8210 1876
rect 8176 1810 8210 1826
rect 9808 1860 9842 1876
rect 9808 1810 9842 1826
rect 11440 1860 11474 1876
rect 11440 1810 11474 1826
rect 13072 1860 13106 1876
rect 13072 1810 13106 1826
rect 16 1656 50 1672
rect 16 1606 50 1622
rect 1648 1656 1682 1672
rect 1648 1606 1682 1622
rect 3280 1656 3314 1672
rect 3280 1606 3314 1622
rect 4912 1656 4946 1672
rect 4912 1606 4946 1622
rect 6544 1656 6578 1672
rect 6544 1606 6578 1622
rect 8176 1656 8210 1672
rect 8176 1606 8210 1622
rect 9808 1656 9842 1672
rect 9808 1606 9842 1622
rect 11440 1656 11474 1672
rect 11440 1606 11474 1622
rect 13072 1656 13106 1672
rect 13072 1606 13106 1622
rect 16 1452 50 1468
rect 16 1402 50 1418
rect 1648 1452 1682 1468
rect 1648 1402 1682 1418
rect 3280 1452 3314 1468
rect 3280 1402 3314 1418
rect 4912 1452 4946 1468
rect 4912 1402 4946 1418
rect 6544 1452 6578 1468
rect 6544 1402 6578 1418
rect 8176 1452 8210 1468
rect 8176 1402 8210 1418
rect 9808 1452 9842 1468
rect 9808 1402 9842 1418
rect 11440 1452 11474 1468
rect 11440 1402 11474 1418
rect 13072 1452 13106 1468
rect 13072 1402 13106 1418
rect 16 1248 50 1264
rect 16 1198 50 1214
rect 1648 1248 1682 1264
rect 1648 1198 1682 1214
rect 3280 1248 3314 1264
rect 3280 1198 3314 1214
rect 4912 1248 4946 1264
rect 4912 1198 4946 1214
rect 6544 1248 6578 1264
rect 6544 1198 6578 1214
rect 8176 1248 8210 1264
rect 8176 1198 8210 1214
rect 9808 1248 9842 1264
rect 9808 1198 9842 1214
rect 11440 1248 11474 1264
rect 11440 1198 11474 1214
rect 13072 1248 13106 1264
rect 13072 1198 13106 1214
rect 16 1044 50 1060
rect 16 994 50 1010
rect 1648 1044 1682 1060
rect 1648 994 1682 1010
rect 3280 1044 3314 1060
rect 3280 994 3314 1010
rect 4912 1044 4946 1060
rect 4912 994 4946 1010
rect 6544 1044 6578 1060
rect 6544 994 6578 1010
rect 8176 1044 8210 1060
rect 8176 994 8210 1010
rect 9808 1044 9842 1060
rect 9808 994 9842 1010
rect 11440 1044 11474 1060
rect 11440 994 11474 1010
rect 13072 1044 13106 1060
rect 13072 994 13106 1010
rect 211 856 227 890
rect 261 856 277 890
rect 415 856 431 890
rect 465 856 481 890
rect 619 856 635 890
rect 669 856 685 890
rect 823 856 839 890
rect 873 856 889 890
rect 1027 856 1043 890
rect 1077 856 1093 890
rect 1231 856 1247 890
rect 1281 856 1297 890
rect 1435 856 1451 890
rect 1485 856 1501 890
rect 1639 856 1655 890
rect 1689 856 1705 890
rect 1843 856 1859 890
rect 1893 856 1909 890
rect 2047 856 2063 890
rect 2097 856 2113 890
rect 2251 856 2267 890
rect 2301 856 2317 890
rect 2455 856 2471 890
rect 2505 856 2521 890
rect 2659 856 2675 890
rect 2709 856 2725 890
rect 2863 856 2879 890
rect 2913 856 2929 890
rect 3067 856 3083 890
rect 3117 856 3133 890
rect 3271 856 3287 890
rect 3321 856 3337 890
rect 3475 856 3491 890
rect 3525 856 3541 890
rect 3679 856 3695 890
rect 3729 856 3745 890
rect 3883 856 3899 890
rect 3933 856 3949 890
rect 4087 856 4103 890
rect 4137 856 4153 890
rect 4291 856 4307 890
rect 4341 856 4357 890
rect 4495 856 4511 890
rect 4545 856 4561 890
rect 4699 856 4715 890
rect 4749 856 4765 890
rect 4903 856 4919 890
rect 4953 856 4969 890
rect 5107 856 5123 890
rect 5157 856 5173 890
rect 5311 856 5327 890
rect 5361 856 5377 890
rect 5515 856 5531 890
rect 5565 856 5581 890
rect 5719 856 5735 890
rect 5769 856 5785 890
rect 5923 856 5939 890
rect 5973 856 5989 890
rect 6127 856 6143 890
rect 6177 856 6193 890
rect 6331 856 6347 890
rect 6381 856 6397 890
rect 6535 856 6551 890
rect 6585 856 6601 890
rect 6739 856 6755 890
rect 6789 856 6805 890
rect 6943 856 6959 890
rect 6993 856 7009 890
rect 7147 856 7163 890
rect 7197 856 7213 890
rect 7351 856 7367 890
rect 7401 856 7417 890
rect 7555 856 7571 890
rect 7605 856 7621 890
rect 7759 856 7775 890
rect 7809 856 7825 890
rect 7963 856 7979 890
rect 8013 856 8029 890
rect 8167 856 8183 890
rect 8217 856 8233 890
rect 8371 856 8387 890
rect 8421 856 8437 890
rect 8575 856 8591 890
rect 8625 856 8641 890
rect 8779 856 8795 890
rect 8829 856 8845 890
rect 8983 856 8999 890
rect 9033 856 9049 890
rect 9187 856 9203 890
rect 9237 856 9253 890
rect 9391 856 9407 890
rect 9441 856 9457 890
rect 9595 856 9611 890
rect 9645 856 9661 890
rect 9799 856 9815 890
rect 9849 856 9865 890
rect 10003 856 10019 890
rect 10053 856 10069 890
rect 10207 856 10223 890
rect 10257 856 10273 890
rect 10411 856 10427 890
rect 10461 856 10477 890
rect 10615 856 10631 890
rect 10665 856 10681 890
rect 10819 856 10835 890
rect 10869 856 10885 890
rect 11023 856 11039 890
rect 11073 856 11089 890
rect 11227 856 11243 890
rect 11277 856 11293 890
rect 11431 856 11447 890
rect 11481 856 11497 890
rect 11635 856 11651 890
rect 11685 856 11701 890
rect 11839 856 11855 890
rect 11889 856 11905 890
rect 12043 856 12059 890
rect 12093 856 12109 890
rect 12247 856 12263 890
rect 12297 856 12313 890
rect 12451 856 12467 890
rect 12501 856 12517 890
rect 12655 856 12671 890
rect 12705 856 12721 890
rect 12859 856 12875 890
rect 12909 856 12925 890
rect 13077 856 13093 890
rect 13127 856 13143 890
<< viali >>
rect 16 7850 50 7884
rect 1648 7850 1682 7884
rect 3280 7850 3314 7884
rect 4912 7850 4946 7884
rect 6544 7850 6578 7884
rect 8176 7850 8210 7884
rect 9808 7850 9842 7884
rect 11440 7850 11474 7884
rect 13072 7850 13106 7884
rect 16 7646 50 7680
rect 1648 7646 1682 7680
rect 3280 7646 3314 7680
rect 4912 7646 4946 7680
rect 6544 7646 6578 7680
rect 8176 7646 8210 7680
rect 9808 7646 9842 7680
rect 11440 7646 11474 7680
rect 13072 7646 13106 7680
rect 16 7442 50 7476
rect 1648 7442 1682 7476
rect 3280 7442 3314 7476
rect 4912 7442 4946 7476
rect 6544 7442 6578 7476
rect 8176 7442 8210 7476
rect 9808 7442 9842 7476
rect 11440 7442 11474 7476
rect 13072 7442 13106 7476
rect 16 7238 50 7272
rect 1648 7238 1682 7272
rect 3280 7238 3314 7272
rect 4912 7238 4946 7272
rect 6544 7238 6578 7272
rect 8176 7238 8210 7272
rect 9808 7238 9842 7272
rect 11440 7238 11474 7272
rect 13072 7238 13106 7272
rect 16 7034 50 7068
rect 1648 7034 1682 7068
rect 3280 7034 3314 7068
rect 4912 7034 4946 7068
rect 6544 7034 6578 7068
rect 8176 7034 8210 7068
rect 9808 7034 9842 7068
rect 11440 7034 11474 7068
rect 13072 7034 13106 7068
rect 16 6830 50 6864
rect 1648 6830 1682 6864
rect 3280 6830 3314 6864
rect 4912 6830 4946 6864
rect 6544 6830 6578 6864
rect 8176 6830 8210 6864
rect 9808 6830 9842 6864
rect 11440 6830 11474 6864
rect 13072 6830 13106 6864
rect 16 6626 50 6660
rect 1648 6626 1682 6660
rect 3280 6626 3314 6660
rect 4912 6626 4946 6660
rect 6544 6626 6578 6660
rect 8176 6626 8210 6660
rect 9808 6626 9842 6660
rect 11440 6626 11474 6660
rect 13072 6626 13106 6660
rect 16 6422 50 6456
rect 1648 6422 1682 6456
rect 3280 6422 3314 6456
rect 4912 6422 4946 6456
rect 6544 6422 6578 6456
rect 8176 6422 8210 6456
rect 9808 6422 9842 6456
rect 11440 6422 11474 6456
rect 13072 6422 13106 6456
rect 16 6218 50 6252
rect 1648 6218 1682 6252
rect 3280 6218 3314 6252
rect 4912 6218 4946 6252
rect 6544 6218 6578 6252
rect 8176 6218 8210 6252
rect 9808 6218 9842 6252
rect 11440 6218 11474 6252
rect 13072 6218 13106 6252
rect 227 6064 261 6098
rect 431 6064 465 6098
rect 635 6064 669 6098
rect 839 6064 873 6098
rect 1043 6064 1077 6098
rect 1247 6064 1281 6098
rect 1451 6064 1485 6098
rect 1655 6064 1689 6098
rect 1859 6064 1893 6098
rect 2063 6064 2097 6098
rect 2267 6064 2301 6098
rect 2471 6064 2505 6098
rect 2675 6064 2709 6098
rect 2879 6064 2913 6098
rect 3083 6064 3117 6098
rect 3287 6064 3321 6098
rect 3491 6064 3525 6098
rect 3695 6064 3729 6098
rect 3899 6064 3933 6098
rect 4103 6064 4137 6098
rect 4307 6064 4341 6098
rect 4511 6064 4545 6098
rect 4715 6064 4749 6098
rect 4919 6064 4953 6098
rect 5123 6064 5157 6098
rect 5327 6064 5361 6098
rect 5531 6064 5565 6098
rect 5735 6064 5769 6098
rect 5939 6064 5973 6098
rect 6143 6064 6177 6098
rect 6347 6064 6381 6098
rect 6551 6064 6585 6098
rect 6755 6064 6789 6098
rect 6959 6064 6993 6098
rect 7163 6064 7197 6098
rect 7367 6064 7401 6098
rect 7571 6064 7605 6098
rect 7775 6064 7809 6098
rect 7979 6064 8013 6098
rect 8183 6064 8217 6098
rect 8387 6064 8421 6098
rect 8591 6064 8625 6098
rect 8795 6064 8829 6098
rect 8999 6064 9033 6098
rect 9203 6064 9237 6098
rect 9407 6064 9441 6098
rect 9611 6064 9645 6098
rect 9815 6064 9849 6098
rect 10019 6064 10053 6098
rect 10223 6064 10257 6098
rect 10427 6064 10461 6098
rect 10631 6064 10665 6098
rect 10835 6064 10869 6098
rect 11039 6064 11073 6098
rect 11243 6064 11277 6098
rect 11447 6064 11481 6098
rect 11651 6064 11685 6098
rect 11855 6064 11889 6098
rect 12059 6064 12093 6098
rect 12263 6064 12297 6098
rect 12467 6064 12501 6098
rect 12671 6064 12705 6098
rect 12875 6064 12909 6098
rect 13093 6064 13127 6098
rect 16 5910 50 5944
rect 1648 5910 1682 5944
rect 3280 5910 3314 5944
rect 4912 5910 4946 5944
rect 6544 5910 6578 5944
rect 8176 5910 8210 5944
rect 9808 5910 9842 5944
rect 11440 5910 11474 5944
rect 13072 5910 13106 5944
rect 16 5706 50 5740
rect 1648 5706 1682 5740
rect 3280 5706 3314 5740
rect 4912 5706 4946 5740
rect 6544 5706 6578 5740
rect 8176 5706 8210 5740
rect 9808 5706 9842 5740
rect 11440 5706 11474 5740
rect 13072 5706 13106 5740
rect 16 5502 50 5536
rect 1648 5502 1682 5536
rect 3280 5502 3314 5536
rect 4912 5502 4946 5536
rect 6544 5502 6578 5536
rect 8176 5502 8210 5536
rect 9808 5502 9842 5536
rect 11440 5502 11474 5536
rect 13072 5502 13106 5536
rect 16 5298 50 5332
rect 1648 5298 1682 5332
rect 3280 5298 3314 5332
rect 4912 5298 4946 5332
rect 6544 5298 6578 5332
rect 8176 5298 8210 5332
rect 9808 5298 9842 5332
rect 11440 5298 11474 5332
rect 13072 5298 13106 5332
rect 16 5094 50 5128
rect 1648 5094 1682 5128
rect 3280 5094 3314 5128
rect 4912 5094 4946 5128
rect 6544 5094 6578 5128
rect 8176 5094 8210 5128
rect 9808 5094 9842 5128
rect 11440 5094 11474 5128
rect 13072 5094 13106 5128
rect 16 4890 50 4924
rect 1648 4890 1682 4924
rect 3280 4890 3314 4924
rect 4912 4890 4946 4924
rect 6544 4890 6578 4924
rect 8176 4890 8210 4924
rect 9808 4890 9842 4924
rect 11440 4890 11474 4924
rect 13072 4890 13106 4924
rect 16 4686 50 4720
rect 1648 4686 1682 4720
rect 3280 4686 3314 4720
rect 4912 4686 4946 4720
rect 6544 4686 6578 4720
rect 8176 4686 8210 4720
rect 9808 4686 9842 4720
rect 11440 4686 11474 4720
rect 13072 4686 13106 4720
rect 16 4482 50 4516
rect 1648 4482 1682 4516
rect 3280 4482 3314 4516
rect 4912 4482 4946 4516
rect 6544 4482 6578 4516
rect 8176 4482 8210 4516
rect 9808 4482 9842 4516
rect 11440 4482 11474 4516
rect 13072 4482 13106 4516
rect 227 4328 261 4362
rect 431 4328 465 4362
rect 635 4328 669 4362
rect 839 4328 873 4362
rect 1043 4328 1077 4362
rect 1247 4328 1281 4362
rect 1451 4328 1485 4362
rect 1655 4328 1689 4362
rect 1859 4328 1893 4362
rect 2063 4328 2097 4362
rect 2267 4328 2301 4362
rect 2471 4328 2505 4362
rect 2675 4328 2709 4362
rect 2879 4328 2913 4362
rect 3083 4328 3117 4362
rect 3287 4328 3321 4362
rect 3491 4328 3525 4362
rect 3695 4328 3729 4362
rect 3899 4328 3933 4362
rect 4103 4328 4137 4362
rect 4307 4328 4341 4362
rect 4511 4328 4545 4362
rect 4715 4328 4749 4362
rect 4919 4328 4953 4362
rect 5123 4328 5157 4362
rect 5327 4328 5361 4362
rect 5531 4328 5565 4362
rect 5735 4328 5769 4362
rect 5939 4328 5973 4362
rect 6143 4328 6177 4362
rect 6347 4328 6381 4362
rect 6551 4328 6585 4362
rect 6755 4328 6789 4362
rect 6959 4328 6993 4362
rect 7163 4328 7197 4362
rect 7367 4328 7401 4362
rect 7571 4328 7605 4362
rect 7775 4328 7809 4362
rect 7979 4328 8013 4362
rect 8183 4328 8217 4362
rect 8387 4328 8421 4362
rect 8591 4328 8625 4362
rect 8795 4328 8829 4362
rect 8999 4328 9033 4362
rect 9203 4328 9237 4362
rect 9407 4328 9441 4362
rect 9611 4328 9645 4362
rect 9815 4328 9849 4362
rect 10019 4328 10053 4362
rect 10223 4328 10257 4362
rect 10427 4328 10461 4362
rect 10631 4328 10665 4362
rect 10835 4328 10869 4362
rect 11039 4328 11073 4362
rect 11243 4328 11277 4362
rect 11447 4328 11481 4362
rect 11651 4328 11685 4362
rect 11855 4328 11889 4362
rect 12059 4328 12093 4362
rect 12263 4328 12297 4362
rect 12467 4328 12501 4362
rect 12671 4328 12705 4362
rect 12875 4328 12909 4362
rect 13093 4328 13127 4362
rect 16 4174 50 4208
rect 1648 4174 1682 4208
rect 3280 4174 3314 4208
rect 4912 4174 4946 4208
rect 6544 4174 6578 4208
rect 8176 4174 8210 4208
rect 9808 4174 9842 4208
rect 11440 4174 11474 4208
rect 13072 4174 13106 4208
rect 16 3970 50 4004
rect 1648 3970 1682 4004
rect 3280 3970 3314 4004
rect 4912 3970 4946 4004
rect 6544 3970 6578 4004
rect 8176 3970 8210 4004
rect 9808 3970 9842 4004
rect 11440 3970 11474 4004
rect 13072 3970 13106 4004
rect 16 3766 50 3800
rect 1648 3766 1682 3800
rect 3280 3766 3314 3800
rect 4912 3766 4946 3800
rect 6544 3766 6578 3800
rect 8176 3766 8210 3800
rect 9808 3766 9842 3800
rect 11440 3766 11474 3800
rect 13072 3766 13106 3800
rect 16 3562 50 3596
rect 1648 3562 1682 3596
rect 3280 3562 3314 3596
rect 4912 3562 4946 3596
rect 6544 3562 6578 3596
rect 8176 3562 8210 3596
rect 9808 3562 9842 3596
rect 11440 3562 11474 3596
rect 13072 3562 13106 3596
rect 16 3358 50 3392
rect 1648 3358 1682 3392
rect 3280 3358 3314 3392
rect 4912 3358 4946 3392
rect 6544 3358 6578 3392
rect 8176 3358 8210 3392
rect 9808 3358 9842 3392
rect 11440 3358 11474 3392
rect 13072 3358 13106 3392
rect 16 3154 50 3188
rect 1648 3154 1682 3188
rect 3280 3154 3314 3188
rect 4912 3154 4946 3188
rect 6544 3154 6578 3188
rect 8176 3154 8210 3188
rect 9808 3154 9842 3188
rect 11440 3154 11474 3188
rect 13072 3154 13106 3188
rect 16 2950 50 2984
rect 1648 2950 1682 2984
rect 3280 2950 3314 2984
rect 4912 2950 4946 2984
rect 6544 2950 6578 2984
rect 8176 2950 8210 2984
rect 9808 2950 9842 2984
rect 11440 2950 11474 2984
rect 13072 2950 13106 2984
rect 16 2746 50 2780
rect 1648 2746 1682 2780
rect 3280 2746 3314 2780
rect 4912 2746 4946 2780
rect 6544 2746 6578 2780
rect 8176 2746 8210 2780
rect 9808 2746 9842 2780
rect 11440 2746 11474 2780
rect 13072 2746 13106 2780
rect 227 2592 261 2626
rect 431 2592 465 2626
rect 635 2592 669 2626
rect 839 2592 873 2626
rect 1043 2592 1077 2626
rect 1247 2592 1281 2626
rect 1451 2592 1485 2626
rect 1655 2592 1689 2626
rect 1859 2592 1893 2626
rect 2063 2592 2097 2626
rect 2267 2592 2301 2626
rect 2471 2592 2505 2626
rect 2675 2592 2709 2626
rect 2879 2592 2913 2626
rect 3083 2592 3117 2626
rect 3287 2592 3321 2626
rect 3491 2592 3525 2626
rect 3695 2592 3729 2626
rect 3899 2592 3933 2626
rect 4103 2592 4137 2626
rect 4307 2592 4341 2626
rect 4511 2592 4545 2626
rect 4715 2592 4749 2626
rect 4919 2592 4953 2626
rect 5123 2592 5157 2626
rect 5327 2592 5361 2626
rect 5531 2592 5565 2626
rect 5735 2592 5769 2626
rect 5939 2592 5973 2626
rect 6143 2592 6177 2626
rect 6347 2592 6381 2626
rect 6551 2592 6585 2626
rect 6755 2592 6789 2626
rect 6959 2592 6993 2626
rect 7163 2592 7197 2626
rect 7367 2592 7401 2626
rect 7571 2592 7605 2626
rect 7775 2592 7809 2626
rect 7979 2592 8013 2626
rect 8183 2592 8217 2626
rect 8387 2592 8421 2626
rect 8591 2592 8625 2626
rect 8795 2592 8829 2626
rect 8999 2592 9033 2626
rect 9203 2592 9237 2626
rect 9407 2592 9441 2626
rect 9611 2592 9645 2626
rect 9815 2592 9849 2626
rect 10019 2592 10053 2626
rect 10223 2592 10257 2626
rect 10427 2592 10461 2626
rect 10631 2592 10665 2626
rect 10835 2592 10869 2626
rect 11039 2592 11073 2626
rect 11243 2592 11277 2626
rect 11447 2592 11481 2626
rect 11651 2592 11685 2626
rect 11855 2592 11889 2626
rect 12059 2592 12093 2626
rect 12263 2592 12297 2626
rect 12467 2592 12501 2626
rect 12671 2592 12705 2626
rect 12875 2592 12909 2626
rect 13093 2592 13127 2626
rect 16 2438 50 2472
rect 1648 2438 1682 2472
rect 3280 2438 3314 2472
rect 4912 2438 4946 2472
rect 6544 2438 6578 2472
rect 8176 2438 8210 2472
rect 9808 2438 9842 2472
rect 11440 2438 11474 2472
rect 13072 2438 13106 2472
rect 16 2234 50 2268
rect 1648 2234 1682 2268
rect 3280 2234 3314 2268
rect 4912 2234 4946 2268
rect 6544 2234 6578 2268
rect 8176 2234 8210 2268
rect 9808 2234 9842 2268
rect 11440 2234 11474 2268
rect 13072 2234 13106 2268
rect 16 2030 50 2064
rect 1648 2030 1682 2064
rect 3280 2030 3314 2064
rect 4912 2030 4946 2064
rect 6544 2030 6578 2064
rect 8176 2030 8210 2064
rect 9808 2030 9842 2064
rect 11440 2030 11474 2064
rect 13072 2030 13106 2064
rect 16 1826 50 1860
rect 1648 1826 1682 1860
rect 3280 1826 3314 1860
rect 4912 1826 4946 1860
rect 6544 1826 6578 1860
rect 8176 1826 8210 1860
rect 9808 1826 9842 1860
rect 11440 1826 11474 1860
rect 13072 1826 13106 1860
rect 16 1622 50 1656
rect 1648 1622 1682 1656
rect 3280 1622 3314 1656
rect 4912 1622 4946 1656
rect 6544 1622 6578 1656
rect 8176 1622 8210 1656
rect 9808 1622 9842 1656
rect 11440 1622 11474 1656
rect 13072 1622 13106 1656
rect 16 1418 50 1452
rect 1648 1418 1682 1452
rect 3280 1418 3314 1452
rect 4912 1418 4946 1452
rect 6544 1418 6578 1452
rect 8176 1418 8210 1452
rect 9808 1418 9842 1452
rect 11440 1418 11474 1452
rect 13072 1418 13106 1452
rect 16 1214 50 1248
rect 1648 1214 1682 1248
rect 3280 1214 3314 1248
rect 4912 1214 4946 1248
rect 6544 1214 6578 1248
rect 8176 1214 8210 1248
rect 9808 1214 9842 1248
rect 11440 1214 11474 1248
rect 13072 1214 13106 1248
rect 16 1010 50 1044
rect 1648 1010 1682 1044
rect 3280 1010 3314 1044
rect 4912 1010 4946 1044
rect 6544 1010 6578 1044
rect 8176 1010 8210 1044
rect 9808 1010 9842 1044
rect 11440 1010 11474 1044
rect 13072 1010 13106 1044
rect 227 856 261 890
rect 431 856 465 890
rect 635 856 669 890
rect 839 856 873 890
rect 1043 856 1077 890
rect 1247 856 1281 890
rect 1451 856 1485 890
rect 1655 856 1689 890
rect 1859 856 1893 890
rect 2063 856 2097 890
rect 2267 856 2301 890
rect 2471 856 2505 890
rect 2675 856 2709 890
rect 2879 856 2913 890
rect 3083 856 3117 890
rect 3287 856 3321 890
rect 3491 856 3525 890
rect 3695 856 3729 890
rect 3899 856 3933 890
rect 4103 856 4137 890
rect 4307 856 4341 890
rect 4511 856 4545 890
rect 4715 856 4749 890
rect 4919 856 4953 890
rect 5123 856 5157 890
rect 5327 856 5361 890
rect 5531 856 5565 890
rect 5735 856 5769 890
rect 5939 856 5973 890
rect 6143 856 6177 890
rect 6347 856 6381 890
rect 6551 856 6585 890
rect 6755 856 6789 890
rect 6959 856 6993 890
rect 7163 856 7197 890
rect 7367 856 7401 890
rect 7571 856 7605 890
rect 7775 856 7809 890
rect 7979 856 8013 890
rect 8183 856 8217 890
rect 8387 856 8421 890
rect 8591 856 8625 890
rect 8795 856 8829 890
rect 8999 856 9033 890
rect 9203 856 9237 890
rect 9407 856 9441 890
rect 9611 856 9645 890
rect 9815 856 9849 890
rect 10019 856 10053 890
rect 10223 856 10257 890
rect 10427 856 10461 890
rect 10631 856 10665 890
rect 10835 856 10869 890
rect 11039 856 11073 890
rect 11243 856 11277 890
rect 11447 856 11481 890
rect 11651 856 11685 890
rect 11855 856 11889 890
rect 12059 856 12093 890
rect 12263 856 12297 890
rect 12467 856 12501 890
rect 12671 856 12705 890
rect 12875 856 12909 890
rect 13093 856 13127 890
<< metal1 >>
rect 114 7980 13022 8008
rect 8 7893 59 7900
rect 1640 7893 1691 7900
rect 3272 7893 3323 7900
rect 4904 7893 4955 7900
rect 6536 7893 6587 7900
rect 8168 7893 8219 7900
rect 9800 7893 9851 7900
rect 11432 7893 11483 7900
rect 13064 7893 13115 7900
rect 1 7841 7 7893
rect 59 7841 65 7893
rect 1633 7841 1639 7893
rect 1691 7841 1697 7893
rect 3265 7841 3271 7893
rect 3323 7841 3329 7893
rect 4897 7841 4903 7893
rect 4955 7841 4961 7893
rect 6529 7841 6535 7893
rect 6587 7841 6593 7893
rect 8161 7841 8167 7893
rect 8219 7841 8225 7893
rect 9793 7841 9799 7893
rect 9851 7841 9857 7893
rect 11425 7841 11431 7893
rect 11483 7841 11489 7893
rect 13057 7841 13063 7893
rect 13115 7881 13121 7893
rect 13115 7853 13305 7881
rect 13115 7841 13121 7853
rect 8 7834 59 7841
rect 1640 7834 1691 7841
rect 3272 7834 3323 7841
rect 4904 7834 4955 7841
rect 6536 7834 6587 7841
rect 8168 7834 8219 7841
rect 9800 7834 9851 7841
rect 11432 7834 11483 7841
rect 13064 7834 13115 7841
rect 8 7689 59 7696
rect 1640 7689 1691 7696
rect 3272 7689 3323 7696
rect 4904 7689 4955 7696
rect 6536 7689 6587 7696
rect 8168 7689 8219 7696
rect 9800 7689 9851 7696
rect 11432 7689 11483 7696
rect 13064 7689 13115 7696
rect 1 7637 7 7689
rect 59 7637 65 7689
rect 1633 7637 1639 7689
rect 1691 7637 1697 7689
rect 3265 7637 3271 7689
rect 3323 7637 3329 7689
rect 4897 7637 4903 7689
rect 4955 7637 4961 7689
rect 6529 7637 6535 7689
rect 6587 7637 6593 7689
rect 8161 7637 8167 7689
rect 8219 7637 8225 7689
rect 9793 7637 9799 7689
rect 9851 7637 9857 7689
rect 11425 7637 11431 7689
rect 11483 7637 11489 7689
rect 13057 7637 13063 7689
rect 13115 7637 13121 7689
rect 8 7630 59 7637
rect 1640 7630 1691 7637
rect 3272 7630 3323 7637
rect 4904 7630 4955 7637
rect 6536 7630 6587 7637
rect 8168 7630 8219 7637
rect 9800 7630 9851 7637
rect 11432 7630 11483 7637
rect 13064 7630 13115 7637
rect 8 7485 59 7492
rect 1640 7485 1691 7492
rect 3272 7485 3323 7492
rect 4904 7485 4955 7492
rect 6536 7485 6587 7492
rect 8168 7485 8219 7492
rect 9800 7485 9851 7492
rect 11432 7485 11483 7492
rect 13064 7485 13115 7492
rect 1 7433 7 7485
rect 59 7433 65 7485
rect 1633 7433 1639 7485
rect 1691 7433 1697 7485
rect 3265 7433 3271 7485
rect 3323 7433 3329 7485
rect 4897 7433 4903 7485
rect 4955 7433 4961 7485
rect 6529 7433 6535 7485
rect 6587 7433 6593 7485
rect 8161 7433 8167 7485
rect 8219 7433 8225 7485
rect 9793 7433 9799 7485
rect 9851 7433 9857 7485
rect 11425 7433 11431 7485
rect 11483 7433 11489 7485
rect 13057 7433 13063 7485
rect 13115 7433 13121 7485
rect 8 7426 59 7433
rect 1640 7426 1691 7433
rect 3272 7426 3323 7433
rect 4904 7426 4955 7433
rect 6536 7426 6587 7433
rect 8168 7426 8219 7433
rect 9800 7426 9851 7433
rect 11432 7426 11483 7433
rect 13064 7426 13115 7433
rect 8 7281 59 7288
rect 1640 7281 1691 7288
rect 3272 7281 3323 7288
rect 4904 7281 4955 7288
rect 6536 7281 6587 7288
rect 8168 7281 8219 7288
rect 9800 7281 9851 7288
rect 11432 7281 11483 7288
rect 13064 7281 13115 7288
rect 1 7229 7 7281
rect 59 7229 65 7281
rect 1633 7229 1639 7281
rect 1691 7229 1697 7281
rect 3265 7229 3271 7281
rect 3323 7229 3329 7281
rect 4897 7229 4903 7281
rect 4955 7229 4961 7281
rect 6529 7229 6535 7281
rect 6587 7229 6593 7281
rect 8161 7229 8167 7281
rect 8219 7229 8225 7281
rect 9793 7229 9799 7281
rect 9851 7229 9857 7281
rect 11425 7229 11431 7281
rect 11483 7229 11489 7281
rect 13057 7229 13063 7281
rect 13115 7229 13121 7281
rect 8 7222 59 7229
rect 1640 7222 1691 7229
rect 3272 7222 3323 7229
rect 4904 7222 4955 7229
rect 6536 7222 6587 7229
rect 8168 7222 8219 7229
rect 9800 7222 9851 7229
rect 11432 7222 11483 7229
rect 13064 7222 13115 7229
rect 8 7077 59 7084
rect 1640 7077 1691 7084
rect 3272 7077 3323 7084
rect 4904 7077 4955 7084
rect 6536 7077 6587 7084
rect 8168 7077 8219 7084
rect 9800 7077 9851 7084
rect 11432 7077 11483 7084
rect 13064 7077 13115 7084
rect 1 7025 7 7077
rect 59 7025 65 7077
rect 1633 7025 1639 7077
rect 1691 7025 1697 7077
rect 3265 7025 3271 7077
rect 3323 7025 3329 7077
rect 4897 7025 4903 7077
rect 4955 7025 4961 7077
rect 6529 7025 6535 7077
rect 6587 7025 6593 7077
rect 8161 7025 8167 7077
rect 8219 7025 8225 7077
rect 9793 7025 9799 7077
rect 9851 7025 9857 7077
rect 11425 7025 11431 7077
rect 11483 7025 11489 7077
rect 13057 7025 13063 7077
rect 13115 7025 13121 7077
rect 8 7018 59 7025
rect 1640 7018 1691 7025
rect 3272 7018 3323 7025
rect 4904 7018 4955 7025
rect 6536 7018 6587 7025
rect 8168 7018 8219 7025
rect 9800 7018 9851 7025
rect 11432 7018 11483 7025
rect 13064 7018 13115 7025
rect 8 6873 59 6880
rect 1640 6873 1691 6880
rect 3272 6873 3323 6880
rect 4904 6873 4955 6880
rect 6536 6873 6587 6880
rect 8168 6873 8219 6880
rect 9800 6873 9851 6880
rect 11432 6873 11483 6880
rect 13064 6873 13115 6880
rect 1 6821 7 6873
rect 59 6821 65 6873
rect 1633 6821 1639 6873
rect 1691 6821 1697 6873
rect 3265 6821 3271 6873
rect 3323 6821 3329 6873
rect 4897 6821 4903 6873
rect 4955 6821 4961 6873
rect 6529 6821 6535 6873
rect 6587 6821 6593 6873
rect 8161 6821 8167 6873
rect 8219 6821 8225 6873
rect 9793 6821 9799 6873
rect 9851 6821 9857 6873
rect 11425 6821 11431 6873
rect 11483 6821 11489 6873
rect 13057 6821 13063 6873
rect 13115 6821 13121 6873
rect 8 6814 59 6821
rect 1640 6814 1691 6821
rect 3272 6814 3323 6821
rect 4904 6814 4955 6821
rect 6536 6814 6587 6821
rect 8168 6814 8219 6821
rect 9800 6814 9851 6821
rect 11432 6814 11483 6821
rect 13064 6814 13115 6821
rect 8 6669 59 6676
rect 1640 6669 1691 6676
rect 3272 6669 3323 6676
rect 4904 6669 4955 6676
rect 6536 6669 6587 6676
rect 8168 6669 8219 6676
rect 9800 6669 9851 6676
rect 11432 6669 11483 6676
rect 13064 6669 13115 6676
rect 1 6617 7 6669
rect 59 6617 65 6669
rect 1633 6617 1639 6669
rect 1691 6617 1697 6669
rect 3265 6617 3271 6669
rect 3323 6617 3329 6669
rect 4897 6617 4903 6669
rect 4955 6617 4961 6669
rect 6529 6617 6535 6669
rect 6587 6617 6593 6669
rect 8161 6617 8167 6669
rect 8219 6617 8225 6669
rect 9793 6617 9799 6669
rect 9851 6617 9857 6669
rect 11425 6617 11431 6669
rect 11483 6617 11489 6669
rect 13057 6617 13063 6669
rect 13115 6617 13121 6669
rect 8 6610 59 6617
rect 1640 6610 1691 6617
rect 3272 6610 3323 6617
rect 4904 6610 4955 6617
rect 6536 6610 6587 6617
rect 8168 6610 8219 6617
rect 9800 6610 9851 6617
rect 11432 6610 11483 6617
rect 13064 6610 13115 6617
rect 8 6465 59 6472
rect 1640 6465 1691 6472
rect 3272 6465 3323 6472
rect 4904 6465 4955 6472
rect 6536 6465 6587 6472
rect 8168 6465 8219 6472
rect 9800 6465 9851 6472
rect 11432 6465 11483 6472
rect 13064 6465 13115 6472
rect 1 6413 7 6465
rect 59 6413 65 6465
rect 1633 6413 1639 6465
rect 1691 6413 1697 6465
rect 3265 6413 3271 6465
rect 3323 6413 3329 6465
rect 4897 6413 4903 6465
rect 4955 6413 4961 6465
rect 6529 6413 6535 6465
rect 6587 6413 6593 6465
rect 8161 6413 8167 6465
rect 8219 6413 8225 6465
rect 9793 6413 9799 6465
rect 9851 6413 9857 6465
rect 11425 6413 11431 6465
rect 11483 6413 11489 6465
rect 13057 6413 13063 6465
rect 13115 6413 13121 6465
rect 8 6406 59 6413
rect 1640 6406 1691 6413
rect 3272 6406 3323 6413
rect 4904 6406 4955 6413
rect 6536 6406 6587 6413
rect 8168 6406 8219 6413
rect 9800 6406 9851 6413
rect 11432 6406 11483 6413
rect 13064 6406 13115 6413
rect 8 6261 59 6268
rect 1640 6261 1691 6268
rect 3272 6261 3323 6268
rect 4904 6261 4955 6268
rect 6536 6261 6587 6268
rect 8168 6261 8219 6268
rect 9800 6261 9851 6268
rect 11432 6261 11483 6268
rect 13064 6261 13115 6268
rect 1 6209 7 6261
rect 59 6209 65 6261
rect 1633 6209 1639 6261
rect 1691 6209 1697 6261
rect 3265 6209 3271 6261
rect 3323 6209 3329 6261
rect 4897 6209 4903 6261
rect 4955 6209 4961 6261
rect 6529 6209 6535 6261
rect 6587 6209 6593 6261
rect 8161 6209 8167 6261
rect 8219 6209 8225 6261
rect 9793 6209 9799 6261
rect 9851 6209 9857 6261
rect 11425 6209 11431 6261
rect 11483 6209 11489 6261
rect 13057 6209 13063 6261
rect 13115 6209 13121 6261
rect 8 6202 59 6209
rect 1640 6202 1691 6209
rect 3272 6202 3323 6209
rect 4904 6202 4955 6209
rect 6536 6202 6587 6209
rect 8168 6202 8219 6209
rect 9800 6202 9851 6209
rect 11432 6202 11483 6209
rect 13064 6202 13115 6209
rect 128 5977 156 6185
rect 218 6107 270 6113
rect 218 6049 270 6055
rect 332 5977 360 6185
rect 422 6107 474 6113
rect 422 6049 474 6055
rect 536 5977 564 6185
rect 626 6107 678 6113
rect 626 6049 678 6055
rect 740 5977 768 6185
rect 830 6107 882 6113
rect 830 6049 882 6055
rect 944 5977 972 6185
rect 1034 6107 1086 6113
rect 1034 6049 1086 6055
rect 1148 5977 1176 6185
rect 1238 6107 1290 6113
rect 1238 6049 1290 6055
rect 1352 5977 1380 6185
rect 1442 6107 1494 6113
rect 1442 6049 1494 6055
rect 1556 5977 1584 6185
rect 1646 6107 1698 6113
rect 1646 6049 1698 6055
rect 1760 5977 1788 6185
rect 1850 6107 1902 6113
rect 1850 6049 1902 6055
rect 1964 5977 1992 6185
rect 2054 6107 2106 6113
rect 2054 6049 2106 6055
rect 2168 5977 2196 6185
rect 2258 6107 2310 6113
rect 2258 6049 2310 6055
rect 2372 5977 2400 6185
rect 2462 6107 2514 6113
rect 2462 6049 2514 6055
rect 2576 5977 2604 6185
rect 2666 6107 2718 6113
rect 2666 6049 2718 6055
rect 2780 5977 2808 6185
rect 2870 6107 2922 6113
rect 2870 6049 2922 6055
rect 2984 5977 3012 6185
rect 3074 6107 3126 6113
rect 3074 6049 3126 6055
rect 3188 5977 3216 6185
rect 3278 6107 3330 6113
rect 3278 6049 3330 6055
rect 3392 5977 3420 6185
rect 3482 6107 3534 6113
rect 3482 6049 3534 6055
rect 3596 5977 3624 6185
rect 3686 6107 3738 6113
rect 3686 6049 3738 6055
rect 3800 5977 3828 6185
rect 3890 6107 3942 6113
rect 3890 6049 3942 6055
rect 4004 5977 4032 6185
rect 4094 6107 4146 6113
rect 4094 6049 4146 6055
rect 4208 5977 4236 6185
rect 4298 6107 4350 6113
rect 4298 6049 4350 6055
rect 4412 5977 4440 6185
rect 4502 6107 4554 6113
rect 4502 6049 4554 6055
rect 4616 5977 4644 6185
rect 4706 6107 4758 6113
rect 4706 6049 4758 6055
rect 4820 5977 4848 6185
rect 4910 6107 4962 6113
rect 4910 6049 4962 6055
rect 5024 5977 5052 6185
rect 5114 6107 5166 6113
rect 5114 6049 5166 6055
rect 5228 5977 5256 6185
rect 5318 6107 5370 6113
rect 5318 6049 5370 6055
rect 5432 5977 5460 6185
rect 5522 6107 5574 6113
rect 5522 6049 5574 6055
rect 5636 5977 5664 6185
rect 5726 6107 5778 6113
rect 5726 6049 5778 6055
rect 5840 5977 5868 6185
rect 5930 6107 5982 6113
rect 5930 6049 5982 6055
rect 6044 5977 6072 6185
rect 6134 6107 6186 6113
rect 6134 6049 6186 6055
rect 6248 5977 6276 6185
rect 6338 6107 6390 6113
rect 6338 6049 6390 6055
rect 6452 5977 6480 6185
rect 6542 6107 6594 6113
rect 6542 6049 6594 6055
rect 6656 5977 6684 6185
rect 6746 6107 6798 6113
rect 6746 6049 6798 6055
rect 6860 5977 6888 6185
rect 6950 6107 7002 6113
rect 6950 6049 7002 6055
rect 7064 5977 7092 6185
rect 7154 6107 7206 6113
rect 7154 6049 7206 6055
rect 7268 5977 7296 6185
rect 7358 6107 7410 6113
rect 7358 6049 7410 6055
rect 7472 5977 7500 6185
rect 7562 6107 7614 6113
rect 7562 6049 7614 6055
rect 7676 5977 7704 6185
rect 7766 6107 7818 6113
rect 7766 6049 7818 6055
rect 7880 5977 7908 6185
rect 7970 6107 8022 6113
rect 7970 6049 8022 6055
rect 8084 5977 8112 6185
rect 8174 6107 8226 6113
rect 8174 6049 8226 6055
rect 8288 5977 8316 6185
rect 8378 6107 8430 6113
rect 8378 6049 8430 6055
rect 8492 5977 8520 6185
rect 8582 6107 8634 6113
rect 8582 6049 8634 6055
rect 8696 5977 8724 6185
rect 8786 6107 8838 6113
rect 8786 6049 8838 6055
rect 8900 5977 8928 6185
rect 8990 6107 9042 6113
rect 8990 6049 9042 6055
rect 9104 5977 9132 6185
rect 9194 6107 9246 6113
rect 9194 6049 9246 6055
rect 9308 5977 9336 6185
rect 9398 6107 9450 6113
rect 9398 6049 9450 6055
rect 9512 5977 9540 6185
rect 9602 6107 9654 6113
rect 9602 6049 9654 6055
rect 9716 5977 9744 6185
rect 9806 6107 9858 6113
rect 9806 6049 9858 6055
rect 9920 5977 9948 6185
rect 10010 6107 10062 6113
rect 10010 6049 10062 6055
rect 10124 5977 10152 6185
rect 10214 6107 10266 6113
rect 10214 6049 10266 6055
rect 10328 5977 10356 6185
rect 10418 6107 10470 6113
rect 10418 6049 10470 6055
rect 10532 5977 10560 6185
rect 10622 6107 10674 6113
rect 10622 6049 10674 6055
rect 10736 5977 10764 6185
rect 10826 6107 10878 6113
rect 10826 6049 10878 6055
rect 10940 5977 10968 6185
rect 11030 6107 11082 6113
rect 11030 6049 11082 6055
rect 11144 5977 11172 6185
rect 11234 6107 11286 6113
rect 11234 6049 11286 6055
rect 11348 5977 11376 6185
rect 11438 6107 11490 6113
rect 11438 6049 11490 6055
rect 11552 5977 11580 6185
rect 11642 6107 11694 6113
rect 11642 6049 11694 6055
rect 11756 5977 11784 6185
rect 11846 6107 11898 6113
rect 11846 6049 11898 6055
rect 11960 5977 11988 6185
rect 12050 6107 12102 6113
rect 12050 6049 12102 6055
rect 12164 5977 12192 6185
rect 12254 6107 12306 6113
rect 12254 6049 12306 6055
rect 12368 5977 12396 6185
rect 12458 6107 12510 6113
rect 12458 6049 12510 6055
rect 12572 5977 12600 6185
rect 12662 6107 12714 6113
rect 12662 6049 12714 6055
rect 12776 5977 12804 6185
rect 12866 6107 12918 6113
rect 12866 6049 12918 6055
rect 12980 5977 13008 6185
rect 13084 6107 13136 6113
rect 13084 6049 13136 6055
rect 8 5953 59 5960
rect 1640 5953 1691 5960
rect 3272 5953 3323 5960
rect 4904 5953 4955 5960
rect 6536 5953 6587 5960
rect 8168 5953 8219 5960
rect 9800 5953 9851 5960
rect 11432 5953 11483 5960
rect 13064 5953 13115 5960
rect 1 5901 7 5953
rect 59 5901 65 5953
rect 1633 5901 1639 5953
rect 1691 5901 1697 5953
rect 3265 5901 3271 5953
rect 3323 5901 3329 5953
rect 4897 5901 4903 5953
rect 4955 5901 4961 5953
rect 6529 5901 6535 5953
rect 6587 5901 6593 5953
rect 8161 5901 8167 5953
rect 8219 5901 8225 5953
rect 9793 5901 9799 5953
rect 9851 5901 9857 5953
rect 11425 5901 11431 5953
rect 11483 5901 11489 5953
rect 13057 5901 13063 5953
rect 13115 5901 13121 5953
rect 8 5894 59 5901
rect 1640 5894 1691 5901
rect 3272 5894 3323 5901
rect 4904 5894 4955 5901
rect 6536 5894 6587 5901
rect 8168 5894 8219 5901
rect 9800 5894 9851 5901
rect 11432 5894 11483 5901
rect 13064 5894 13115 5901
rect 8 5749 59 5756
rect 1640 5749 1691 5756
rect 3272 5749 3323 5756
rect 4904 5749 4955 5756
rect 6536 5749 6587 5756
rect 8168 5749 8219 5756
rect 9800 5749 9851 5756
rect 11432 5749 11483 5756
rect 13064 5749 13115 5756
rect 1 5697 7 5749
rect 59 5697 65 5749
rect 1633 5697 1639 5749
rect 1691 5697 1697 5749
rect 3265 5697 3271 5749
rect 3323 5697 3329 5749
rect 4897 5697 4903 5749
rect 4955 5697 4961 5749
rect 6529 5697 6535 5749
rect 6587 5697 6593 5749
rect 8161 5697 8167 5749
rect 8219 5697 8225 5749
rect 9793 5697 9799 5749
rect 9851 5697 9857 5749
rect 11425 5697 11431 5749
rect 11483 5697 11489 5749
rect 13057 5697 13063 5749
rect 13115 5697 13121 5749
rect 8 5690 59 5697
rect 1640 5690 1691 5697
rect 3272 5690 3323 5697
rect 4904 5690 4955 5697
rect 6536 5690 6587 5697
rect 8168 5690 8219 5697
rect 9800 5690 9851 5697
rect 11432 5690 11483 5697
rect 13064 5690 13115 5697
rect 8 5545 59 5552
rect 1640 5545 1691 5552
rect 3272 5545 3323 5552
rect 4904 5545 4955 5552
rect 6536 5545 6587 5552
rect 8168 5545 8219 5552
rect 9800 5545 9851 5552
rect 11432 5545 11483 5552
rect 13064 5545 13115 5552
rect 1 5493 7 5545
rect 59 5493 65 5545
rect 1633 5493 1639 5545
rect 1691 5493 1697 5545
rect 3265 5493 3271 5545
rect 3323 5493 3329 5545
rect 4897 5493 4903 5545
rect 4955 5493 4961 5545
rect 6529 5493 6535 5545
rect 6587 5493 6593 5545
rect 8161 5493 8167 5545
rect 8219 5493 8225 5545
rect 9793 5493 9799 5545
rect 9851 5493 9857 5545
rect 11425 5493 11431 5545
rect 11483 5493 11489 5545
rect 13057 5493 13063 5545
rect 13115 5493 13121 5545
rect 8 5486 59 5493
rect 1640 5486 1691 5493
rect 3272 5486 3323 5493
rect 4904 5486 4955 5493
rect 6536 5486 6587 5493
rect 8168 5486 8219 5493
rect 9800 5486 9851 5493
rect 11432 5486 11483 5493
rect 13064 5486 13115 5493
rect 8 5341 59 5348
rect 1640 5341 1691 5348
rect 3272 5341 3323 5348
rect 4904 5341 4955 5348
rect 6536 5341 6587 5348
rect 8168 5341 8219 5348
rect 9800 5341 9851 5348
rect 11432 5341 11483 5348
rect 13064 5341 13115 5348
rect 1 5289 7 5341
rect 59 5289 65 5341
rect 1633 5289 1639 5341
rect 1691 5289 1697 5341
rect 3265 5289 3271 5341
rect 3323 5289 3329 5341
rect 4897 5289 4903 5341
rect 4955 5289 4961 5341
rect 6529 5289 6535 5341
rect 6587 5289 6593 5341
rect 8161 5289 8167 5341
rect 8219 5289 8225 5341
rect 9793 5289 9799 5341
rect 9851 5289 9857 5341
rect 11425 5289 11431 5341
rect 11483 5289 11489 5341
rect 13057 5289 13063 5341
rect 13115 5289 13121 5341
rect 8 5282 59 5289
rect 1640 5282 1691 5289
rect 3272 5282 3323 5289
rect 4904 5282 4955 5289
rect 6536 5282 6587 5289
rect 8168 5282 8219 5289
rect 9800 5282 9851 5289
rect 11432 5282 11483 5289
rect 13064 5282 13115 5289
rect 8 5137 59 5144
rect 1640 5137 1691 5144
rect 3272 5137 3323 5144
rect 4904 5137 4955 5144
rect 6536 5137 6587 5144
rect 8168 5137 8219 5144
rect 9800 5137 9851 5144
rect 11432 5137 11483 5144
rect 13064 5137 13115 5144
rect 1 5085 7 5137
rect 59 5085 65 5137
rect 1633 5085 1639 5137
rect 1691 5085 1697 5137
rect 3265 5085 3271 5137
rect 3323 5085 3329 5137
rect 4897 5085 4903 5137
rect 4955 5085 4961 5137
rect 6529 5085 6535 5137
rect 6587 5085 6593 5137
rect 8161 5085 8167 5137
rect 8219 5085 8225 5137
rect 9793 5085 9799 5137
rect 9851 5085 9857 5137
rect 11425 5085 11431 5137
rect 11483 5085 11489 5137
rect 13057 5085 13063 5137
rect 13115 5085 13121 5137
rect 8 5078 59 5085
rect 1640 5078 1691 5085
rect 3272 5078 3323 5085
rect 4904 5078 4955 5085
rect 6536 5078 6587 5085
rect 8168 5078 8219 5085
rect 9800 5078 9851 5085
rect 11432 5078 11483 5085
rect 13064 5078 13115 5085
rect 8 4933 59 4940
rect 1640 4933 1691 4940
rect 3272 4933 3323 4940
rect 4904 4933 4955 4940
rect 6536 4933 6587 4940
rect 8168 4933 8219 4940
rect 9800 4933 9851 4940
rect 11432 4933 11483 4940
rect 13064 4933 13115 4940
rect 1 4881 7 4933
rect 59 4881 65 4933
rect 1633 4881 1639 4933
rect 1691 4881 1697 4933
rect 3265 4881 3271 4933
rect 3323 4881 3329 4933
rect 4897 4881 4903 4933
rect 4955 4881 4961 4933
rect 6529 4881 6535 4933
rect 6587 4881 6593 4933
rect 8161 4881 8167 4933
rect 8219 4881 8225 4933
rect 9793 4881 9799 4933
rect 9851 4881 9857 4933
rect 11425 4881 11431 4933
rect 11483 4881 11489 4933
rect 13057 4881 13063 4933
rect 13115 4881 13121 4933
rect 8 4874 59 4881
rect 1640 4874 1691 4881
rect 3272 4874 3323 4881
rect 4904 4874 4955 4881
rect 6536 4874 6587 4881
rect 8168 4874 8219 4881
rect 9800 4874 9851 4881
rect 11432 4874 11483 4881
rect 13064 4874 13115 4881
rect 8 4729 59 4736
rect 1640 4729 1691 4736
rect 3272 4729 3323 4736
rect 4904 4729 4955 4736
rect 6536 4729 6587 4736
rect 8168 4729 8219 4736
rect 9800 4729 9851 4736
rect 11432 4729 11483 4736
rect 13064 4729 13115 4736
rect 1 4677 7 4729
rect 59 4677 65 4729
rect 1633 4677 1639 4729
rect 1691 4677 1697 4729
rect 3265 4677 3271 4729
rect 3323 4677 3329 4729
rect 4897 4677 4903 4729
rect 4955 4677 4961 4729
rect 6529 4677 6535 4729
rect 6587 4677 6593 4729
rect 8161 4677 8167 4729
rect 8219 4677 8225 4729
rect 9793 4677 9799 4729
rect 9851 4677 9857 4729
rect 11425 4677 11431 4729
rect 11483 4677 11489 4729
rect 13057 4677 13063 4729
rect 13115 4677 13121 4729
rect 8 4670 59 4677
rect 1640 4670 1691 4677
rect 3272 4670 3323 4677
rect 4904 4670 4955 4677
rect 6536 4670 6587 4677
rect 8168 4670 8219 4677
rect 9800 4670 9851 4677
rect 11432 4670 11483 4677
rect 13064 4670 13115 4677
rect 8 4525 59 4532
rect 1640 4525 1691 4532
rect 3272 4525 3323 4532
rect 4904 4525 4955 4532
rect 6536 4525 6587 4532
rect 8168 4525 8219 4532
rect 9800 4525 9851 4532
rect 11432 4525 11483 4532
rect 13064 4525 13115 4532
rect 1 4473 7 4525
rect 59 4473 65 4525
rect 1633 4473 1639 4525
rect 1691 4473 1697 4525
rect 3265 4473 3271 4525
rect 3323 4473 3329 4525
rect 4897 4473 4903 4525
rect 4955 4473 4961 4525
rect 6529 4473 6535 4525
rect 6587 4473 6593 4525
rect 8161 4473 8167 4525
rect 8219 4473 8225 4525
rect 9793 4473 9799 4525
rect 9851 4473 9857 4525
rect 11425 4473 11431 4525
rect 11483 4473 11489 4525
rect 13057 4473 13063 4525
rect 13115 4473 13121 4525
rect 8 4466 59 4473
rect 1640 4466 1691 4473
rect 3272 4466 3323 4473
rect 4904 4466 4955 4473
rect 6536 4466 6587 4473
rect 8168 4466 8219 4473
rect 9800 4466 9851 4473
rect 11432 4466 11483 4473
rect 13064 4466 13115 4473
rect 128 4241 156 4449
rect 218 4371 270 4377
rect 218 4313 270 4319
rect 332 4241 360 4449
rect 422 4371 474 4377
rect 422 4313 474 4319
rect 536 4241 564 4449
rect 626 4371 678 4377
rect 626 4313 678 4319
rect 740 4241 768 4449
rect 830 4371 882 4377
rect 830 4313 882 4319
rect 944 4241 972 4449
rect 1034 4371 1086 4377
rect 1034 4313 1086 4319
rect 1148 4241 1176 4449
rect 1238 4371 1290 4377
rect 1238 4313 1290 4319
rect 1352 4241 1380 4449
rect 1442 4371 1494 4377
rect 1442 4313 1494 4319
rect 1556 4241 1584 4449
rect 1646 4371 1698 4377
rect 1646 4313 1698 4319
rect 1760 4241 1788 4449
rect 1850 4371 1902 4377
rect 1850 4313 1902 4319
rect 1964 4241 1992 4449
rect 2054 4371 2106 4377
rect 2054 4313 2106 4319
rect 2168 4241 2196 4449
rect 2258 4371 2310 4377
rect 2258 4313 2310 4319
rect 2372 4241 2400 4449
rect 2462 4371 2514 4377
rect 2462 4313 2514 4319
rect 2576 4241 2604 4449
rect 2666 4371 2718 4377
rect 2666 4313 2718 4319
rect 2780 4241 2808 4449
rect 2870 4371 2922 4377
rect 2870 4313 2922 4319
rect 2984 4241 3012 4449
rect 3074 4371 3126 4377
rect 3074 4313 3126 4319
rect 3188 4241 3216 4449
rect 3278 4371 3330 4377
rect 3278 4313 3330 4319
rect 3392 4241 3420 4449
rect 3482 4371 3534 4377
rect 3482 4313 3534 4319
rect 3596 4241 3624 4449
rect 3686 4371 3738 4377
rect 3686 4313 3738 4319
rect 3800 4241 3828 4449
rect 3890 4371 3942 4377
rect 3890 4313 3942 4319
rect 4004 4241 4032 4449
rect 4094 4371 4146 4377
rect 4094 4313 4146 4319
rect 4208 4241 4236 4449
rect 4298 4371 4350 4377
rect 4298 4313 4350 4319
rect 4412 4241 4440 4449
rect 4502 4371 4554 4377
rect 4502 4313 4554 4319
rect 4616 4241 4644 4449
rect 4706 4371 4758 4377
rect 4706 4313 4758 4319
rect 4820 4241 4848 4449
rect 4910 4371 4962 4377
rect 4910 4313 4962 4319
rect 5024 4241 5052 4449
rect 5114 4371 5166 4377
rect 5114 4313 5166 4319
rect 5228 4241 5256 4449
rect 5318 4371 5370 4377
rect 5318 4313 5370 4319
rect 5432 4241 5460 4449
rect 5522 4371 5574 4377
rect 5522 4313 5574 4319
rect 5636 4241 5664 4449
rect 5726 4371 5778 4377
rect 5726 4313 5778 4319
rect 5840 4241 5868 4449
rect 5930 4371 5982 4377
rect 5930 4313 5982 4319
rect 6044 4241 6072 4449
rect 6134 4371 6186 4377
rect 6134 4313 6186 4319
rect 6248 4241 6276 4449
rect 6338 4371 6390 4377
rect 6338 4313 6390 4319
rect 6452 4241 6480 4449
rect 6542 4371 6594 4377
rect 6542 4313 6594 4319
rect 6656 4241 6684 4449
rect 6746 4371 6798 4377
rect 6746 4313 6798 4319
rect 6860 4241 6888 4449
rect 6950 4371 7002 4377
rect 6950 4313 7002 4319
rect 7064 4241 7092 4449
rect 7154 4371 7206 4377
rect 7154 4313 7206 4319
rect 7268 4241 7296 4449
rect 7358 4371 7410 4377
rect 7358 4313 7410 4319
rect 7472 4241 7500 4449
rect 7562 4371 7614 4377
rect 7562 4313 7614 4319
rect 7676 4241 7704 4449
rect 7766 4371 7818 4377
rect 7766 4313 7818 4319
rect 7880 4241 7908 4449
rect 7970 4371 8022 4377
rect 7970 4313 8022 4319
rect 8084 4241 8112 4449
rect 8174 4371 8226 4377
rect 8174 4313 8226 4319
rect 8288 4241 8316 4449
rect 8378 4371 8430 4377
rect 8378 4313 8430 4319
rect 8492 4241 8520 4449
rect 8582 4371 8634 4377
rect 8582 4313 8634 4319
rect 8696 4241 8724 4449
rect 8786 4371 8838 4377
rect 8786 4313 8838 4319
rect 8900 4241 8928 4449
rect 8990 4371 9042 4377
rect 8990 4313 9042 4319
rect 9104 4241 9132 4449
rect 9194 4371 9246 4377
rect 9194 4313 9246 4319
rect 9308 4241 9336 4449
rect 9398 4371 9450 4377
rect 9398 4313 9450 4319
rect 9512 4241 9540 4449
rect 9602 4371 9654 4377
rect 9602 4313 9654 4319
rect 9716 4241 9744 4449
rect 9806 4371 9858 4377
rect 9806 4313 9858 4319
rect 9920 4241 9948 4449
rect 10010 4371 10062 4377
rect 10010 4313 10062 4319
rect 10124 4241 10152 4449
rect 10214 4371 10266 4377
rect 10214 4313 10266 4319
rect 10328 4241 10356 4449
rect 10418 4371 10470 4377
rect 10418 4313 10470 4319
rect 10532 4241 10560 4449
rect 10622 4371 10674 4377
rect 10622 4313 10674 4319
rect 10736 4241 10764 4449
rect 10826 4371 10878 4377
rect 10826 4313 10878 4319
rect 10940 4241 10968 4449
rect 11030 4371 11082 4377
rect 11030 4313 11082 4319
rect 11144 4241 11172 4449
rect 11234 4371 11286 4377
rect 11234 4313 11286 4319
rect 11348 4241 11376 4449
rect 11438 4371 11490 4377
rect 11438 4313 11490 4319
rect 11552 4241 11580 4449
rect 11642 4371 11694 4377
rect 11642 4313 11694 4319
rect 11756 4241 11784 4449
rect 11846 4371 11898 4377
rect 11846 4313 11898 4319
rect 11960 4241 11988 4449
rect 12050 4371 12102 4377
rect 12050 4313 12102 4319
rect 12164 4241 12192 4449
rect 12254 4371 12306 4377
rect 12254 4313 12306 4319
rect 12368 4241 12396 4449
rect 12458 4371 12510 4377
rect 12458 4313 12510 4319
rect 12572 4241 12600 4449
rect 12662 4371 12714 4377
rect 12662 4313 12714 4319
rect 12776 4241 12804 4449
rect 12866 4371 12918 4377
rect 12866 4313 12918 4319
rect 12980 4241 13008 4449
rect 13084 4371 13136 4377
rect 13084 4313 13136 4319
rect 8 4217 59 4224
rect 1640 4217 1691 4224
rect 3272 4217 3323 4224
rect 4904 4217 4955 4224
rect 6536 4217 6587 4224
rect 8168 4217 8219 4224
rect 9800 4217 9851 4224
rect 11432 4217 11483 4224
rect 13064 4217 13115 4224
rect 1 4165 7 4217
rect 59 4165 65 4217
rect 1633 4165 1639 4217
rect 1691 4165 1697 4217
rect 3265 4165 3271 4217
rect 3323 4165 3329 4217
rect 4897 4165 4903 4217
rect 4955 4165 4961 4217
rect 6529 4165 6535 4217
rect 6587 4165 6593 4217
rect 8161 4165 8167 4217
rect 8219 4165 8225 4217
rect 9793 4165 9799 4217
rect 9851 4165 9857 4217
rect 11425 4165 11431 4217
rect 11483 4165 11489 4217
rect 13057 4165 13063 4217
rect 13115 4165 13121 4217
rect 8 4158 59 4165
rect 1640 4158 1691 4165
rect 3272 4158 3323 4165
rect 4904 4158 4955 4165
rect 6536 4158 6587 4165
rect 8168 4158 8219 4165
rect 9800 4158 9851 4165
rect 11432 4158 11483 4165
rect 13064 4158 13115 4165
rect 8 4013 59 4020
rect 1640 4013 1691 4020
rect 3272 4013 3323 4020
rect 4904 4013 4955 4020
rect 6536 4013 6587 4020
rect 8168 4013 8219 4020
rect 9800 4013 9851 4020
rect 11432 4013 11483 4020
rect 13064 4013 13115 4020
rect 1 3961 7 4013
rect 59 3961 65 4013
rect 1633 3961 1639 4013
rect 1691 3961 1697 4013
rect 3265 3961 3271 4013
rect 3323 3961 3329 4013
rect 4897 3961 4903 4013
rect 4955 3961 4961 4013
rect 6529 3961 6535 4013
rect 6587 3961 6593 4013
rect 8161 3961 8167 4013
rect 8219 3961 8225 4013
rect 9793 3961 9799 4013
rect 9851 3961 9857 4013
rect 11425 3961 11431 4013
rect 11483 3961 11489 4013
rect 13057 3961 13063 4013
rect 13115 3961 13121 4013
rect 8 3954 59 3961
rect 1640 3954 1691 3961
rect 3272 3954 3323 3961
rect 4904 3954 4955 3961
rect 6536 3954 6587 3961
rect 8168 3954 8219 3961
rect 9800 3954 9851 3961
rect 11432 3954 11483 3961
rect 13064 3954 13115 3961
rect 8 3809 59 3816
rect 1640 3809 1691 3816
rect 3272 3809 3323 3816
rect 4904 3809 4955 3816
rect 6536 3809 6587 3816
rect 8168 3809 8219 3816
rect 9800 3809 9851 3816
rect 11432 3809 11483 3816
rect 13064 3809 13115 3816
rect 1 3757 7 3809
rect 59 3757 65 3809
rect 1633 3757 1639 3809
rect 1691 3757 1697 3809
rect 3265 3757 3271 3809
rect 3323 3757 3329 3809
rect 4897 3757 4903 3809
rect 4955 3757 4961 3809
rect 6529 3757 6535 3809
rect 6587 3757 6593 3809
rect 8161 3757 8167 3809
rect 8219 3757 8225 3809
rect 9793 3757 9799 3809
rect 9851 3757 9857 3809
rect 11425 3757 11431 3809
rect 11483 3757 11489 3809
rect 13057 3757 13063 3809
rect 13115 3757 13121 3809
rect 8 3750 59 3757
rect 1640 3750 1691 3757
rect 3272 3750 3323 3757
rect 4904 3750 4955 3757
rect 6536 3750 6587 3757
rect 8168 3750 8219 3757
rect 9800 3750 9851 3757
rect 11432 3750 11483 3757
rect 13064 3750 13115 3757
rect 8 3605 59 3612
rect 1640 3605 1691 3612
rect 3272 3605 3323 3612
rect 4904 3605 4955 3612
rect 6536 3605 6587 3612
rect 8168 3605 8219 3612
rect 9800 3605 9851 3612
rect 11432 3605 11483 3612
rect 13064 3605 13115 3612
rect 1 3553 7 3605
rect 59 3553 65 3605
rect 1633 3553 1639 3605
rect 1691 3553 1697 3605
rect 3265 3553 3271 3605
rect 3323 3553 3329 3605
rect 4897 3553 4903 3605
rect 4955 3553 4961 3605
rect 6529 3553 6535 3605
rect 6587 3553 6593 3605
rect 8161 3553 8167 3605
rect 8219 3553 8225 3605
rect 9793 3553 9799 3605
rect 9851 3553 9857 3605
rect 11425 3553 11431 3605
rect 11483 3553 11489 3605
rect 13057 3553 13063 3605
rect 13115 3553 13121 3605
rect 8 3546 59 3553
rect 1640 3546 1691 3553
rect 3272 3546 3323 3553
rect 4904 3546 4955 3553
rect 6536 3546 6587 3553
rect 8168 3546 8219 3553
rect 9800 3546 9851 3553
rect 11432 3546 11483 3553
rect 13064 3546 13115 3553
rect 8 3401 59 3408
rect 1640 3401 1691 3408
rect 3272 3401 3323 3408
rect 4904 3401 4955 3408
rect 6536 3401 6587 3408
rect 8168 3401 8219 3408
rect 9800 3401 9851 3408
rect 11432 3401 11483 3408
rect 13064 3401 13115 3408
rect 1 3349 7 3401
rect 59 3349 65 3401
rect 1633 3349 1639 3401
rect 1691 3349 1697 3401
rect 3265 3349 3271 3401
rect 3323 3349 3329 3401
rect 4897 3349 4903 3401
rect 4955 3349 4961 3401
rect 6529 3349 6535 3401
rect 6587 3349 6593 3401
rect 8161 3349 8167 3401
rect 8219 3349 8225 3401
rect 9793 3349 9799 3401
rect 9851 3349 9857 3401
rect 11425 3349 11431 3401
rect 11483 3349 11489 3401
rect 13057 3349 13063 3401
rect 13115 3349 13121 3401
rect 8 3342 59 3349
rect 1640 3342 1691 3349
rect 3272 3342 3323 3349
rect 4904 3342 4955 3349
rect 6536 3342 6587 3349
rect 8168 3342 8219 3349
rect 9800 3342 9851 3349
rect 11432 3342 11483 3349
rect 13064 3342 13115 3349
rect 8 3197 59 3204
rect 1640 3197 1691 3204
rect 3272 3197 3323 3204
rect 4904 3197 4955 3204
rect 6536 3197 6587 3204
rect 8168 3197 8219 3204
rect 9800 3197 9851 3204
rect 11432 3197 11483 3204
rect 13064 3197 13115 3204
rect 1 3145 7 3197
rect 59 3145 65 3197
rect 1633 3145 1639 3197
rect 1691 3145 1697 3197
rect 3265 3145 3271 3197
rect 3323 3145 3329 3197
rect 4897 3145 4903 3197
rect 4955 3145 4961 3197
rect 6529 3145 6535 3197
rect 6587 3145 6593 3197
rect 8161 3145 8167 3197
rect 8219 3145 8225 3197
rect 9793 3145 9799 3197
rect 9851 3145 9857 3197
rect 11425 3145 11431 3197
rect 11483 3145 11489 3197
rect 13057 3145 13063 3197
rect 13115 3145 13121 3197
rect 8 3138 59 3145
rect 1640 3138 1691 3145
rect 3272 3138 3323 3145
rect 4904 3138 4955 3145
rect 6536 3138 6587 3145
rect 8168 3138 8219 3145
rect 9800 3138 9851 3145
rect 11432 3138 11483 3145
rect 13064 3138 13115 3145
rect 8 2993 59 3000
rect 1640 2993 1691 3000
rect 3272 2993 3323 3000
rect 4904 2993 4955 3000
rect 6536 2993 6587 3000
rect 8168 2993 8219 3000
rect 9800 2993 9851 3000
rect 11432 2993 11483 3000
rect 13064 2993 13115 3000
rect 1 2941 7 2993
rect 59 2941 65 2993
rect 1633 2941 1639 2993
rect 1691 2941 1697 2993
rect 3265 2941 3271 2993
rect 3323 2941 3329 2993
rect 4897 2941 4903 2993
rect 4955 2941 4961 2993
rect 6529 2941 6535 2993
rect 6587 2941 6593 2993
rect 8161 2941 8167 2993
rect 8219 2941 8225 2993
rect 9793 2941 9799 2993
rect 9851 2941 9857 2993
rect 11425 2941 11431 2993
rect 11483 2941 11489 2993
rect 13057 2941 13063 2993
rect 13115 2941 13121 2993
rect 8 2934 59 2941
rect 1640 2934 1691 2941
rect 3272 2934 3323 2941
rect 4904 2934 4955 2941
rect 6536 2934 6587 2941
rect 8168 2934 8219 2941
rect 9800 2934 9851 2941
rect 11432 2934 11483 2941
rect 13064 2934 13115 2941
rect 8 2789 59 2796
rect 1640 2789 1691 2796
rect 3272 2789 3323 2796
rect 4904 2789 4955 2796
rect 6536 2789 6587 2796
rect 8168 2789 8219 2796
rect 9800 2789 9851 2796
rect 11432 2789 11483 2796
rect 13064 2789 13115 2796
rect 1 2737 7 2789
rect 59 2737 65 2789
rect 1633 2737 1639 2789
rect 1691 2737 1697 2789
rect 3265 2737 3271 2789
rect 3323 2737 3329 2789
rect 4897 2737 4903 2789
rect 4955 2737 4961 2789
rect 6529 2737 6535 2789
rect 6587 2737 6593 2789
rect 8161 2737 8167 2789
rect 8219 2737 8225 2789
rect 9793 2737 9799 2789
rect 9851 2737 9857 2789
rect 11425 2737 11431 2789
rect 11483 2737 11489 2789
rect 13057 2737 13063 2789
rect 13115 2737 13121 2789
rect 8 2730 59 2737
rect 1640 2730 1691 2737
rect 3272 2730 3323 2737
rect 4904 2730 4955 2737
rect 6536 2730 6587 2737
rect 8168 2730 8219 2737
rect 9800 2730 9851 2737
rect 11432 2730 11483 2737
rect 13064 2730 13115 2737
rect 128 2505 156 2713
rect 218 2635 270 2641
rect 218 2577 270 2583
rect 332 2505 360 2713
rect 422 2635 474 2641
rect 422 2577 474 2583
rect 536 2505 564 2713
rect 626 2635 678 2641
rect 626 2577 678 2583
rect 740 2505 768 2713
rect 830 2635 882 2641
rect 830 2577 882 2583
rect 944 2505 972 2713
rect 1034 2635 1086 2641
rect 1034 2577 1086 2583
rect 1148 2505 1176 2713
rect 1238 2635 1290 2641
rect 1238 2577 1290 2583
rect 1352 2505 1380 2713
rect 1442 2635 1494 2641
rect 1442 2577 1494 2583
rect 1556 2505 1584 2713
rect 1646 2635 1698 2641
rect 1646 2577 1698 2583
rect 1760 2505 1788 2713
rect 1850 2635 1902 2641
rect 1850 2577 1902 2583
rect 1964 2505 1992 2713
rect 2054 2635 2106 2641
rect 2054 2577 2106 2583
rect 2168 2505 2196 2713
rect 2258 2635 2310 2641
rect 2258 2577 2310 2583
rect 2372 2505 2400 2713
rect 2462 2635 2514 2641
rect 2462 2577 2514 2583
rect 2576 2505 2604 2713
rect 2666 2635 2718 2641
rect 2666 2577 2718 2583
rect 2780 2505 2808 2713
rect 2870 2635 2922 2641
rect 2870 2577 2922 2583
rect 2984 2505 3012 2713
rect 3074 2635 3126 2641
rect 3074 2577 3126 2583
rect 3188 2505 3216 2713
rect 3278 2635 3330 2641
rect 3278 2577 3330 2583
rect 3392 2505 3420 2713
rect 3482 2635 3534 2641
rect 3482 2577 3534 2583
rect 3596 2505 3624 2713
rect 3686 2635 3738 2641
rect 3686 2577 3738 2583
rect 3800 2505 3828 2713
rect 3890 2635 3942 2641
rect 3890 2577 3942 2583
rect 4004 2505 4032 2713
rect 4094 2635 4146 2641
rect 4094 2577 4146 2583
rect 4208 2505 4236 2713
rect 4298 2635 4350 2641
rect 4298 2577 4350 2583
rect 4412 2505 4440 2713
rect 4502 2635 4554 2641
rect 4502 2577 4554 2583
rect 4616 2505 4644 2713
rect 4706 2635 4758 2641
rect 4706 2577 4758 2583
rect 4820 2505 4848 2713
rect 4910 2635 4962 2641
rect 4910 2577 4962 2583
rect 5024 2505 5052 2713
rect 5114 2635 5166 2641
rect 5114 2577 5166 2583
rect 5228 2505 5256 2713
rect 5318 2635 5370 2641
rect 5318 2577 5370 2583
rect 5432 2505 5460 2713
rect 5522 2635 5574 2641
rect 5522 2577 5574 2583
rect 5636 2505 5664 2713
rect 5726 2635 5778 2641
rect 5726 2577 5778 2583
rect 5840 2505 5868 2713
rect 5930 2635 5982 2641
rect 5930 2577 5982 2583
rect 6044 2505 6072 2713
rect 6134 2635 6186 2641
rect 6134 2577 6186 2583
rect 6248 2505 6276 2713
rect 6338 2635 6390 2641
rect 6338 2577 6390 2583
rect 6452 2505 6480 2713
rect 6542 2635 6594 2641
rect 6542 2577 6594 2583
rect 6656 2505 6684 2713
rect 6746 2635 6798 2641
rect 6746 2577 6798 2583
rect 6860 2505 6888 2713
rect 6950 2635 7002 2641
rect 6950 2577 7002 2583
rect 7064 2505 7092 2713
rect 7154 2635 7206 2641
rect 7154 2577 7206 2583
rect 7268 2505 7296 2713
rect 7358 2635 7410 2641
rect 7358 2577 7410 2583
rect 7472 2505 7500 2713
rect 7562 2635 7614 2641
rect 7562 2577 7614 2583
rect 7676 2505 7704 2713
rect 7766 2635 7818 2641
rect 7766 2577 7818 2583
rect 7880 2505 7908 2713
rect 7970 2635 8022 2641
rect 7970 2577 8022 2583
rect 8084 2505 8112 2713
rect 8174 2635 8226 2641
rect 8174 2577 8226 2583
rect 8288 2505 8316 2713
rect 8378 2635 8430 2641
rect 8378 2577 8430 2583
rect 8492 2505 8520 2713
rect 8582 2635 8634 2641
rect 8582 2577 8634 2583
rect 8696 2505 8724 2713
rect 8786 2635 8838 2641
rect 8786 2577 8838 2583
rect 8900 2505 8928 2713
rect 8990 2635 9042 2641
rect 8990 2577 9042 2583
rect 9104 2505 9132 2713
rect 9194 2635 9246 2641
rect 9194 2577 9246 2583
rect 9308 2505 9336 2713
rect 9398 2635 9450 2641
rect 9398 2577 9450 2583
rect 9512 2505 9540 2713
rect 9602 2635 9654 2641
rect 9602 2577 9654 2583
rect 9716 2505 9744 2713
rect 9806 2635 9858 2641
rect 9806 2577 9858 2583
rect 9920 2505 9948 2713
rect 10010 2635 10062 2641
rect 10010 2577 10062 2583
rect 10124 2505 10152 2713
rect 10214 2635 10266 2641
rect 10214 2577 10266 2583
rect 10328 2505 10356 2713
rect 10418 2635 10470 2641
rect 10418 2577 10470 2583
rect 10532 2505 10560 2713
rect 10622 2635 10674 2641
rect 10622 2577 10674 2583
rect 10736 2505 10764 2713
rect 10826 2635 10878 2641
rect 10826 2577 10878 2583
rect 10940 2505 10968 2713
rect 11030 2635 11082 2641
rect 11030 2577 11082 2583
rect 11144 2505 11172 2713
rect 11234 2635 11286 2641
rect 11234 2577 11286 2583
rect 11348 2505 11376 2713
rect 11438 2635 11490 2641
rect 11438 2577 11490 2583
rect 11552 2505 11580 2713
rect 11642 2635 11694 2641
rect 11642 2577 11694 2583
rect 11756 2505 11784 2713
rect 11846 2635 11898 2641
rect 11846 2577 11898 2583
rect 11960 2505 11988 2713
rect 12050 2635 12102 2641
rect 12050 2577 12102 2583
rect 12164 2505 12192 2713
rect 12254 2635 12306 2641
rect 12254 2577 12306 2583
rect 12368 2505 12396 2713
rect 12458 2635 12510 2641
rect 12458 2577 12510 2583
rect 12572 2505 12600 2713
rect 12662 2635 12714 2641
rect 12662 2577 12714 2583
rect 12776 2505 12804 2713
rect 12866 2635 12918 2641
rect 12866 2577 12918 2583
rect 12980 2505 13008 2713
rect 13084 2635 13136 2641
rect 13084 2577 13136 2583
rect 8 2481 59 2488
rect 1640 2481 1691 2488
rect 3272 2481 3323 2488
rect 4904 2481 4955 2488
rect 6536 2481 6587 2488
rect 8168 2481 8219 2488
rect 9800 2481 9851 2488
rect 11432 2481 11483 2488
rect 13064 2481 13115 2488
rect 1 2429 7 2481
rect 59 2429 65 2481
rect 1633 2429 1639 2481
rect 1691 2429 1697 2481
rect 3265 2429 3271 2481
rect 3323 2429 3329 2481
rect 4897 2429 4903 2481
rect 4955 2429 4961 2481
rect 6529 2429 6535 2481
rect 6587 2429 6593 2481
rect 8161 2429 8167 2481
rect 8219 2429 8225 2481
rect 9793 2429 9799 2481
rect 9851 2429 9857 2481
rect 11425 2429 11431 2481
rect 11483 2429 11489 2481
rect 13057 2429 13063 2481
rect 13115 2429 13121 2481
rect 8 2422 59 2429
rect 1640 2422 1691 2429
rect 3272 2422 3323 2429
rect 4904 2422 4955 2429
rect 6536 2422 6587 2429
rect 8168 2422 8219 2429
rect 9800 2422 9851 2429
rect 11432 2422 11483 2429
rect 13064 2422 13115 2429
rect 8 2277 59 2284
rect 1640 2277 1691 2284
rect 3272 2277 3323 2284
rect 4904 2277 4955 2284
rect 6536 2277 6587 2284
rect 8168 2277 8219 2284
rect 9800 2277 9851 2284
rect 11432 2277 11483 2284
rect 13064 2277 13115 2284
rect 1 2225 7 2277
rect 59 2225 65 2277
rect 1633 2225 1639 2277
rect 1691 2225 1697 2277
rect 3265 2225 3271 2277
rect 3323 2225 3329 2277
rect 4897 2225 4903 2277
rect 4955 2225 4961 2277
rect 6529 2225 6535 2277
rect 6587 2225 6593 2277
rect 8161 2225 8167 2277
rect 8219 2225 8225 2277
rect 9793 2225 9799 2277
rect 9851 2225 9857 2277
rect 11425 2225 11431 2277
rect 11483 2225 11489 2277
rect 13057 2225 13063 2277
rect 13115 2225 13121 2277
rect 8 2218 59 2225
rect 1640 2218 1691 2225
rect 3272 2218 3323 2225
rect 4904 2218 4955 2225
rect 6536 2218 6587 2225
rect 8168 2218 8219 2225
rect 9800 2218 9851 2225
rect 11432 2218 11483 2225
rect 13064 2218 13115 2225
rect 8 2073 59 2080
rect 1640 2073 1691 2080
rect 3272 2073 3323 2080
rect 4904 2073 4955 2080
rect 6536 2073 6587 2080
rect 8168 2073 8219 2080
rect 9800 2073 9851 2080
rect 11432 2073 11483 2080
rect 13064 2073 13115 2080
rect 1 2021 7 2073
rect 59 2021 65 2073
rect 1633 2021 1639 2073
rect 1691 2021 1697 2073
rect 3265 2021 3271 2073
rect 3323 2021 3329 2073
rect 4897 2021 4903 2073
rect 4955 2021 4961 2073
rect 6529 2021 6535 2073
rect 6587 2021 6593 2073
rect 8161 2021 8167 2073
rect 8219 2021 8225 2073
rect 9793 2021 9799 2073
rect 9851 2021 9857 2073
rect 11425 2021 11431 2073
rect 11483 2021 11489 2073
rect 13057 2021 13063 2073
rect 13115 2021 13121 2073
rect 8 2014 59 2021
rect 1640 2014 1691 2021
rect 3272 2014 3323 2021
rect 4904 2014 4955 2021
rect 6536 2014 6587 2021
rect 8168 2014 8219 2021
rect 9800 2014 9851 2021
rect 11432 2014 11483 2021
rect 13064 2014 13115 2021
rect 8 1869 59 1876
rect 1640 1869 1691 1876
rect 3272 1869 3323 1876
rect 4904 1869 4955 1876
rect 6536 1869 6587 1876
rect 8168 1869 8219 1876
rect 9800 1869 9851 1876
rect 11432 1869 11483 1876
rect 13064 1869 13115 1876
rect 1 1817 7 1869
rect 59 1817 65 1869
rect 1633 1817 1639 1869
rect 1691 1817 1697 1869
rect 3265 1817 3271 1869
rect 3323 1817 3329 1869
rect 4897 1817 4903 1869
rect 4955 1817 4961 1869
rect 6529 1817 6535 1869
rect 6587 1817 6593 1869
rect 8161 1817 8167 1869
rect 8219 1817 8225 1869
rect 9793 1817 9799 1869
rect 9851 1817 9857 1869
rect 11425 1817 11431 1869
rect 11483 1817 11489 1869
rect 13057 1817 13063 1869
rect 13115 1817 13121 1869
rect 8 1810 59 1817
rect 1640 1810 1691 1817
rect 3272 1810 3323 1817
rect 4904 1810 4955 1817
rect 6536 1810 6587 1817
rect 8168 1810 8219 1817
rect 9800 1810 9851 1817
rect 11432 1810 11483 1817
rect 13064 1810 13115 1817
rect 8 1665 59 1672
rect 1640 1665 1691 1672
rect 3272 1665 3323 1672
rect 4904 1665 4955 1672
rect 6536 1665 6587 1672
rect 8168 1665 8219 1672
rect 9800 1665 9851 1672
rect 11432 1665 11483 1672
rect 13064 1665 13115 1672
rect 1 1613 7 1665
rect 59 1613 65 1665
rect 1633 1613 1639 1665
rect 1691 1613 1697 1665
rect 3265 1613 3271 1665
rect 3323 1613 3329 1665
rect 4897 1613 4903 1665
rect 4955 1613 4961 1665
rect 6529 1613 6535 1665
rect 6587 1613 6593 1665
rect 8161 1613 8167 1665
rect 8219 1613 8225 1665
rect 9793 1613 9799 1665
rect 9851 1613 9857 1665
rect 11425 1613 11431 1665
rect 11483 1613 11489 1665
rect 13057 1613 13063 1665
rect 13115 1613 13121 1665
rect 8 1606 59 1613
rect 1640 1606 1691 1613
rect 3272 1606 3323 1613
rect 4904 1606 4955 1613
rect 6536 1606 6587 1613
rect 8168 1606 8219 1613
rect 9800 1606 9851 1613
rect 11432 1606 11483 1613
rect 13064 1606 13115 1613
rect 8 1461 59 1468
rect 1640 1461 1691 1468
rect 3272 1461 3323 1468
rect 4904 1461 4955 1468
rect 6536 1461 6587 1468
rect 8168 1461 8219 1468
rect 9800 1461 9851 1468
rect 11432 1461 11483 1468
rect 13064 1461 13115 1468
rect 1 1409 7 1461
rect 59 1409 65 1461
rect 1633 1409 1639 1461
rect 1691 1409 1697 1461
rect 3265 1409 3271 1461
rect 3323 1409 3329 1461
rect 4897 1409 4903 1461
rect 4955 1409 4961 1461
rect 6529 1409 6535 1461
rect 6587 1409 6593 1461
rect 8161 1409 8167 1461
rect 8219 1409 8225 1461
rect 9793 1409 9799 1461
rect 9851 1409 9857 1461
rect 11425 1409 11431 1461
rect 11483 1409 11489 1461
rect 13057 1409 13063 1461
rect 13115 1409 13121 1461
rect 8 1402 59 1409
rect 1640 1402 1691 1409
rect 3272 1402 3323 1409
rect 4904 1402 4955 1409
rect 6536 1402 6587 1409
rect 8168 1402 8219 1409
rect 9800 1402 9851 1409
rect 11432 1402 11483 1409
rect 13064 1402 13115 1409
rect 8 1257 59 1264
rect 1640 1257 1691 1264
rect 3272 1257 3323 1264
rect 4904 1257 4955 1264
rect 6536 1257 6587 1264
rect 8168 1257 8219 1264
rect 9800 1257 9851 1264
rect 11432 1257 11483 1264
rect 13064 1257 13115 1264
rect 1 1205 7 1257
rect 59 1205 65 1257
rect 1633 1205 1639 1257
rect 1691 1205 1697 1257
rect 3265 1205 3271 1257
rect 3323 1205 3329 1257
rect 4897 1205 4903 1257
rect 4955 1205 4961 1257
rect 6529 1205 6535 1257
rect 6587 1205 6593 1257
rect 8161 1205 8167 1257
rect 8219 1205 8225 1257
rect 9793 1205 9799 1257
rect 9851 1205 9857 1257
rect 11425 1205 11431 1257
rect 11483 1205 11489 1257
rect 13057 1205 13063 1257
rect 13115 1205 13121 1257
rect 8 1198 59 1205
rect 1640 1198 1691 1205
rect 3272 1198 3323 1205
rect 4904 1198 4955 1205
rect 6536 1198 6587 1205
rect 8168 1198 8219 1205
rect 9800 1198 9851 1205
rect 11432 1198 11483 1205
rect 13064 1198 13115 1205
rect 8 1053 59 1060
rect 1640 1053 1691 1060
rect 3272 1053 3323 1060
rect 4904 1053 4955 1060
rect 6536 1053 6587 1060
rect 8168 1053 8219 1060
rect 9800 1053 9851 1060
rect 11432 1053 11483 1060
rect 13064 1053 13115 1060
rect 1 1001 7 1053
rect 59 1001 65 1053
rect 1633 1001 1639 1053
rect 1691 1001 1697 1053
rect 3265 1001 3271 1053
rect 3323 1001 3329 1053
rect 4897 1001 4903 1053
rect 4955 1001 4961 1053
rect 6529 1001 6535 1053
rect 6587 1001 6593 1053
rect 8161 1001 8167 1053
rect 8219 1001 8225 1053
rect 9793 1001 9799 1053
rect 9851 1001 9857 1053
rect 11425 1001 11431 1053
rect 11483 1001 11489 1053
rect 13057 1001 13063 1053
rect 13115 1001 13121 1053
rect 8 994 59 1001
rect 1640 994 1691 1001
rect 3272 994 3323 1001
rect 4904 994 4955 1001
rect 6536 994 6587 1001
rect 8168 994 8219 1001
rect 9800 994 9851 1001
rect 11432 994 11483 1001
rect 13064 994 13115 1001
rect 128 -14 156 977
rect 218 899 270 905
rect 218 841 270 847
rect 332 -14 360 977
rect 422 899 474 905
rect 422 841 474 847
rect 536 -14 564 977
rect 626 899 678 905
rect 626 841 678 847
rect 740 -14 768 977
rect 830 899 882 905
rect 830 841 882 847
rect 944 -14 972 977
rect 1034 899 1086 905
rect 1034 841 1086 847
rect 1148 -14 1176 977
rect 1238 899 1290 905
rect 1238 841 1290 847
rect 1352 -14 1380 977
rect 1442 899 1494 905
rect 1442 841 1494 847
rect 1556 -14 1584 977
rect 1646 899 1698 905
rect 1646 841 1698 847
rect 1760 -14 1788 977
rect 1850 899 1902 905
rect 1850 841 1902 847
rect 1964 -14 1992 977
rect 2054 899 2106 905
rect 2054 841 2106 847
rect 2168 -14 2196 977
rect 2258 899 2310 905
rect 2258 841 2310 847
rect 2372 -14 2400 977
rect 2462 899 2514 905
rect 2462 841 2514 847
rect 2576 -14 2604 977
rect 2666 899 2718 905
rect 2666 841 2718 847
rect 2780 -14 2808 977
rect 2870 899 2922 905
rect 2870 841 2922 847
rect 2984 -14 3012 977
rect 3074 899 3126 905
rect 3074 841 3126 847
rect 3188 -14 3216 977
rect 3278 899 3330 905
rect 3278 841 3330 847
rect 3392 -14 3420 977
rect 3482 899 3534 905
rect 3482 841 3534 847
rect 3596 -14 3624 977
rect 3686 899 3738 905
rect 3686 841 3738 847
rect 3800 -14 3828 977
rect 3890 899 3942 905
rect 3890 841 3942 847
rect 4004 -14 4032 977
rect 4094 899 4146 905
rect 4094 841 4146 847
rect 4208 -14 4236 977
rect 4298 899 4350 905
rect 4298 841 4350 847
rect 4412 -14 4440 977
rect 4502 899 4554 905
rect 4502 841 4554 847
rect 4616 -14 4644 977
rect 4706 899 4758 905
rect 4706 841 4758 847
rect 4820 -14 4848 977
rect 4910 899 4962 905
rect 4910 841 4962 847
rect 5024 -14 5052 977
rect 5114 899 5166 905
rect 5114 841 5166 847
rect 5228 -14 5256 977
rect 5318 899 5370 905
rect 5318 841 5370 847
rect 5432 -14 5460 977
rect 5522 899 5574 905
rect 5522 841 5574 847
rect 5636 -14 5664 977
rect 5726 899 5778 905
rect 5726 841 5778 847
rect 5840 -14 5868 977
rect 5930 899 5982 905
rect 5930 841 5982 847
rect 6044 -14 6072 977
rect 6134 899 6186 905
rect 6134 841 6186 847
rect 6248 -14 6276 977
rect 6338 899 6390 905
rect 6338 841 6390 847
rect 6452 -14 6480 977
rect 6542 899 6594 905
rect 6542 841 6594 847
rect 6656 -14 6684 977
rect 6746 899 6798 905
rect 6746 841 6798 847
rect 6860 -14 6888 977
rect 6950 899 7002 905
rect 6950 841 7002 847
rect 7064 -14 7092 977
rect 7154 899 7206 905
rect 7154 841 7206 847
rect 7268 -14 7296 977
rect 7358 899 7410 905
rect 7358 841 7410 847
rect 7472 -14 7500 977
rect 7562 899 7614 905
rect 7562 841 7614 847
rect 7676 -14 7704 977
rect 7766 899 7818 905
rect 7766 841 7818 847
rect 7880 -14 7908 977
rect 7970 899 8022 905
rect 7970 841 8022 847
rect 8084 -14 8112 977
rect 8174 899 8226 905
rect 8174 841 8226 847
rect 8288 -14 8316 977
rect 8378 899 8430 905
rect 8378 841 8430 847
rect 8492 -14 8520 977
rect 8582 899 8634 905
rect 8582 841 8634 847
rect 8696 -14 8724 977
rect 8786 899 8838 905
rect 8786 841 8838 847
rect 8900 -14 8928 977
rect 8990 899 9042 905
rect 8990 841 9042 847
rect 9104 -14 9132 977
rect 9194 899 9246 905
rect 9194 841 9246 847
rect 9308 -14 9336 977
rect 9398 899 9450 905
rect 9398 841 9450 847
rect 9512 -14 9540 977
rect 9602 899 9654 905
rect 9602 841 9654 847
rect 9716 -14 9744 977
rect 9806 899 9858 905
rect 9806 841 9858 847
rect 9920 -14 9948 977
rect 10010 899 10062 905
rect 10010 841 10062 847
rect 10124 -14 10152 977
rect 10214 899 10266 905
rect 10214 841 10266 847
rect 10328 -14 10356 977
rect 10418 899 10470 905
rect 10418 841 10470 847
rect 10532 -14 10560 977
rect 10622 899 10674 905
rect 10622 841 10674 847
rect 10736 -14 10764 977
rect 10826 899 10878 905
rect 10826 841 10878 847
rect 10940 -14 10968 977
rect 11030 899 11082 905
rect 11030 841 11082 847
rect 11144 -14 11172 977
rect 11234 899 11286 905
rect 11234 841 11286 847
rect 11348 -14 11376 977
rect 11438 899 11490 905
rect 11438 841 11490 847
rect 11552 -14 11580 977
rect 11642 899 11694 905
rect 11642 841 11694 847
rect 11756 -14 11784 977
rect 11846 899 11898 905
rect 11846 841 11898 847
rect 11960 -14 11988 977
rect 12050 899 12102 905
rect 12050 841 12102 847
rect 12164 -14 12192 977
rect 12254 899 12306 905
rect 12254 841 12306 847
rect 12368 -14 12396 977
rect 12458 899 12510 905
rect 12458 841 12510 847
rect 12572 -14 12600 977
rect 12662 899 12714 905
rect 12662 841 12714 847
rect 12776 -14 12804 977
rect 12866 899 12918 905
rect 12866 841 12918 847
rect 12980 -14 13008 977
rect 13084 899 13136 905
rect 13084 841 13136 847
rect 13277 396 13305 7853
rect 13131 368 13305 396
<< via1 >>
rect 7 7884 59 7893
rect 7 7850 16 7884
rect 16 7850 50 7884
rect 50 7850 59 7884
rect 7 7841 59 7850
rect 1639 7884 1691 7893
rect 1639 7850 1648 7884
rect 1648 7850 1682 7884
rect 1682 7850 1691 7884
rect 1639 7841 1691 7850
rect 3271 7884 3323 7893
rect 3271 7850 3280 7884
rect 3280 7850 3314 7884
rect 3314 7850 3323 7884
rect 3271 7841 3323 7850
rect 4903 7884 4955 7893
rect 4903 7850 4912 7884
rect 4912 7850 4946 7884
rect 4946 7850 4955 7884
rect 4903 7841 4955 7850
rect 6535 7884 6587 7893
rect 6535 7850 6544 7884
rect 6544 7850 6578 7884
rect 6578 7850 6587 7884
rect 6535 7841 6587 7850
rect 8167 7884 8219 7893
rect 8167 7850 8176 7884
rect 8176 7850 8210 7884
rect 8210 7850 8219 7884
rect 8167 7841 8219 7850
rect 9799 7884 9851 7893
rect 9799 7850 9808 7884
rect 9808 7850 9842 7884
rect 9842 7850 9851 7884
rect 9799 7841 9851 7850
rect 11431 7884 11483 7893
rect 11431 7850 11440 7884
rect 11440 7850 11474 7884
rect 11474 7850 11483 7884
rect 11431 7841 11483 7850
rect 13063 7884 13115 7893
rect 13063 7850 13072 7884
rect 13072 7850 13106 7884
rect 13106 7850 13115 7884
rect 13063 7841 13115 7850
rect 7 7680 59 7689
rect 7 7646 16 7680
rect 16 7646 50 7680
rect 50 7646 59 7680
rect 7 7637 59 7646
rect 1639 7680 1691 7689
rect 1639 7646 1648 7680
rect 1648 7646 1682 7680
rect 1682 7646 1691 7680
rect 1639 7637 1691 7646
rect 3271 7680 3323 7689
rect 3271 7646 3280 7680
rect 3280 7646 3314 7680
rect 3314 7646 3323 7680
rect 3271 7637 3323 7646
rect 4903 7680 4955 7689
rect 4903 7646 4912 7680
rect 4912 7646 4946 7680
rect 4946 7646 4955 7680
rect 4903 7637 4955 7646
rect 6535 7680 6587 7689
rect 6535 7646 6544 7680
rect 6544 7646 6578 7680
rect 6578 7646 6587 7680
rect 6535 7637 6587 7646
rect 8167 7680 8219 7689
rect 8167 7646 8176 7680
rect 8176 7646 8210 7680
rect 8210 7646 8219 7680
rect 8167 7637 8219 7646
rect 9799 7680 9851 7689
rect 9799 7646 9808 7680
rect 9808 7646 9842 7680
rect 9842 7646 9851 7680
rect 9799 7637 9851 7646
rect 11431 7680 11483 7689
rect 11431 7646 11440 7680
rect 11440 7646 11474 7680
rect 11474 7646 11483 7680
rect 11431 7637 11483 7646
rect 13063 7680 13115 7689
rect 13063 7646 13072 7680
rect 13072 7646 13106 7680
rect 13106 7646 13115 7680
rect 13063 7637 13115 7646
rect 7 7476 59 7485
rect 7 7442 16 7476
rect 16 7442 50 7476
rect 50 7442 59 7476
rect 7 7433 59 7442
rect 1639 7476 1691 7485
rect 1639 7442 1648 7476
rect 1648 7442 1682 7476
rect 1682 7442 1691 7476
rect 1639 7433 1691 7442
rect 3271 7476 3323 7485
rect 3271 7442 3280 7476
rect 3280 7442 3314 7476
rect 3314 7442 3323 7476
rect 3271 7433 3323 7442
rect 4903 7476 4955 7485
rect 4903 7442 4912 7476
rect 4912 7442 4946 7476
rect 4946 7442 4955 7476
rect 4903 7433 4955 7442
rect 6535 7476 6587 7485
rect 6535 7442 6544 7476
rect 6544 7442 6578 7476
rect 6578 7442 6587 7476
rect 6535 7433 6587 7442
rect 8167 7476 8219 7485
rect 8167 7442 8176 7476
rect 8176 7442 8210 7476
rect 8210 7442 8219 7476
rect 8167 7433 8219 7442
rect 9799 7476 9851 7485
rect 9799 7442 9808 7476
rect 9808 7442 9842 7476
rect 9842 7442 9851 7476
rect 9799 7433 9851 7442
rect 11431 7476 11483 7485
rect 11431 7442 11440 7476
rect 11440 7442 11474 7476
rect 11474 7442 11483 7476
rect 11431 7433 11483 7442
rect 13063 7476 13115 7485
rect 13063 7442 13072 7476
rect 13072 7442 13106 7476
rect 13106 7442 13115 7476
rect 13063 7433 13115 7442
rect 7 7272 59 7281
rect 7 7238 16 7272
rect 16 7238 50 7272
rect 50 7238 59 7272
rect 7 7229 59 7238
rect 1639 7272 1691 7281
rect 1639 7238 1648 7272
rect 1648 7238 1682 7272
rect 1682 7238 1691 7272
rect 1639 7229 1691 7238
rect 3271 7272 3323 7281
rect 3271 7238 3280 7272
rect 3280 7238 3314 7272
rect 3314 7238 3323 7272
rect 3271 7229 3323 7238
rect 4903 7272 4955 7281
rect 4903 7238 4912 7272
rect 4912 7238 4946 7272
rect 4946 7238 4955 7272
rect 4903 7229 4955 7238
rect 6535 7272 6587 7281
rect 6535 7238 6544 7272
rect 6544 7238 6578 7272
rect 6578 7238 6587 7272
rect 6535 7229 6587 7238
rect 8167 7272 8219 7281
rect 8167 7238 8176 7272
rect 8176 7238 8210 7272
rect 8210 7238 8219 7272
rect 8167 7229 8219 7238
rect 9799 7272 9851 7281
rect 9799 7238 9808 7272
rect 9808 7238 9842 7272
rect 9842 7238 9851 7272
rect 9799 7229 9851 7238
rect 11431 7272 11483 7281
rect 11431 7238 11440 7272
rect 11440 7238 11474 7272
rect 11474 7238 11483 7272
rect 11431 7229 11483 7238
rect 13063 7272 13115 7281
rect 13063 7238 13072 7272
rect 13072 7238 13106 7272
rect 13106 7238 13115 7272
rect 13063 7229 13115 7238
rect 7 7068 59 7077
rect 7 7034 16 7068
rect 16 7034 50 7068
rect 50 7034 59 7068
rect 7 7025 59 7034
rect 1639 7068 1691 7077
rect 1639 7034 1648 7068
rect 1648 7034 1682 7068
rect 1682 7034 1691 7068
rect 1639 7025 1691 7034
rect 3271 7068 3323 7077
rect 3271 7034 3280 7068
rect 3280 7034 3314 7068
rect 3314 7034 3323 7068
rect 3271 7025 3323 7034
rect 4903 7068 4955 7077
rect 4903 7034 4912 7068
rect 4912 7034 4946 7068
rect 4946 7034 4955 7068
rect 4903 7025 4955 7034
rect 6535 7068 6587 7077
rect 6535 7034 6544 7068
rect 6544 7034 6578 7068
rect 6578 7034 6587 7068
rect 6535 7025 6587 7034
rect 8167 7068 8219 7077
rect 8167 7034 8176 7068
rect 8176 7034 8210 7068
rect 8210 7034 8219 7068
rect 8167 7025 8219 7034
rect 9799 7068 9851 7077
rect 9799 7034 9808 7068
rect 9808 7034 9842 7068
rect 9842 7034 9851 7068
rect 9799 7025 9851 7034
rect 11431 7068 11483 7077
rect 11431 7034 11440 7068
rect 11440 7034 11474 7068
rect 11474 7034 11483 7068
rect 11431 7025 11483 7034
rect 13063 7068 13115 7077
rect 13063 7034 13072 7068
rect 13072 7034 13106 7068
rect 13106 7034 13115 7068
rect 13063 7025 13115 7034
rect 7 6864 59 6873
rect 7 6830 16 6864
rect 16 6830 50 6864
rect 50 6830 59 6864
rect 7 6821 59 6830
rect 1639 6864 1691 6873
rect 1639 6830 1648 6864
rect 1648 6830 1682 6864
rect 1682 6830 1691 6864
rect 1639 6821 1691 6830
rect 3271 6864 3323 6873
rect 3271 6830 3280 6864
rect 3280 6830 3314 6864
rect 3314 6830 3323 6864
rect 3271 6821 3323 6830
rect 4903 6864 4955 6873
rect 4903 6830 4912 6864
rect 4912 6830 4946 6864
rect 4946 6830 4955 6864
rect 4903 6821 4955 6830
rect 6535 6864 6587 6873
rect 6535 6830 6544 6864
rect 6544 6830 6578 6864
rect 6578 6830 6587 6864
rect 6535 6821 6587 6830
rect 8167 6864 8219 6873
rect 8167 6830 8176 6864
rect 8176 6830 8210 6864
rect 8210 6830 8219 6864
rect 8167 6821 8219 6830
rect 9799 6864 9851 6873
rect 9799 6830 9808 6864
rect 9808 6830 9842 6864
rect 9842 6830 9851 6864
rect 9799 6821 9851 6830
rect 11431 6864 11483 6873
rect 11431 6830 11440 6864
rect 11440 6830 11474 6864
rect 11474 6830 11483 6864
rect 11431 6821 11483 6830
rect 13063 6864 13115 6873
rect 13063 6830 13072 6864
rect 13072 6830 13106 6864
rect 13106 6830 13115 6864
rect 13063 6821 13115 6830
rect 7 6660 59 6669
rect 7 6626 16 6660
rect 16 6626 50 6660
rect 50 6626 59 6660
rect 7 6617 59 6626
rect 1639 6660 1691 6669
rect 1639 6626 1648 6660
rect 1648 6626 1682 6660
rect 1682 6626 1691 6660
rect 1639 6617 1691 6626
rect 3271 6660 3323 6669
rect 3271 6626 3280 6660
rect 3280 6626 3314 6660
rect 3314 6626 3323 6660
rect 3271 6617 3323 6626
rect 4903 6660 4955 6669
rect 4903 6626 4912 6660
rect 4912 6626 4946 6660
rect 4946 6626 4955 6660
rect 4903 6617 4955 6626
rect 6535 6660 6587 6669
rect 6535 6626 6544 6660
rect 6544 6626 6578 6660
rect 6578 6626 6587 6660
rect 6535 6617 6587 6626
rect 8167 6660 8219 6669
rect 8167 6626 8176 6660
rect 8176 6626 8210 6660
rect 8210 6626 8219 6660
rect 8167 6617 8219 6626
rect 9799 6660 9851 6669
rect 9799 6626 9808 6660
rect 9808 6626 9842 6660
rect 9842 6626 9851 6660
rect 9799 6617 9851 6626
rect 11431 6660 11483 6669
rect 11431 6626 11440 6660
rect 11440 6626 11474 6660
rect 11474 6626 11483 6660
rect 11431 6617 11483 6626
rect 13063 6660 13115 6669
rect 13063 6626 13072 6660
rect 13072 6626 13106 6660
rect 13106 6626 13115 6660
rect 13063 6617 13115 6626
rect 7 6456 59 6465
rect 7 6422 16 6456
rect 16 6422 50 6456
rect 50 6422 59 6456
rect 7 6413 59 6422
rect 1639 6456 1691 6465
rect 1639 6422 1648 6456
rect 1648 6422 1682 6456
rect 1682 6422 1691 6456
rect 1639 6413 1691 6422
rect 3271 6456 3323 6465
rect 3271 6422 3280 6456
rect 3280 6422 3314 6456
rect 3314 6422 3323 6456
rect 3271 6413 3323 6422
rect 4903 6456 4955 6465
rect 4903 6422 4912 6456
rect 4912 6422 4946 6456
rect 4946 6422 4955 6456
rect 4903 6413 4955 6422
rect 6535 6456 6587 6465
rect 6535 6422 6544 6456
rect 6544 6422 6578 6456
rect 6578 6422 6587 6456
rect 6535 6413 6587 6422
rect 8167 6456 8219 6465
rect 8167 6422 8176 6456
rect 8176 6422 8210 6456
rect 8210 6422 8219 6456
rect 8167 6413 8219 6422
rect 9799 6456 9851 6465
rect 9799 6422 9808 6456
rect 9808 6422 9842 6456
rect 9842 6422 9851 6456
rect 9799 6413 9851 6422
rect 11431 6456 11483 6465
rect 11431 6422 11440 6456
rect 11440 6422 11474 6456
rect 11474 6422 11483 6456
rect 11431 6413 11483 6422
rect 13063 6456 13115 6465
rect 13063 6422 13072 6456
rect 13072 6422 13106 6456
rect 13106 6422 13115 6456
rect 13063 6413 13115 6422
rect 7 6252 59 6261
rect 7 6218 16 6252
rect 16 6218 50 6252
rect 50 6218 59 6252
rect 7 6209 59 6218
rect 1639 6252 1691 6261
rect 1639 6218 1648 6252
rect 1648 6218 1682 6252
rect 1682 6218 1691 6252
rect 1639 6209 1691 6218
rect 3271 6252 3323 6261
rect 3271 6218 3280 6252
rect 3280 6218 3314 6252
rect 3314 6218 3323 6252
rect 3271 6209 3323 6218
rect 4903 6252 4955 6261
rect 4903 6218 4912 6252
rect 4912 6218 4946 6252
rect 4946 6218 4955 6252
rect 4903 6209 4955 6218
rect 6535 6252 6587 6261
rect 6535 6218 6544 6252
rect 6544 6218 6578 6252
rect 6578 6218 6587 6252
rect 6535 6209 6587 6218
rect 8167 6252 8219 6261
rect 8167 6218 8176 6252
rect 8176 6218 8210 6252
rect 8210 6218 8219 6252
rect 8167 6209 8219 6218
rect 9799 6252 9851 6261
rect 9799 6218 9808 6252
rect 9808 6218 9842 6252
rect 9842 6218 9851 6252
rect 9799 6209 9851 6218
rect 11431 6252 11483 6261
rect 11431 6218 11440 6252
rect 11440 6218 11474 6252
rect 11474 6218 11483 6252
rect 11431 6209 11483 6218
rect 13063 6252 13115 6261
rect 13063 6218 13072 6252
rect 13072 6218 13106 6252
rect 13106 6218 13115 6252
rect 13063 6209 13115 6218
rect 218 6098 270 6107
rect 218 6064 227 6098
rect 227 6064 261 6098
rect 261 6064 270 6098
rect 218 6055 270 6064
rect 422 6098 474 6107
rect 422 6064 431 6098
rect 431 6064 465 6098
rect 465 6064 474 6098
rect 422 6055 474 6064
rect 626 6098 678 6107
rect 626 6064 635 6098
rect 635 6064 669 6098
rect 669 6064 678 6098
rect 626 6055 678 6064
rect 830 6098 882 6107
rect 830 6064 839 6098
rect 839 6064 873 6098
rect 873 6064 882 6098
rect 830 6055 882 6064
rect 1034 6098 1086 6107
rect 1034 6064 1043 6098
rect 1043 6064 1077 6098
rect 1077 6064 1086 6098
rect 1034 6055 1086 6064
rect 1238 6098 1290 6107
rect 1238 6064 1247 6098
rect 1247 6064 1281 6098
rect 1281 6064 1290 6098
rect 1238 6055 1290 6064
rect 1442 6098 1494 6107
rect 1442 6064 1451 6098
rect 1451 6064 1485 6098
rect 1485 6064 1494 6098
rect 1442 6055 1494 6064
rect 1646 6098 1698 6107
rect 1646 6064 1655 6098
rect 1655 6064 1689 6098
rect 1689 6064 1698 6098
rect 1646 6055 1698 6064
rect 1850 6098 1902 6107
rect 1850 6064 1859 6098
rect 1859 6064 1893 6098
rect 1893 6064 1902 6098
rect 1850 6055 1902 6064
rect 2054 6098 2106 6107
rect 2054 6064 2063 6098
rect 2063 6064 2097 6098
rect 2097 6064 2106 6098
rect 2054 6055 2106 6064
rect 2258 6098 2310 6107
rect 2258 6064 2267 6098
rect 2267 6064 2301 6098
rect 2301 6064 2310 6098
rect 2258 6055 2310 6064
rect 2462 6098 2514 6107
rect 2462 6064 2471 6098
rect 2471 6064 2505 6098
rect 2505 6064 2514 6098
rect 2462 6055 2514 6064
rect 2666 6098 2718 6107
rect 2666 6064 2675 6098
rect 2675 6064 2709 6098
rect 2709 6064 2718 6098
rect 2666 6055 2718 6064
rect 2870 6098 2922 6107
rect 2870 6064 2879 6098
rect 2879 6064 2913 6098
rect 2913 6064 2922 6098
rect 2870 6055 2922 6064
rect 3074 6098 3126 6107
rect 3074 6064 3083 6098
rect 3083 6064 3117 6098
rect 3117 6064 3126 6098
rect 3074 6055 3126 6064
rect 3278 6098 3330 6107
rect 3278 6064 3287 6098
rect 3287 6064 3321 6098
rect 3321 6064 3330 6098
rect 3278 6055 3330 6064
rect 3482 6098 3534 6107
rect 3482 6064 3491 6098
rect 3491 6064 3525 6098
rect 3525 6064 3534 6098
rect 3482 6055 3534 6064
rect 3686 6098 3738 6107
rect 3686 6064 3695 6098
rect 3695 6064 3729 6098
rect 3729 6064 3738 6098
rect 3686 6055 3738 6064
rect 3890 6098 3942 6107
rect 3890 6064 3899 6098
rect 3899 6064 3933 6098
rect 3933 6064 3942 6098
rect 3890 6055 3942 6064
rect 4094 6098 4146 6107
rect 4094 6064 4103 6098
rect 4103 6064 4137 6098
rect 4137 6064 4146 6098
rect 4094 6055 4146 6064
rect 4298 6098 4350 6107
rect 4298 6064 4307 6098
rect 4307 6064 4341 6098
rect 4341 6064 4350 6098
rect 4298 6055 4350 6064
rect 4502 6098 4554 6107
rect 4502 6064 4511 6098
rect 4511 6064 4545 6098
rect 4545 6064 4554 6098
rect 4502 6055 4554 6064
rect 4706 6098 4758 6107
rect 4706 6064 4715 6098
rect 4715 6064 4749 6098
rect 4749 6064 4758 6098
rect 4706 6055 4758 6064
rect 4910 6098 4962 6107
rect 4910 6064 4919 6098
rect 4919 6064 4953 6098
rect 4953 6064 4962 6098
rect 4910 6055 4962 6064
rect 5114 6098 5166 6107
rect 5114 6064 5123 6098
rect 5123 6064 5157 6098
rect 5157 6064 5166 6098
rect 5114 6055 5166 6064
rect 5318 6098 5370 6107
rect 5318 6064 5327 6098
rect 5327 6064 5361 6098
rect 5361 6064 5370 6098
rect 5318 6055 5370 6064
rect 5522 6098 5574 6107
rect 5522 6064 5531 6098
rect 5531 6064 5565 6098
rect 5565 6064 5574 6098
rect 5522 6055 5574 6064
rect 5726 6098 5778 6107
rect 5726 6064 5735 6098
rect 5735 6064 5769 6098
rect 5769 6064 5778 6098
rect 5726 6055 5778 6064
rect 5930 6098 5982 6107
rect 5930 6064 5939 6098
rect 5939 6064 5973 6098
rect 5973 6064 5982 6098
rect 5930 6055 5982 6064
rect 6134 6098 6186 6107
rect 6134 6064 6143 6098
rect 6143 6064 6177 6098
rect 6177 6064 6186 6098
rect 6134 6055 6186 6064
rect 6338 6098 6390 6107
rect 6338 6064 6347 6098
rect 6347 6064 6381 6098
rect 6381 6064 6390 6098
rect 6338 6055 6390 6064
rect 6542 6098 6594 6107
rect 6542 6064 6551 6098
rect 6551 6064 6585 6098
rect 6585 6064 6594 6098
rect 6542 6055 6594 6064
rect 6746 6098 6798 6107
rect 6746 6064 6755 6098
rect 6755 6064 6789 6098
rect 6789 6064 6798 6098
rect 6746 6055 6798 6064
rect 6950 6098 7002 6107
rect 6950 6064 6959 6098
rect 6959 6064 6993 6098
rect 6993 6064 7002 6098
rect 6950 6055 7002 6064
rect 7154 6098 7206 6107
rect 7154 6064 7163 6098
rect 7163 6064 7197 6098
rect 7197 6064 7206 6098
rect 7154 6055 7206 6064
rect 7358 6098 7410 6107
rect 7358 6064 7367 6098
rect 7367 6064 7401 6098
rect 7401 6064 7410 6098
rect 7358 6055 7410 6064
rect 7562 6098 7614 6107
rect 7562 6064 7571 6098
rect 7571 6064 7605 6098
rect 7605 6064 7614 6098
rect 7562 6055 7614 6064
rect 7766 6098 7818 6107
rect 7766 6064 7775 6098
rect 7775 6064 7809 6098
rect 7809 6064 7818 6098
rect 7766 6055 7818 6064
rect 7970 6098 8022 6107
rect 7970 6064 7979 6098
rect 7979 6064 8013 6098
rect 8013 6064 8022 6098
rect 7970 6055 8022 6064
rect 8174 6098 8226 6107
rect 8174 6064 8183 6098
rect 8183 6064 8217 6098
rect 8217 6064 8226 6098
rect 8174 6055 8226 6064
rect 8378 6098 8430 6107
rect 8378 6064 8387 6098
rect 8387 6064 8421 6098
rect 8421 6064 8430 6098
rect 8378 6055 8430 6064
rect 8582 6098 8634 6107
rect 8582 6064 8591 6098
rect 8591 6064 8625 6098
rect 8625 6064 8634 6098
rect 8582 6055 8634 6064
rect 8786 6098 8838 6107
rect 8786 6064 8795 6098
rect 8795 6064 8829 6098
rect 8829 6064 8838 6098
rect 8786 6055 8838 6064
rect 8990 6098 9042 6107
rect 8990 6064 8999 6098
rect 8999 6064 9033 6098
rect 9033 6064 9042 6098
rect 8990 6055 9042 6064
rect 9194 6098 9246 6107
rect 9194 6064 9203 6098
rect 9203 6064 9237 6098
rect 9237 6064 9246 6098
rect 9194 6055 9246 6064
rect 9398 6098 9450 6107
rect 9398 6064 9407 6098
rect 9407 6064 9441 6098
rect 9441 6064 9450 6098
rect 9398 6055 9450 6064
rect 9602 6098 9654 6107
rect 9602 6064 9611 6098
rect 9611 6064 9645 6098
rect 9645 6064 9654 6098
rect 9602 6055 9654 6064
rect 9806 6098 9858 6107
rect 9806 6064 9815 6098
rect 9815 6064 9849 6098
rect 9849 6064 9858 6098
rect 9806 6055 9858 6064
rect 10010 6098 10062 6107
rect 10010 6064 10019 6098
rect 10019 6064 10053 6098
rect 10053 6064 10062 6098
rect 10010 6055 10062 6064
rect 10214 6098 10266 6107
rect 10214 6064 10223 6098
rect 10223 6064 10257 6098
rect 10257 6064 10266 6098
rect 10214 6055 10266 6064
rect 10418 6098 10470 6107
rect 10418 6064 10427 6098
rect 10427 6064 10461 6098
rect 10461 6064 10470 6098
rect 10418 6055 10470 6064
rect 10622 6098 10674 6107
rect 10622 6064 10631 6098
rect 10631 6064 10665 6098
rect 10665 6064 10674 6098
rect 10622 6055 10674 6064
rect 10826 6098 10878 6107
rect 10826 6064 10835 6098
rect 10835 6064 10869 6098
rect 10869 6064 10878 6098
rect 10826 6055 10878 6064
rect 11030 6098 11082 6107
rect 11030 6064 11039 6098
rect 11039 6064 11073 6098
rect 11073 6064 11082 6098
rect 11030 6055 11082 6064
rect 11234 6098 11286 6107
rect 11234 6064 11243 6098
rect 11243 6064 11277 6098
rect 11277 6064 11286 6098
rect 11234 6055 11286 6064
rect 11438 6098 11490 6107
rect 11438 6064 11447 6098
rect 11447 6064 11481 6098
rect 11481 6064 11490 6098
rect 11438 6055 11490 6064
rect 11642 6098 11694 6107
rect 11642 6064 11651 6098
rect 11651 6064 11685 6098
rect 11685 6064 11694 6098
rect 11642 6055 11694 6064
rect 11846 6098 11898 6107
rect 11846 6064 11855 6098
rect 11855 6064 11889 6098
rect 11889 6064 11898 6098
rect 11846 6055 11898 6064
rect 12050 6098 12102 6107
rect 12050 6064 12059 6098
rect 12059 6064 12093 6098
rect 12093 6064 12102 6098
rect 12050 6055 12102 6064
rect 12254 6098 12306 6107
rect 12254 6064 12263 6098
rect 12263 6064 12297 6098
rect 12297 6064 12306 6098
rect 12254 6055 12306 6064
rect 12458 6098 12510 6107
rect 12458 6064 12467 6098
rect 12467 6064 12501 6098
rect 12501 6064 12510 6098
rect 12458 6055 12510 6064
rect 12662 6098 12714 6107
rect 12662 6064 12671 6098
rect 12671 6064 12705 6098
rect 12705 6064 12714 6098
rect 12662 6055 12714 6064
rect 12866 6098 12918 6107
rect 12866 6064 12875 6098
rect 12875 6064 12909 6098
rect 12909 6064 12918 6098
rect 12866 6055 12918 6064
rect 13084 6098 13136 6107
rect 13084 6064 13093 6098
rect 13093 6064 13127 6098
rect 13127 6064 13136 6098
rect 13084 6055 13136 6064
rect 7 5944 59 5953
rect 7 5910 16 5944
rect 16 5910 50 5944
rect 50 5910 59 5944
rect 7 5901 59 5910
rect 1639 5944 1691 5953
rect 1639 5910 1648 5944
rect 1648 5910 1682 5944
rect 1682 5910 1691 5944
rect 1639 5901 1691 5910
rect 3271 5944 3323 5953
rect 3271 5910 3280 5944
rect 3280 5910 3314 5944
rect 3314 5910 3323 5944
rect 3271 5901 3323 5910
rect 4903 5944 4955 5953
rect 4903 5910 4912 5944
rect 4912 5910 4946 5944
rect 4946 5910 4955 5944
rect 4903 5901 4955 5910
rect 6535 5944 6587 5953
rect 6535 5910 6544 5944
rect 6544 5910 6578 5944
rect 6578 5910 6587 5944
rect 6535 5901 6587 5910
rect 8167 5944 8219 5953
rect 8167 5910 8176 5944
rect 8176 5910 8210 5944
rect 8210 5910 8219 5944
rect 8167 5901 8219 5910
rect 9799 5944 9851 5953
rect 9799 5910 9808 5944
rect 9808 5910 9842 5944
rect 9842 5910 9851 5944
rect 9799 5901 9851 5910
rect 11431 5944 11483 5953
rect 11431 5910 11440 5944
rect 11440 5910 11474 5944
rect 11474 5910 11483 5944
rect 11431 5901 11483 5910
rect 13063 5944 13115 5953
rect 13063 5910 13072 5944
rect 13072 5910 13106 5944
rect 13106 5910 13115 5944
rect 13063 5901 13115 5910
rect 7 5740 59 5749
rect 7 5706 16 5740
rect 16 5706 50 5740
rect 50 5706 59 5740
rect 7 5697 59 5706
rect 1639 5740 1691 5749
rect 1639 5706 1648 5740
rect 1648 5706 1682 5740
rect 1682 5706 1691 5740
rect 1639 5697 1691 5706
rect 3271 5740 3323 5749
rect 3271 5706 3280 5740
rect 3280 5706 3314 5740
rect 3314 5706 3323 5740
rect 3271 5697 3323 5706
rect 4903 5740 4955 5749
rect 4903 5706 4912 5740
rect 4912 5706 4946 5740
rect 4946 5706 4955 5740
rect 4903 5697 4955 5706
rect 6535 5740 6587 5749
rect 6535 5706 6544 5740
rect 6544 5706 6578 5740
rect 6578 5706 6587 5740
rect 6535 5697 6587 5706
rect 8167 5740 8219 5749
rect 8167 5706 8176 5740
rect 8176 5706 8210 5740
rect 8210 5706 8219 5740
rect 8167 5697 8219 5706
rect 9799 5740 9851 5749
rect 9799 5706 9808 5740
rect 9808 5706 9842 5740
rect 9842 5706 9851 5740
rect 9799 5697 9851 5706
rect 11431 5740 11483 5749
rect 11431 5706 11440 5740
rect 11440 5706 11474 5740
rect 11474 5706 11483 5740
rect 11431 5697 11483 5706
rect 13063 5740 13115 5749
rect 13063 5706 13072 5740
rect 13072 5706 13106 5740
rect 13106 5706 13115 5740
rect 13063 5697 13115 5706
rect 7 5536 59 5545
rect 7 5502 16 5536
rect 16 5502 50 5536
rect 50 5502 59 5536
rect 7 5493 59 5502
rect 1639 5536 1691 5545
rect 1639 5502 1648 5536
rect 1648 5502 1682 5536
rect 1682 5502 1691 5536
rect 1639 5493 1691 5502
rect 3271 5536 3323 5545
rect 3271 5502 3280 5536
rect 3280 5502 3314 5536
rect 3314 5502 3323 5536
rect 3271 5493 3323 5502
rect 4903 5536 4955 5545
rect 4903 5502 4912 5536
rect 4912 5502 4946 5536
rect 4946 5502 4955 5536
rect 4903 5493 4955 5502
rect 6535 5536 6587 5545
rect 6535 5502 6544 5536
rect 6544 5502 6578 5536
rect 6578 5502 6587 5536
rect 6535 5493 6587 5502
rect 8167 5536 8219 5545
rect 8167 5502 8176 5536
rect 8176 5502 8210 5536
rect 8210 5502 8219 5536
rect 8167 5493 8219 5502
rect 9799 5536 9851 5545
rect 9799 5502 9808 5536
rect 9808 5502 9842 5536
rect 9842 5502 9851 5536
rect 9799 5493 9851 5502
rect 11431 5536 11483 5545
rect 11431 5502 11440 5536
rect 11440 5502 11474 5536
rect 11474 5502 11483 5536
rect 11431 5493 11483 5502
rect 13063 5536 13115 5545
rect 13063 5502 13072 5536
rect 13072 5502 13106 5536
rect 13106 5502 13115 5536
rect 13063 5493 13115 5502
rect 7 5332 59 5341
rect 7 5298 16 5332
rect 16 5298 50 5332
rect 50 5298 59 5332
rect 7 5289 59 5298
rect 1639 5332 1691 5341
rect 1639 5298 1648 5332
rect 1648 5298 1682 5332
rect 1682 5298 1691 5332
rect 1639 5289 1691 5298
rect 3271 5332 3323 5341
rect 3271 5298 3280 5332
rect 3280 5298 3314 5332
rect 3314 5298 3323 5332
rect 3271 5289 3323 5298
rect 4903 5332 4955 5341
rect 4903 5298 4912 5332
rect 4912 5298 4946 5332
rect 4946 5298 4955 5332
rect 4903 5289 4955 5298
rect 6535 5332 6587 5341
rect 6535 5298 6544 5332
rect 6544 5298 6578 5332
rect 6578 5298 6587 5332
rect 6535 5289 6587 5298
rect 8167 5332 8219 5341
rect 8167 5298 8176 5332
rect 8176 5298 8210 5332
rect 8210 5298 8219 5332
rect 8167 5289 8219 5298
rect 9799 5332 9851 5341
rect 9799 5298 9808 5332
rect 9808 5298 9842 5332
rect 9842 5298 9851 5332
rect 9799 5289 9851 5298
rect 11431 5332 11483 5341
rect 11431 5298 11440 5332
rect 11440 5298 11474 5332
rect 11474 5298 11483 5332
rect 11431 5289 11483 5298
rect 13063 5332 13115 5341
rect 13063 5298 13072 5332
rect 13072 5298 13106 5332
rect 13106 5298 13115 5332
rect 13063 5289 13115 5298
rect 7 5128 59 5137
rect 7 5094 16 5128
rect 16 5094 50 5128
rect 50 5094 59 5128
rect 7 5085 59 5094
rect 1639 5128 1691 5137
rect 1639 5094 1648 5128
rect 1648 5094 1682 5128
rect 1682 5094 1691 5128
rect 1639 5085 1691 5094
rect 3271 5128 3323 5137
rect 3271 5094 3280 5128
rect 3280 5094 3314 5128
rect 3314 5094 3323 5128
rect 3271 5085 3323 5094
rect 4903 5128 4955 5137
rect 4903 5094 4912 5128
rect 4912 5094 4946 5128
rect 4946 5094 4955 5128
rect 4903 5085 4955 5094
rect 6535 5128 6587 5137
rect 6535 5094 6544 5128
rect 6544 5094 6578 5128
rect 6578 5094 6587 5128
rect 6535 5085 6587 5094
rect 8167 5128 8219 5137
rect 8167 5094 8176 5128
rect 8176 5094 8210 5128
rect 8210 5094 8219 5128
rect 8167 5085 8219 5094
rect 9799 5128 9851 5137
rect 9799 5094 9808 5128
rect 9808 5094 9842 5128
rect 9842 5094 9851 5128
rect 9799 5085 9851 5094
rect 11431 5128 11483 5137
rect 11431 5094 11440 5128
rect 11440 5094 11474 5128
rect 11474 5094 11483 5128
rect 11431 5085 11483 5094
rect 13063 5128 13115 5137
rect 13063 5094 13072 5128
rect 13072 5094 13106 5128
rect 13106 5094 13115 5128
rect 13063 5085 13115 5094
rect 7 4924 59 4933
rect 7 4890 16 4924
rect 16 4890 50 4924
rect 50 4890 59 4924
rect 7 4881 59 4890
rect 1639 4924 1691 4933
rect 1639 4890 1648 4924
rect 1648 4890 1682 4924
rect 1682 4890 1691 4924
rect 1639 4881 1691 4890
rect 3271 4924 3323 4933
rect 3271 4890 3280 4924
rect 3280 4890 3314 4924
rect 3314 4890 3323 4924
rect 3271 4881 3323 4890
rect 4903 4924 4955 4933
rect 4903 4890 4912 4924
rect 4912 4890 4946 4924
rect 4946 4890 4955 4924
rect 4903 4881 4955 4890
rect 6535 4924 6587 4933
rect 6535 4890 6544 4924
rect 6544 4890 6578 4924
rect 6578 4890 6587 4924
rect 6535 4881 6587 4890
rect 8167 4924 8219 4933
rect 8167 4890 8176 4924
rect 8176 4890 8210 4924
rect 8210 4890 8219 4924
rect 8167 4881 8219 4890
rect 9799 4924 9851 4933
rect 9799 4890 9808 4924
rect 9808 4890 9842 4924
rect 9842 4890 9851 4924
rect 9799 4881 9851 4890
rect 11431 4924 11483 4933
rect 11431 4890 11440 4924
rect 11440 4890 11474 4924
rect 11474 4890 11483 4924
rect 11431 4881 11483 4890
rect 13063 4924 13115 4933
rect 13063 4890 13072 4924
rect 13072 4890 13106 4924
rect 13106 4890 13115 4924
rect 13063 4881 13115 4890
rect 7 4720 59 4729
rect 7 4686 16 4720
rect 16 4686 50 4720
rect 50 4686 59 4720
rect 7 4677 59 4686
rect 1639 4720 1691 4729
rect 1639 4686 1648 4720
rect 1648 4686 1682 4720
rect 1682 4686 1691 4720
rect 1639 4677 1691 4686
rect 3271 4720 3323 4729
rect 3271 4686 3280 4720
rect 3280 4686 3314 4720
rect 3314 4686 3323 4720
rect 3271 4677 3323 4686
rect 4903 4720 4955 4729
rect 4903 4686 4912 4720
rect 4912 4686 4946 4720
rect 4946 4686 4955 4720
rect 4903 4677 4955 4686
rect 6535 4720 6587 4729
rect 6535 4686 6544 4720
rect 6544 4686 6578 4720
rect 6578 4686 6587 4720
rect 6535 4677 6587 4686
rect 8167 4720 8219 4729
rect 8167 4686 8176 4720
rect 8176 4686 8210 4720
rect 8210 4686 8219 4720
rect 8167 4677 8219 4686
rect 9799 4720 9851 4729
rect 9799 4686 9808 4720
rect 9808 4686 9842 4720
rect 9842 4686 9851 4720
rect 9799 4677 9851 4686
rect 11431 4720 11483 4729
rect 11431 4686 11440 4720
rect 11440 4686 11474 4720
rect 11474 4686 11483 4720
rect 11431 4677 11483 4686
rect 13063 4720 13115 4729
rect 13063 4686 13072 4720
rect 13072 4686 13106 4720
rect 13106 4686 13115 4720
rect 13063 4677 13115 4686
rect 7 4516 59 4525
rect 7 4482 16 4516
rect 16 4482 50 4516
rect 50 4482 59 4516
rect 7 4473 59 4482
rect 1639 4516 1691 4525
rect 1639 4482 1648 4516
rect 1648 4482 1682 4516
rect 1682 4482 1691 4516
rect 1639 4473 1691 4482
rect 3271 4516 3323 4525
rect 3271 4482 3280 4516
rect 3280 4482 3314 4516
rect 3314 4482 3323 4516
rect 3271 4473 3323 4482
rect 4903 4516 4955 4525
rect 4903 4482 4912 4516
rect 4912 4482 4946 4516
rect 4946 4482 4955 4516
rect 4903 4473 4955 4482
rect 6535 4516 6587 4525
rect 6535 4482 6544 4516
rect 6544 4482 6578 4516
rect 6578 4482 6587 4516
rect 6535 4473 6587 4482
rect 8167 4516 8219 4525
rect 8167 4482 8176 4516
rect 8176 4482 8210 4516
rect 8210 4482 8219 4516
rect 8167 4473 8219 4482
rect 9799 4516 9851 4525
rect 9799 4482 9808 4516
rect 9808 4482 9842 4516
rect 9842 4482 9851 4516
rect 9799 4473 9851 4482
rect 11431 4516 11483 4525
rect 11431 4482 11440 4516
rect 11440 4482 11474 4516
rect 11474 4482 11483 4516
rect 11431 4473 11483 4482
rect 13063 4516 13115 4525
rect 13063 4482 13072 4516
rect 13072 4482 13106 4516
rect 13106 4482 13115 4516
rect 13063 4473 13115 4482
rect 218 4362 270 4371
rect 218 4328 227 4362
rect 227 4328 261 4362
rect 261 4328 270 4362
rect 218 4319 270 4328
rect 422 4362 474 4371
rect 422 4328 431 4362
rect 431 4328 465 4362
rect 465 4328 474 4362
rect 422 4319 474 4328
rect 626 4362 678 4371
rect 626 4328 635 4362
rect 635 4328 669 4362
rect 669 4328 678 4362
rect 626 4319 678 4328
rect 830 4362 882 4371
rect 830 4328 839 4362
rect 839 4328 873 4362
rect 873 4328 882 4362
rect 830 4319 882 4328
rect 1034 4362 1086 4371
rect 1034 4328 1043 4362
rect 1043 4328 1077 4362
rect 1077 4328 1086 4362
rect 1034 4319 1086 4328
rect 1238 4362 1290 4371
rect 1238 4328 1247 4362
rect 1247 4328 1281 4362
rect 1281 4328 1290 4362
rect 1238 4319 1290 4328
rect 1442 4362 1494 4371
rect 1442 4328 1451 4362
rect 1451 4328 1485 4362
rect 1485 4328 1494 4362
rect 1442 4319 1494 4328
rect 1646 4362 1698 4371
rect 1646 4328 1655 4362
rect 1655 4328 1689 4362
rect 1689 4328 1698 4362
rect 1646 4319 1698 4328
rect 1850 4362 1902 4371
rect 1850 4328 1859 4362
rect 1859 4328 1893 4362
rect 1893 4328 1902 4362
rect 1850 4319 1902 4328
rect 2054 4362 2106 4371
rect 2054 4328 2063 4362
rect 2063 4328 2097 4362
rect 2097 4328 2106 4362
rect 2054 4319 2106 4328
rect 2258 4362 2310 4371
rect 2258 4328 2267 4362
rect 2267 4328 2301 4362
rect 2301 4328 2310 4362
rect 2258 4319 2310 4328
rect 2462 4362 2514 4371
rect 2462 4328 2471 4362
rect 2471 4328 2505 4362
rect 2505 4328 2514 4362
rect 2462 4319 2514 4328
rect 2666 4362 2718 4371
rect 2666 4328 2675 4362
rect 2675 4328 2709 4362
rect 2709 4328 2718 4362
rect 2666 4319 2718 4328
rect 2870 4362 2922 4371
rect 2870 4328 2879 4362
rect 2879 4328 2913 4362
rect 2913 4328 2922 4362
rect 2870 4319 2922 4328
rect 3074 4362 3126 4371
rect 3074 4328 3083 4362
rect 3083 4328 3117 4362
rect 3117 4328 3126 4362
rect 3074 4319 3126 4328
rect 3278 4362 3330 4371
rect 3278 4328 3287 4362
rect 3287 4328 3321 4362
rect 3321 4328 3330 4362
rect 3278 4319 3330 4328
rect 3482 4362 3534 4371
rect 3482 4328 3491 4362
rect 3491 4328 3525 4362
rect 3525 4328 3534 4362
rect 3482 4319 3534 4328
rect 3686 4362 3738 4371
rect 3686 4328 3695 4362
rect 3695 4328 3729 4362
rect 3729 4328 3738 4362
rect 3686 4319 3738 4328
rect 3890 4362 3942 4371
rect 3890 4328 3899 4362
rect 3899 4328 3933 4362
rect 3933 4328 3942 4362
rect 3890 4319 3942 4328
rect 4094 4362 4146 4371
rect 4094 4328 4103 4362
rect 4103 4328 4137 4362
rect 4137 4328 4146 4362
rect 4094 4319 4146 4328
rect 4298 4362 4350 4371
rect 4298 4328 4307 4362
rect 4307 4328 4341 4362
rect 4341 4328 4350 4362
rect 4298 4319 4350 4328
rect 4502 4362 4554 4371
rect 4502 4328 4511 4362
rect 4511 4328 4545 4362
rect 4545 4328 4554 4362
rect 4502 4319 4554 4328
rect 4706 4362 4758 4371
rect 4706 4328 4715 4362
rect 4715 4328 4749 4362
rect 4749 4328 4758 4362
rect 4706 4319 4758 4328
rect 4910 4362 4962 4371
rect 4910 4328 4919 4362
rect 4919 4328 4953 4362
rect 4953 4328 4962 4362
rect 4910 4319 4962 4328
rect 5114 4362 5166 4371
rect 5114 4328 5123 4362
rect 5123 4328 5157 4362
rect 5157 4328 5166 4362
rect 5114 4319 5166 4328
rect 5318 4362 5370 4371
rect 5318 4328 5327 4362
rect 5327 4328 5361 4362
rect 5361 4328 5370 4362
rect 5318 4319 5370 4328
rect 5522 4362 5574 4371
rect 5522 4328 5531 4362
rect 5531 4328 5565 4362
rect 5565 4328 5574 4362
rect 5522 4319 5574 4328
rect 5726 4362 5778 4371
rect 5726 4328 5735 4362
rect 5735 4328 5769 4362
rect 5769 4328 5778 4362
rect 5726 4319 5778 4328
rect 5930 4362 5982 4371
rect 5930 4328 5939 4362
rect 5939 4328 5973 4362
rect 5973 4328 5982 4362
rect 5930 4319 5982 4328
rect 6134 4362 6186 4371
rect 6134 4328 6143 4362
rect 6143 4328 6177 4362
rect 6177 4328 6186 4362
rect 6134 4319 6186 4328
rect 6338 4362 6390 4371
rect 6338 4328 6347 4362
rect 6347 4328 6381 4362
rect 6381 4328 6390 4362
rect 6338 4319 6390 4328
rect 6542 4362 6594 4371
rect 6542 4328 6551 4362
rect 6551 4328 6585 4362
rect 6585 4328 6594 4362
rect 6542 4319 6594 4328
rect 6746 4362 6798 4371
rect 6746 4328 6755 4362
rect 6755 4328 6789 4362
rect 6789 4328 6798 4362
rect 6746 4319 6798 4328
rect 6950 4362 7002 4371
rect 6950 4328 6959 4362
rect 6959 4328 6993 4362
rect 6993 4328 7002 4362
rect 6950 4319 7002 4328
rect 7154 4362 7206 4371
rect 7154 4328 7163 4362
rect 7163 4328 7197 4362
rect 7197 4328 7206 4362
rect 7154 4319 7206 4328
rect 7358 4362 7410 4371
rect 7358 4328 7367 4362
rect 7367 4328 7401 4362
rect 7401 4328 7410 4362
rect 7358 4319 7410 4328
rect 7562 4362 7614 4371
rect 7562 4328 7571 4362
rect 7571 4328 7605 4362
rect 7605 4328 7614 4362
rect 7562 4319 7614 4328
rect 7766 4362 7818 4371
rect 7766 4328 7775 4362
rect 7775 4328 7809 4362
rect 7809 4328 7818 4362
rect 7766 4319 7818 4328
rect 7970 4362 8022 4371
rect 7970 4328 7979 4362
rect 7979 4328 8013 4362
rect 8013 4328 8022 4362
rect 7970 4319 8022 4328
rect 8174 4362 8226 4371
rect 8174 4328 8183 4362
rect 8183 4328 8217 4362
rect 8217 4328 8226 4362
rect 8174 4319 8226 4328
rect 8378 4362 8430 4371
rect 8378 4328 8387 4362
rect 8387 4328 8421 4362
rect 8421 4328 8430 4362
rect 8378 4319 8430 4328
rect 8582 4362 8634 4371
rect 8582 4328 8591 4362
rect 8591 4328 8625 4362
rect 8625 4328 8634 4362
rect 8582 4319 8634 4328
rect 8786 4362 8838 4371
rect 8786 4328 8795 4362
rect 8795 4328 8829 4362
rect 8829 4328 8838 4362
rect 8786 4319 8838 4328
rect 8990 4362 9042 4371
rect 8990 4328 8999 4362
rect 8999 4328 9033 4362
rect 9033 4328 9042 4362
rect 8990 4319 9042 4328
rect 9194 4362 9246 4371
rect 9194 4328 9203 4362
rect 9203 4328 9237 4362
rect 9237 4328 9246 4362
rect 9194 4319 9246 4328
rect 9398 4362 9450 4371
rect 9398 4328 9407 4362
rect 9407 4328 9441 4362
rect 9441 4328 9450 4362
rect 9398 4319 9450 4328
rect 9602 4362 9654 4371
rect 9602 4328 9611 4362
rect 9611 4328 9645 4362
rect 9645 4328 9654 4362
rect 9602 4319 9654 4328
rect 9806 4362 9858 4371
rect 9806 4328 9815 4362
rect 9815 4328 9849 4362
rect 9849 4328 9858 4362
rect 9806 4319 9858 4328
rect 10010 4362 10062 4371
rect 10010 4328 10019 4362
rect 10019 4328 10053 4362
rect 10053 4328 10062 4362
rect 10010 4319 10062 4328
rect 10214 4362 10266 4371
rect 10214 4328 10223 4362
rect 10223 4328 10257 4362
rect 10257 4328 10266 4362
rect 10214 4319 10266 4328
rect 10418 4362 10470 4371
rect 10418 4328 10427 4362
rect 10427 4328 10461 4362
rect 10461 4328 10470 4362
rect 10418 4319 10470 4328
rect 10622 4362 10674 4371
rect 10622 4328 10631 4362
rect 10631 4328 10665 4362
rect 10665 4328 10674 4362
rect 10622 4319 10674 4328
rect 10826 4362 10878 4371
rect 10826 4328 10835 4362
rect 10835 4328 10869 4362
rect 10869 4328 10878 4362
rect 10826 4319 10878 4328
rect 11030 4362 11082 4371
rect 11030 4328 11039 4362
rect 11039 4328 11073 4362
rect 11073 4328 11082 4362
rect 11030 4319 11082 4328
rect 11234 4362 11286 4371
rect 11234 4328 11243 4362
rect 11243 4328 11277 4362
rect 11277 4328 11286 4362
rect 11234 4319 11286 4328
rect 11438 4362 11490 4371
rect 11438 4328 11447 4362
rect 11447 4328 11481 4362
rect 11481 4328 11490 4362
rect 11438 4319 11490 4328
rect 11642 4362 11694 4371
rect 11642 4328 11651 4362
rect 11651 4328 11685 4362
rect 11685 4328 11694 4362
rect 11642 4319 11694 4328
rect 11846 4362 11898 4371
rect 11846 4328 11855 4362
rect 11855 4328 11889 4362
rect 11889 4328 11898 4362
rect 11846 4319 11898 4328
rect 12050 4362 12102 4371
rect 12050 4328 12059 4362
rect 12059 4328 12093 4362
rect 12093 4328 12102 4362
rect 12050 4319 12102 4328
rect 12254 4362 12306 4371
rect 12254 4328 12263 4362
rect 12263 4328 12297 4362
rect 12297 4328 12306 4362
rect 12254 4319 12306 4328
rect 12458 4362 12510 4371
rect 12458 4328 12467 4362
rect 12467 4328 12501 4362
rect 12501 4328 12510 4362
rect 12458 4319 12510 4328
rect 12662 4362 12714 4371
rect 12662 4328 12671 4362
rect 12671 4328 12705 4362
rect 12705 4328 12714 4362
rect 12662 4319 12714 4328
rect 12866 4362 12918 4371
rect 12866 4328 12875 4362
rect 12875 4328 12909 4362
rect 12909 4328 12918 4362
rect 12866 4319 12918 4328
rect 13084 4362 13136 4371
rect 13084 4328 13093 4362
rect 13093 4328 13127 4362
rect 13127 4328 13136 4362
rect 13084 4319 13136 4328
rect 7 4208 59 4217
rect 7 4174 16 4208
rect 16 4174 50 4208
rect 50 4174 59 4208
rect 7 4165 59 4174
rect 1639 4208 1691 4217
rect 1639 4174 1648 4208
rect 1648 4174 1682 4208
rect 1682 4174 1691 4208
rect 1639 4165 1691 4174
rect 3271 4208 3323 4217
rect 3271 4174 3280 4208
rect 3280 4174 3314 4208
rect 3314 4174 3323 4208
rect 3271 4165 3323 4174
rect 4903 4208 4955 4217
rect 4903 4174 4912 4208
rect 4912 4174 4946 4208
rect 4946 4174 4955 4208
rect 4903 4165 4955 4174
rect 6535 4208 6587 4217
rect 6535 4174 6544 4208
rect 6544 4174 6578 4208
rect 6578 4174 6587 4208
rect 6535 4165 6587 4174
rect 8167 4208 8219 4217
rect 8167 4174 8176 4208
rect 8176 4174 8210 4208
rect 8210 4174 8219 4208
rect 8167 4165 8219 4174
rect 9799 4208 9851 4217
rect 9799 4174 9808 4208
rect 9808 4174 9842 4208
rect 9842 4174 9851 4208
rect 9799 4165 9851 4174
rect 11431 4208 11483 4217
rect 11431 4174 11440 4208
rect 11440 4174 11474 4208
rect 11474 4174 11483 4208
rect 11431 4165 11483 4174
rect 13063 4208 13115 4217
rect 13063 4174 13072 4208
rect 13072 4174 13106 4208
rect 13106 4174 13115 4208
rect 13063 4165 13115 4174
rect 7 4004 59 4013
rect 7 3970 16 4004
rect 16 3970 50 4004
rect 50 3970 59 4004
rect 7 3961 59 3970
rect 1639 4004 1691 4013
rect 1639 3970 1648 4004
rect 1648 3970 1682 4004
rect 1682 3970 1691 4004
rect 1639 3961 1691 3970
rect 3271 4004 3323 4013
rect 3271 3970 3280 4004
rect 3280 3970 3314 4004
rect 3314 3970 3323 4004
rect 3271 3961 3323 3970
rect 4903 4004 4955 4013
rect 4903 3970 4912 4004
rect 4912 3970 4946 4004
rect 4946 3970 4955 4004
rect 4903 3961 4955 3970
rect 6535 4004 6587 4013
rect 6535 3970 6544 4004
rect 6544 3970 6578 4004
rect 6578 3970 6587 4004
rect 6535 3961 6587 3970
rect 8167 4004 8219 4013
rect 8167 3970 8176 4004
rect 8176 3970 8210 4004
rect 8210 3970 8219 4004
rect 8167 3961 8219 3970
rect 9799 4004 9851 4013
rect 9799 3970 9808 4004
rect 9808 3970 9842 4004
rect 9842 3970 9851 4004
rect 9799 3961 9851 3970
rect 11431 4004 11483 4013
rect 11431 3970 11440 4004
rect 11440 3970 11474 4004
rect 11474 3970 11483 4004
rect 11431 3961 11483 3970
rect 13063 4004 13115 4013
rect 13063 3970 13072 4004
rect 13072 3970 13106 4004
rect 13106 3970 13115 4004
rect 13063 3961 13115 3970
rect 7 3800 59 3809
rect 7 3766 16 3800
rect 16 3766 50 3800
rect 50 3766 59 3800
rect 7 3757 59 3766
rect 1639 3800 1691 3809
rect 1639 3766 1648 3800
rect 1648 3766 1682 3800
rect 1682 3766 1691 3800
rect 1639 3757 1691 3766
rect 3271 3800 3323 3809
rect 3271 3766 3280 3800
rect 3280 3766 3314 3800
rect 3314 3766 3323 3800
rect 3271 3757 3323 3766
rect 4903 3800 4955 3809
rect 4903 3766 4912 3800
rect 4912 3766 4946 3800
rect 4946 3766 4955 3800
rect 4903 3757 4955 3766
rect 6535 3800 6587 3809
rect 6535 3766 6544 3800
rect 6544 3766 6578 3800
rect 6578 3766 6587 3800
rect 6535 3757 6587 3766
rect 8167 3800 8219 3809
rect 8167 3766 8176 3800
rect 8176 3766 8210 3800
rect 8210 3766 8219 3800
rect 8167 3757 8219 3766
rect 9799 3800 9851 3809
rect 9799 3766 9808 3800
rect 9808 3766 9842 3800
rect 9842 3766 9851 3800
rect 9799 3757 9851 3766
rect 11431 3800 11483 3809
rect 11431 3766 11440 3800
rect 11440 3766 11474 3800
rect 11474 3766 11483 3800
rect 11431 3757 11483 3766
rect 13063 3800 13115 3809
rect 13063 3766 13072 3800
rect 13072 3766 13106 3800
rect 13106 3766 13115 3800
rect 13063 3757 13115 3766
rect 7 3596 59 3605
rect 7 3562 16 3596
rect 16 3562 50 3596
rect 50 3562 59 3596
rect 7 3553 59 3562
rect 1639 3596 1691 3605
rect 1639 3562 1648 3596
rect 1648 3562 1682 3596
rect 1682 3562 1691 3596
rect 1639 3553 1691 3562
rect 3271 3596 3323 3605
rect 3271 3562 3280 3596
rect 3280 3562 3314 3596
rect 3314 3562 3323 3596
rect 3271 3553 3323 3562
rect 4903 3596 4955 3605
rect 4903 3562 4912 3596
rect 4912 3562 4946 3596
rect 4946 3562 4955 3596
rect 4903 3553 4955 3562
rect 6535 3596 6587 3605
rect 6535 3562 6544 3596
rect 6544 3562 6578 3596
rect 6578 3562 6587 3596
rect 6535 3553 6587 3562
rect 8167 3596 8219 3605
rect 8167 3562 8176 3596
rect 8176 3562 8210 3596
rect 8210 3562 8219 3596
rect 8167 3553 8219 3562
rect 9799 3596 9851 3605
rect 9799 3562 9808 3596
rect 9808 3562 9842 3596
rect 9842 3562 9851 3596
rect 9799 3553 9851 3562
rect 11431 3596 11483 3605
rect 11431 3562 11440 3596
rect 11440 3562 11474 3596
rect 11474 3562 11483 3596
rect 11431 3553 11483 3562
rect 13063 3596 13115 3605
rect 13063 3562 13072 3596
rect 13072 3562 13106 3596
rect 13106 3562 13115 3596
rect 13063 3553 13115 3562
rect 7 3392 59 3401
rect 7 3358 16 3392
rect 16 3358 50 3392
rect 50 3358 59 3392
rect 7 3349 59 3358
rect 1639 3392 1691 3401
rect 1639 3358 1648 3392
rect 1648 3358 1682 3392
rect 1682 3358 1691 3392
rect 1639 3349 1691 3358
rect 3271 3392 3323 3401
rect 3271 3358 3280 3392
rect 3280 3358 3314 3392
rect 3314 3358 3323 3392
rect 3271 3349 3323 3358
rect 4903 3392 4955 3401
rect 4903 3358 4912 3392
rect 4912 3358 4946 3392
rect 4946 3358 4955 3392
rect 4903 3349 4955 3358
rect 6535 3392 6587 3401
rect 6535 3358 6544 3392
rect 6544 3358 6578 3392
rect 6578 3358 6587 3392
rect 6535 3349 6587 3358
rect 8167 3392 8219 3401
rect 8167 3358 8176 3392
rect 8176 3358 8210 3392
rect 8210 3358 8219 3392
rect 8167 3349 8219 3358
rect 9799 3392 9851 3401
rect 9799 3358 9808 3392
rect 9808 3358 9842 3392
rect 9842 3358 9851 3392
rect 9799 3349 9851 3358
rect 11431 3392 11483 3401
rect 11431 3358 11440 3392
rect 11440 3358 11474 3392
rect 11474 3358 11483 3392
rect 11431 3349 11483 3358
rect 13063 3392 13115 3401
rect 13063 3358 13072 3392
rect 13072 3358 13106 3392
rect 13106 3358 13115 3392
rect 13063 3349 13115 3358
rect 7 3188 59 3197
rect 7 3154 16 3188
rect 16 3154 50 3188
rect 50 3154 59 3188
rect 7 3145 59 3154
rect 1639 3188 1691 3197
rect 1639 3154 1648 3188
rect 1648 3154 1682 3188
rect 1682 3154 1691 3188
rect 1639 3145 1691 3154
rect 3271 3188 3323 3197
rect 3271 3154 3280 3188
rect 3280 3154 3314 3188
rect 3314 3154 3323 3188
rect 3271 3145 3323 3154
rect 4903 3188 4955 3197
rect 4903 3154 4912 3188
rect 4912 3154 4946 3188
rect 4946 3154 4955 3188
rect 4903 3145 4955 3154
rect 6535 3188 6587 3197
rect 6535 3154 6544 3188
rect 6544 3154 6578 3188
rect 6578 3154 6587 3188
rect 6535 3145 6587 3154
rect 8167 3188 8219 3197
rect 8167 3154 8176 3188
rect 8176 3154 8210 3188
rect 8210 3154 8219 3188
rect 8167 3145 8219 3154
rect 9799 3188 9851 3197
rect 9799 3154 9808 3188
rect 9808 3154 9842 3188
rect 9842 3154 9851 3188
rect 9799 3145 9851 3154
rect 11431 3188 11483 3197
rect 11431 3154 11440 3188
rect 11440 3154 11474 3188
rect 11474 3154 11483 3188
rect 11431 3145 11483 3154
rect 13063 3188 13115 3197
rect 13063 3154 13072 3188
rect 13072 3154 13106 3188
rect 13106 3154 13115 3188
rect 13063 3145 13115 3154
rect 7 2984 59 2993
rect 7 2950 16 2984
rect 16 2950 50 2984
rect 50 2950 59 2984
rect 7 2941 59 2950
rect 1639 2984 1691 2993
rect 1639 2950 1648 2984
rect 1648 2950 1682 2984
rect 1682 2950 1691 2984
rect 1639 2941 1691 2950
rect 3271 2984 3323 2993
rect 3271 2950 3280 2984
rect 3280 2950 3314 2984
rect 3314 2950 3323 2984
rect 3271 2941 3323 2950
rect 4903 2984 4955 2993
rect 4903 2950 4912 2984
rect 4912 2950 4946 2984
rect 4946 2950 4955 2984
rect 4903 2941 4955 2950
rect 6535 2984 6587 2993
rect 6535 2950 6544 2984
rect 6544 2950 6578 2984
rect 6578 2950 6587 2984
rect 6535 2941 6587 2950
rect 8167 2984 8219 2993
rect 8167 2950 8176 2984
rect 8176 2950 8210 2984
rect 8210 2950 8219 2984
rect 8167 2941 8219 2950
rect 9799 2984 9851 2993
rect 9799 2950 9808 2984
rect 9808 2950 9842 2984
rect 9842 2950 9851 2984
rect 9799 2941 9851 2950
rect 11431 2984 11483 2993
rect 11431 2950 11440 2984
rect 11440 2950 11474 2984
rect 11474 2950 11483 2984
rect 11431 2941 11483 2950
rect 13063 2984 13115 2993
rect 13063 2950 13072 2984
rect 13072 2950 13106 2984
rect 13106 2950 13115 2984
rect 13063 2941 13115 2950
rect 7 2780 59 2789
rect 7 2746 16 2780
rect 16 2746 50 2780
rect 50 2746 59 2780
rect 7 2737 59 2746
rect 1639 2780 1691 2789
rect 1639 2746 1648 2780
rect 1648 2746 1682 2780
rect 1682 2746 1691 2780
rect 1639 2737 1691 2746
rect 3271 2780 3323 2789
rect 3271 2746 3280 2780
rect 3280 2746 3314 2780
rect 3314 2746 3323 2780
rect 3271 2737 3323 2746
rect 4903 2780 4955 2789
rect 4903 2746 4912 2780
rect 4912 2746 4946 2780
rect 4946 2746 4955 2780
rect 4903 2737 4955 2746
rect 6535 2780 6587 2789
rect 6535 2746 6544 2780
rect 6544 2746 6578 2780
rect 6578 2746 6587 2780
rect 6535 2737 6587 2746
rect 8167 2780 8219 2789
rect 8167 2746 8176 2780
rect 8176 2746 8210 2780
rect 8210 2746 8219 2780
rect 8167 2737 8219 2746
rect 9799 2780 9851 2789
rect 9799 2746 9808 2780
rect 9808 2746 9842 2780
rect 9842 2746 9851 2780
rect 9799 2737 9851 2746
rect 11431 2780 11483 2789
rect 11431 2746 11440 2780
rect 11440 2746 11474 2780
rect 11474 2746 11483 2780
rect 11431 2737 11483 2746
rect 13063 2780 13115 2789
rect 13063 2746 13072 2780
rect 13072 2746 13106 2780
rect 13106 2746 13115 2780
rect 13063 2737 13115 2746
rect 218 2626 270 2635
rect 218 2592 227 2626
rect 227 2592 261 2626
rect 261 2592 270 2626
rect 218 2583 270 2592
rect 422 2626 474 2635
rect 422 2592 431 2626
rect 431 2592 465 2626
rect 465 2592 474 2626
rect 422 2583 474 2592
rect 626 2626 678 2635
rect 626 2592 635 2626
rect 635 2592 669 2626
rect 669 2592 678 2626
rect 626 2583 678 2592
rect 830 2626 882 2635
rect 830 2592 839 2626
rect 839 2592 873 2626
rect 873 2592 882 2626
rect 830 2583 882 2592
rect 1034 2626 1086 2635
rect 1034 2592 1043 2626
rect 1043 2592 1077 2626
rect 1077 2592 1086 2626
rect 1034 2583 1086 2592
rect 1238 2626 1290 2635
rect 1238 2592 1247 2626
rect 1247 2592 1281 2626
rect 1281 2592 1290 2626
rect 1238 2583 1290 2592
rect 1442 2626 1494 2635
rect 1442 2592 1451 2626
rect 1451 2592 1485 2626
rect 1485 2592 1494 2626
rect 1442 2583 1494 2592
rect 1646 2626 1698 2635
rect 1646 2592 1655 2626
rect 1655 2592 1689 2626
rect 1689 2592 1698 2626
rect 1646 2583 1698 2592
rect 1850 2626 1902 2635
rect 1850 2592 1859 2626
rect 1859 2592 1893 2626
rect 1893 2592 1902 2626
rect 1850 2583 1902 2592
rect 2054 2626 2106 2635
rect 2054 2592 2063 2626
rect 2063 2592 2097 2626
rect 2097 2592 2106 2626
rect 2054 2583 2106 2592
rect 2258 2626 2310 2635
rect 2258 2592 2267 2626
rect 2267 2592 2301 2626
rect 2301 2592 2310 2626
rect 2258 2583 2310 2592
rect 2462 2626 2514 2635
rect 2462 2592 2471 2626
rect 2471 2592 2505 2626
rect 2505 2592 2514 2626
rect 2462 2583 2514 2592
rect 2666 2626 2718 2635
rect 2666 2592 2675 2626
rect 2675 2592 2709 2626
rect 2709 2592 2718 2626
rect 2666 2583 2718 2592
rect 2870 2626 2922 2635
rect 2870 2592 2879 2626
rect 2879 2592 2913 2626
rect 2913 2592 2922 2626
rect 2870 2583 2922 2592
rect 3074 2626 3126 2635
rect 3074 2592 3083 2626
rect 3083 2592 3117 2626
rect 3117 2592 3126 2626
rect 3074 2583 3126 2592
rect 3278 2626 3330 2635
rect 3278 2592 3287 2626
rect 3287 2592 3321 2626
rect 3321 2592 3330 2626
rect 3278 2583 3330 2592
rect 3482 2626 3534 2635
rect 3482 2592 3491 2626
rect 3491 2592 3525 2626
rect 3525 2592 3534 2626
rect 3482 2583 3534 2592
rect 3686 2626 3738 2635
rect 3686 2592 3695 2626
rect 3695 2592 3729 2626
rect 3729 2592 3738 2626
rect 3686 2583 3738 2592
rect 3890 2626 3942 2635
rect 3890 2592 3899 2626
rect 3899 2592 3933 2626
rect 3933 2592 3942 2626
rect 3890 2583 3942 2592
rect 4094 2626 4146 2635
rect 4094 2592 4103 2626
rect 4103 2592 4137 2626
rect 4137 2592 4146 2626
rect 4094 2583 4146 2592
rect 4298 2626 4350 2635
rect 4298 2592 4307 2626
rect 4307 2592 4341 2626
rect 4341 2592 4350 2626
rect 4298 2583 4350 2592
rect 4502 2626 4554 2635
rect 4502 2592 4511 2626
rect 4511 2592 4545 2626
rect 4545 2592 4554 2626
rect 4502 2583 4554 2592
rect 4706 2626 4758 2635
rect 4706 2592 4715 2626
rect 4715 2592 4749 2626
rect 4749 2592 4758 2626
rect 4706 2583 4758 2592
rect 4910 2626 4962 2635
rect 4910 2592 4919 2626
rect 4919 2592 4953 2626
rect 4953 2592 4962 2626
rect 4910 2583 4962 2592
rect 5114 2626 5166 2635
rect 5114 2592 5123 2626
rect 5123 2592 5157 2626
rect 5157 2592 5166 2626
rect 5114 2583 5166 2592
rect 5318 2626 5370 2635
rect 5318 2592 5327 2626
rect 5327 2592 5361 2626
rect 5361 2592 5370 2626
rect 5318 2583 5370 2592
rect 5522 2626 5574 2635
rect 5522 2592 5531 2626
rect 5531 2592 5565 2626
rect 5565 2592 5574 2626
rect 5522 2583 5574 2592
rect 5726 2626 5778 2635
rect 5726 2592 5735 2626
rect 5735 2592 5769 2626
rect 5769 2592 5778 2626
rect 5726 2583 5778 2592
rect 5930 2626 5982 2635
rect 5930 2592 5939 2626
rect 5939 2592 5973 2626
rect 5973 2592 5982 2626
rect 5930 2583 5982 2592
rect 6134 2626 6186 2635
rect 6134 2592 6143 2626
rect 6143 2592 6177 2626
rect 6177 2592 6186 2626
rect 6134 2583 6186 2592
rect 6338 2626 6390 2635
rect 6338 2592 6347 2626
rect 6347 2592 6381 2626
rect 6381 2592 6390 2626
rect 6338 2583 6390 2592
rect 6542 2626 6594 2635
rect 6542 2592 6551 2626
rect 6551 2592 6585 2626
rect 6585 2592 6594 2626
rect 6542 2583 6594 2592
rect 6746 2626 6798 2635
rect 6746 2592 6755 2626
rect 6755 2592 6789 2626
rect 6789 2592 6798 2626
rect 6746 2583 6798 2592
rect 6950 2626 7002 2635
rect 6950 2592 6959 2626
rect 6959 2592 6993 2626
rect 6993 2592 7002 2626
rect 6950 2583 7002 2592
rect 7154 2626 7206 2635
rect 7154 2592 7163 2626
rect 7163 2592 7197 2626
rect 7197 2592 7206 2626
rect 7154 2583 7206 2592
rect 7358 2626 7410 2635
rect 7358 2592 7367 2626
rect 7367 2592 7401 2626
rect 7401 2592 7410 2626
rect 7358 2583 7410 2592
rect 7562 2626 7614 2635
rect 7562 2592 7571 2626
rect 7571 2592 7605 2626
rect 7605 2592 7614 2626
rect 7562 2583 7614 2592
rect 7766 2626 7818 2635
rect 7766 2592 7775 2626
rect 7775 2592 7809 2626
rect 7809 2592 7818 2626
rect 7766 2583 7818 2592
rect 7970 2626 8022 2635
rect 7970 2592 7979 2626
rect 7979 2592 8013 2626
rect 8013 2592 8022 2626
rect 7970 2583 8022 2592
rect 8174 2626 8226 2635
rect 8174 2592 8183 2626
rect 8183 2592 8217 2626
rect 8217 2592 8226 2626
rect 8174 2583 8226 2592
rect 8378 2626 8430 2635
rect 8378 2592 8387 2626
rect 8387 2592 8421 2626
rect 8421 2592 8430 2626
rect 8378 2583 8430 2592
rect 8582 2626 8634 2635
rect 8582 2592 8591 2626
rect 8591 2592 8625 2626
rect 8625 2592 8634 2626
rect 8582 2583 8634 2592
rect 8786 2626 8838 2635
rect 8786 2592 8795 2626
rect 8795 2592 8829 2626
rect 8829 2592 8838 2626
rect 8786 2583 8838 2592
rect 8990 2626 9042 2635
rect 8990 2592 8999 2626
rect 8999 2592 9033 2626
rect 9033 2592 9042 2626
rect 8990 2583 9042 2592
rect 9194 2626 9246 2635
rect 9194 2592 9203 2626
rect 9203 2592 9237 2626
rect 9237 2592 9246 2626
rect 9194 2583 9246 2592
rect 9398 2626 9450 2635
rect 9398 2592 9407 2626
rect 9407 2592 9441 2626
rect 9441 2592 9450 2626
rect 9398 2583 9450 2592
rect 9602 2626 9654 2635
rect 9602 2592 9611 2626
rect 9611 2592 9645 2626
rect 9645 2592 9654 2626
rect 9602 2583 9654 2592
rect 9806 2626 9858 2635
rect 9806 2592 9815 2626
rect 9815 2592 9849 2626
rect 9849 2592 9858 2626
rect 9806 2583 9858 2592
rect 10010 2626 10062 2635
rect 10010 2592 10019 2626
rect 10019 2592 10053 2626
rect 10053 2592 10062 2626
rect 10010 2583 10062 2592
rect 10214 2626 10266 2635
rect 10214 2592 10223 2626
rect 10223 2592 10257 2626
rect 10257 2592 10266 2626
rect 10214 2583 10266 2592
rect 10418 2626 10470 2635
rect 10418 2592 10427 2626
rect 10427 2592 10461 2626
rect 10461 2592 10470 2626
rect 10418 2583 10470 2592
rect 10622 2626 10674 2635
rect 10622 2592 10631 2626
rect 10631 2592 10665 2626
rect 10665 2592 10674 2626
rect 10622 2583 10674 2592
rect 10826 2626 10878 2635
rect 10826 2592 10835 2626
rect 10835 2592 10869 2626
rect 10869 2592 10878 2626
rect 10826 2583 10878 2592
rect 11030 2626 11082 2635
rect 11030 2592 11039 2626
rect 11039 2592 11073 2626
rect 11073 2592 11082 2626
rect 11030 2583 11082 2592
rect 11234 2626 11286 2635
rect 11234 2592 11243 2626
rect 11243 2592 11277 2626
rect 11277 2592 11286 2626
rect 11234 2583 11286 2592
rect 11438 2626 11490 2635
rect 11438 2592 11447 2626
rect 11447 2592 11481 2626
rect 11481 2592 11490 2626
rect 11438 2583 11490 2592
rect 11642 2626 11694 2635
rect 11642 2592 11651 2626
rect 11651 2592 11685 2626
rect 11685 2592 11694 2626
rect 11642 2583 11694 2592
rect 11846 2626 11898 2635
rect 11846 2592 11855 2626
rect 11855 2592 11889 2626
rect 11889 2592 11898 2626
rect 11846 2583 11898 2592
rect 12050 2626 12102 2635
rect 12050 2592 12059 2626
rect 12059 2592 12093 2626
rect 12093 2592 12102 2626
rect 12050 2583 12102 2592
rect 12254 2626 12306 2635
rect 12254 2592 12263 2626
rect 12263 2592 12297 2626
rect 12297 2592 12306 2626
rect 12254 2583 12306 2592
rect 12458 2626 12510 2635
rect 12458 2592 12467 2626
rect 12467 2592 12501 2626
rect 12501 2592 12510 2626
rect 12458 2583 12510 2592
rect 12662 2626 12714 2635
rect 12662 2592 12671 2626
rect 12671 2592 12705 2626
rect 12705 2592 12714 2626
rect 12662 2583 12714 2592
rect 12866 2626 12918 2635
rect 12866 2592 12875 2626
rect 12875 2592 12909 2626
rect 12909 2592 12918 2626
rect 12866 2583 12918 2592
rect 13084 2626 13136 2635
rect 13084 2592 13093 2626
rect 13093 2592 13127 2626
rect 13127 2592 13136 2626
rect 13084 2583 13136 2592
rect 7 2472 59 2481
rect 7 2438 16 2472
rect 16 2438 50 2472
rect 50 2438 59 2472
rect 7 2429 59 2438
rect 1639 2472 1691 2481
rect 1639 2438 1648 2472
rect 1648 2438 1682 2472
rect 1682 2438 1691 2472
rect 1639 2429 1691 2438
rect 3271 2472 3323 2481
rect 3271 2438 3280 2472
rect 3280 2438 3314 2472
rect 3314 2438 3323 2472
rect 3271 2429 3323 2438
rect 4903 2472 4955 2481
rect 4903 2438 4912 2472
rect 4912 2438 4946 2472
rect 4946 2438 4955 2472
rect 4903 2429 4955 2438
rect 6535 2472 6587 2481
rect 6535 2438 6544 2472
rect 6544 2438 6578 2472
rect 6578 2438 6587 2472
rect 6535 2429 6587 2438
rect 8167 2472 8219 2481
rect 8167 2438 8176 2472
rect 8176 2438 8210 2472
rect 8210 2438 8219 2472
rect 8167 2429 8219 2438
rect 9799 2472 9851 2481
rect 9799 2438 9808 2472
rect 9808 2438 9842 2472
rect 9842 2438 9851 2472
rect 9799 2429 9851 2438
rect 11431 2472 11483 2481
rect 11431 2438 11440 2472
rect 11440 2438 11474 2472
rect 11474 2438 11483 2472
rect 11431 2429 11483 2438
rect 13063 2472 13115 2481
rect 13063 2438 13072 2472
rect 13072 2438 13106 2472
rect 13106 2438 13115 2472
rect 13063 2429 13115 2438
rect 7 2268 59 2277
rect 7 2234 16 2268
rect 16 2234 50 2268
rect 50 2234 59 2268
rect 7 2225 59 2234
rect 1639 2268 1691 2277
rect 1639 2234 1648 2268
rect 1648 2234 1682 2268
rect 1682 2234 1691 2268
rect 1639 2225 1691 2234
rect 3271 2268 3323 2277
rect 3271 2234 3280 2268
rect 3280 2234 3314 2268
rect 3314 2234 3323 2268
rect 3271 2225 3323 2234
rect 4903 2268 4955 2277
rect 4903 2234 4912 2268
rect 4912 2234 4946 2268
rect 4946 2234 4955 2268
rect 4903 2225 4955 2234
rect 6535 2268 6587 2277
rect 6535 2234 6544 2268
rect 6544 2234 6578 2268
rect 6578 2234 6587 2268
rect 6535 2225 6587 2234
rect 8167 2268 8219 2277
rect 8167 2234 8176 2268
rect 8176 2234 8210 2268
rect 8210 2234 8219 2268
rect 8167 2225 8219 2234
rect 9799 2268 9851 2277
rect 9799 2234 9808 2268
rect 9808 2234 9842 2268
rect 9842 2234 9851 2268
rect 9799 2225 9851 2234
rect 11431 2268 11483 2277
rect 11431 2234 11440 2268
rect 11440 2234 11474 2268
rect 11474 2234 11483 2268
rect 11431 2225 11483 2234
rect 13063 2268 13115 2277
rect 13063 2234 13072 2268
rect 13072 2234 13106 2268
rect 13106 2234 13115 2268
rect 13063 2225 13115 2234
rect 7 2064 59 2073
rect 7 2030 16 2064
rect 16 2030 50 2064
rect 50 2030 59 2064
rect 7 2021 59 2030
rect 1639 2064 1691 2073
rect 1639 2030 1648 2064
rect 1648 2030 1682 2064
rect 1682 2030 1691 2064
rect 1639 2021 1691 2030
rect 3271 2064 3323 2073
rect 3271 2030 3280 2064
rect 3280 2030 3314 2064
rect 3314 2030 3323 2064
rect 3271 2021 3323 2030
rect 4903 2064 4955 2073
rect 4903 2030 4912 2064
rect 4912 2030 4946 2064
rect 4946 2030 4955 2064
rect 4903 2021 4955 2030
rect 6535 2064 6587 2073
rect 6535 2030 6544 2064
rect 6544 2030 6578 2064
rect 6578 2030 6587 2064
rect 6535 2021 6587 2030
rect 8167 2064 8219 2073
rect 8167 2030 8176 2064
rect 8176 2030 8210 2064
rect 8210 2030 8219 2064
rect 8167 2021 8219 2030
rect 9799 2064 9851 2073
rect 9799 2030 9808 2064
rect 9808 2030 9842 2064
rect 9842 2030 9851 2064
rect 9799 2021 9851 2030
rect 11431 2064 11483 2073
rect 11431 2030 11440 2064
rect 11440 2030 11474 2064
rect 11474 2030 11483 2064
rect 11431 2021 11483 2030
rect 13063 2064 13115 2073
rect 13063 2030 13072 2064
rect 13072 2030 13106 2064
rect 13106 2030 13115 2064
rect 13063 2021 13115 2030
rect 7 1860 59 1869
rect 7 1826 16 1860
rect 16 1826 50 1860
rect 50 1826 59 1860
rect 7 1817 59 1826
rect 1639 1860 1691 1869
rect 1639 1826 1648 1860
rect 1648 1826 1682 1860
rect 1682 1826 1691 1860
rect 1639 1817 1691 1826
rect 3271 1860 3323 1869
rect 3271 1826 3280 1860
rect 3280 1826 3314 1860
rect 3314 1826 3323 1860
rect 3271 1817 3323 1826
rect 4903 1860 4955 1869
rect 4903 1826 4912 1860
rect 4912 1826 4946 1860
rect 4946 1826 4955 1860
rect 4903 1817 4955 1826
rect 6535 1860 6587 1869
rect 6535 1826 6544 1860
rect 6544 1826 6578 1860
rect 6578 1826 6587 1860
rect 6535 1817 6587 1826
rect 8167 1860 8219 1869
rect 8167 1826 8176 1860
rect 8176 1826 8210 1860
rect 8210 1826 8219 1860
rect 8167 1817 8219 1826
rect 9799 1860 9851 1869
rect 9799 1826 9808 1860
rect 9808 1826 9842 1860
rect 9842 1826 9851 1860
rect 9799 1817 9851 1826
rect 11431 1860 11483 1869
rect 11431 1826 11440 1860
rect 11440 1826 11474 1860
rect 11474 1826 11483 1860
rect 11431 1817 11483 1826
rect 13063 1860 13115 1869
rect 13063 1826 13072 1860
rect 13072 1826 13106 1860
rect 13106 1826 13115 1860
rect 13063 1817 13115 1826
rect 7 1656 59 1665
rect 7 1622 16 1656
rect 16 1622 50 1656
rect 50 1622 59 1656
rect 7 1613 59 1622
rect 1639 1656 1691 1665
rect 1639 1622 1648 1656
rect 1648 1622 1682 1656
rect 1682 1622 1691 1656
rect 1639 1613 1691 1622
rect 3271 1656 3323 1665
rect 3271 1622 3280 1656
rect 3280 1622 3314 1656
rect 3314 1622 3323 1656
rect 3271 1613 3323 1622
rect 4903 1656 4955 1665
rect 4903 1622 4912 1656
rect 4912 1622 4946 1656
rect 4946 1622 4955 1656
rect 4903 1613 4955 1622
rect 6535 1656 6587 1665
rect 6535 1622 6544 1656
rect 6544 1622 6578 1656
rect 6578 1622 6587 1656
rect 6535 1613 6587 1622
rect 8167 1656 8219 1665
rect 8167 1622 8176 1656
rect 8176 1622 8210 1656
rect 8210 1622 8219 1656
rect 8167 1613 8219 1622
rect 9799 1656 9851 1665
rect 9799 1622 9808 1656
rect 9808 1622 9842 1656
rect 9842 1622 9851 1656
rect 9799 1613 9851 1622
rect 11431 1656 11483 1665
rect 11431 1622 11440 1656
rect 11440 1622 11474 1656
rect 11474 1622 11483 1656
rect 11431 1613 11483 1622
rect 13063 1656 13115 1665
rect 13063 1622 13072 1656
rect 13072 1622 13106 1656
rect 13106 1622 13115 1656
rect 13063 1613 13115 1622
rect 7 1452 59 1461
rect 7 1418 16 1452
rect 16 1418 50 1452
rect 50 1418 59 1452
rect 7 1409 59 1418
rect 1639 1452 1691 1461
rect 1639 1418 1648 1452
rect 1648 1418 1682 1452
rect 1682 1418 1691 1452
rect 1639 1409 1691 1418
rect 3271 1452 3323 1461
rect 3271 1418 3280 1452
rect 3280 1418 3314 1452
rect 3314 1418 3323 1452
rect 3271 1409 3323 1418
rect 4903 1452 4955 1461
rect 4903 1418 4912 1452
rect 4912 1418 4946 1452
rect 4946 1418 4955 1452
rect 4903 1409 4955 1418
rect 6535 1452 6587 1461
rect 6535 1418 6544 1452
rect 6544 1418 6578 1452
rect 6578 1418 6587 1452
rect 6535 1409 6587 1418
rect 8167 1452 8219 1461
rect 8167 1418 8176 1452
rect 8176 1418 8210 1452
rect 8210 1418 8219 1452
rect 8167 1409 8219 1418
rect 9799 1452 9851 1461
rect 9799 1418 9808 1452
rect 9808 1418 9842 1452
rect 9842 1418 9851 1452
rect 9799 1409 9851 1418
rect 11431 1452 11483 1461
rect 11431 1418 11440 1452
rect 11440 1418 11474 1452
rect 11474 1418 11483 1452
rect 11431 1409 11483 1418
rect 13063 1452 13115 1461
rect 13063 1418 13072 1452
rect 13072 1418 13106 1452
rect 13106 1418 13115 1452
rect 13063 1409 13115 1418
rect 7 1248 59 1257
rect 7 1214 16 1248
rect 16 1214 50 1248
rect 50 1214 59 1248
rect 7 1205 59 1214
rect 1639 1248 1691 1257
rect 1639 1214 1648 1248
rect 1648 1214 1682 1248
rect 1682 1214 1691 1248
rect 1639 1205 1691 1214
rect 3271 1248 3323 1257
rect 3271 1214 3280 1248
rect 3280 1214 3314 1248
rect 3314 1214 3323 1248
rect 3271 1205 3323 1214
rect 4903 1248 4955 1257
rect 4903 1214 4912 1248
rect 4912 1214 4946 1248
rect 4946 1214 4955 1248
rect 4903 1205 4955 1214
rect 6535 1248 6587 1257
rect 6535 1214 6544 1248
rect 6544 1214 6578 1248
rect 6578 1214 6587 1248
rect 6535 1205 6587 1214
rect 8167 1248 8219 1257
rect 8167 1214 8176 1248
rect 8176 1214 8210 1248
rect 8210 1214 8219 1248
rect 8167 1205 8219 1214
rect 9799 1248 9851 1257
rect 9799 1214 9808 1248
rect 9808 1214 9842 1248
rect 9842 1214 9851 1248
rect 9799 1205 9851 1214
rect 11431 1248 11483 1257
rect 11431 1214 11440 1248
rect 11440 1214 11474 1248
rect 11474 1214 11483 1248
rect 11431 1205 11483 1214
rect 13063 1248 13115 1257
rect 13063 1214 13072 1248
rect 13072 1214 13106 1248
rect 13106 1214 13115 1248
rect 13063 1205 13115 1214
rect 7 1044 59 1053
rect 7 1010 16 1044
rect 16 1010 50 1044
rect 50 1010 59 1044
rect 7 1001 59 1010
rect 1639 1044 1691 1053
rect 1639 1010 1648 1044
rect 1648 1010 1682 1044
rect 1682 1010 1691 1044
rect 1639 1001 1691 1010
rect 3271 1044 3323 1053
rect 3271 1010 3280 1044
rect 3280 1010 3314 1044
rect 3314 1010 3323 1044
rect 3271 1001 3323 1010
rect 4903 1044 4955 1053
rect 4903 1010 4912 1044
rect 4912 1010 4946 1044
rect 4946 1010 4955 1044
rect 4903 1001 4955 1010
rect 6535 1044 6587 1053
rect 6535 1010 6544 1044
rect 6544 1010 6578 1044
rect 6578 1010 6587 1044
rect 6535 1001 6587 1010
rect 8167 1044 8219 1053
rect 8167 1010 8176 1044
rect 8176 1010 8210 1044
rect 8210 1010 8219 1044
rect 8167 1001 8219 1010
rect 9799 1044 9851 1053
rect 9799 1010 9808 1044
rect 9808 1010 9842 1044
rect 9842 1010 9851 1044
rect 9799 1001 9851 1010
rect 11431 1044 11483 1053
rect 11431 1010 11440 1044
rect 11440 1010 11474 1044
rect 11474 1010 11483 1044
rect 11431 1001 11483 1010
rect 13063 1044 13115 1053
rect 13063 1010 13072 1044
rect 13072 1010 13106 1044
rect 13106 1010 13115 1044
rect 13063 1001 13115 1010
rect 218 890 270 899
rect 218 856 227 890
rect 227 856 261 890
rect 261 856 270 890
rect 218 847 270 856
rect 422 890 474 899
rect 422 856 431 890
rect 431 856 465 890
rect 465 856 474 890
rect 422 847 474 856
rect 626 890 678 899
rect 626 856 635 890
rect 635 856 669 890
rect 669 856 678 890
rect 626 847 678 856
rect 830 890 882 899
rect 830 856 839 890
rect 839 856 873 890
rect 873 856 882 890
rect 830 847 882 856
rect 1034 890 1086 899
rect 1034 856 1043 890
rect 1043 856 1077 890
rect 1077 856 1086 890
rect 1034 847 1086 856
rect 1238 890 1290 899
rect 1238 856 1247 890
rect 1247 856 1281 890
rect 1281 856 1290 890
rect 1238 847 1290 856
rect 1442 890 1494 899
rect 1442 856 1451 890
rect 1451 856 1485 890
rect 1485 856 1494 890
rect 1442 847 1494 856
rect 1646 890 1698 899
rect 1646 856 1655 890
rect 1655 856 1689 890
rect 1689 856 1698 890
rect 1646 847 1698 856
rect 1850 890 1902 899
rect 1850 856 1859 890
rect 1859 856 1893 890
rect 1893 856 1902 890
rect 1850 847 1902 856
rect 2054 890 2106 899
rect 2054 856 2063 890
rect 2063 856 2097 890
rect 2097 856 2106 890
rect 2054 847 2106 856
rect 2258 890 2310 899
rect 2258 856 2267 890
rect 2267 856 2301 890
rect 2301 856 2310 890
rect 2258 847 2310 856
rect 2462 890 2514 899
rect 2462 856 2471 890
rect 2471 856 2505 890
rect 2505 856 2514 890
rect 2462 847 2514 856
rect 2666 890 2718 899
rect 2666 856 2675 890
rect 2675 856 2709 890
rect 2709 856 2718 890
rect 2666 847 2718 856
rect 2870 890 2922 899
rect 2870 856 2879 890
rect 2879 856 2913 890
rect 2913 856 2922 890
rect 2870 847 2922 856
rect 3074 890 3126 899
rect 3074 856 3083 890
rect 3083 856 3117 890
rect 3117 856 3126 890
rect 3074 847 3126 856
rect 3278 890 3330 899
rect 3278 856 3287 890
rect 3287 856 3321 890
rect 3321 856 3330 890
rect 3278 847 3330 856
rect 3482 890 3534 899
rect 3482 856 3491 890
rect 3491 856 3525 890
rect 3525 856 3534 890
rect 3482 847 3534 856
rect 3686 890 3738 899
rect 3686 856 3695 890
rect 3695 856 3729 890
rect 3729 856 3738 890
rect 3686 847 3738 856
rect 3890 890 3942 899
rect 3890 856 3899 890
rect 3899 856 3933 890
rect 3933 856 3942 890
rect 3890 847 3942 856
rect 4094 890 4146 899
rect 4094 856 4103 890
rect 4103 856 4137 890
rect 4137 856 4146 890
rect 4094 847 4146 856
rect 4298 890 4350 899
rect 4298 856 4307 890
rect 4307 856 4341 890
rect 4341 856 4350 890
rect 4298 847 4350 856
rect 4502 890 4554 899
rect 4502 856 4511 890
rect 4511 856 4545 890
rect 4545 856 4554 890
rect 4502 847 4554 856
rect 4706 890 4758 899
rect 4706 856 4715 890
rect 4715 856 4749 890
rect 4749 856 4758 890
rect 4706 847 4758 856
rect 4910 890 4962 899
rect 4910 856 4919 890
rect 4919 856 4953 890
rect 4953 856 4962 890
rect 4910 847 4962 856
rect 5114 890 5166 899
rect 5114 856 5123 890
rect 5123 856 5157 890
rect 5157 856 5166 890
rect 5114 847 5166 856
rect 5318 890 5370 899
rect 5318 856 5327 890
rect 5327 856 5361 890
rect 5361 856 5370 890
rect 5318 847 5370 856
rect 5522 890 5574 899
rect 5522 856 5531 890
rect 5531 856 5565 890
rect 5565 856 5574 890
rect 5522 847 5574 856
rect 5726 890 5778 899
rect 5726 856 5735 890
rect 5735 856 5769 890
rect 5769 856 5778 890
rect 5726 847 5778 856
rect 5930 890 5982 899
rect 5930 856 5939 890
rect 5939 856 5973 890
rect 5973 856 5982 890
rect 5930 847 5982 856
rect 6134 890 6186 899
rect 6134 856 6143 890
rect 6143 856 6177 890
rect 6177 856 6186 890
rect 6134 847 6186 856
rect 6338 890 6390 899
rect 6338 856 6347 890
rect 6347 856 6381 890
rect 6381 856 6390 890
rect 6338 847 6390 856
rect 6542 890 6594 899
rect 6542 856 6551 890
rect 6551 856 6585 890
rect 6585 856 6594 890
rect 6542 847 6594 856
rect 6746 890 6798 899
rect 6746 856 6755 890
rect 6755 856 6789 890
rect 6789 856 6798 890
rect 6746 847 6798 856
rect 6950 890 7002 899
rect 6950 856 6959 890
rect 6959 856 6993 890
rect 6993 856 7002 890
rect 6950 847 7002 856
rect 7154 890 7206 899
rect 7154 856 7163 890
rect 7163 856 7197 890
rect 7197 856 7206 890
rect 7154 847 7206 856
rect 7358 890 7410 899
rect 7358 856 7367 890
rect 7367 856 7401 890
rect 7401 856 7410 890
rect 7358 847 7410 856
rect 7562 890 7614 899
rect 7562 856 7571 890
rect 7571 856 7605 890
rect 7605 856 7614 890
rect 7562 847 7614 856
rect 7766 890 7818 899
rect 7766 856 7775 890
rect 7775 856 7809 890
rect 7809 856 7818 890
rect 7766 847 7818 856
rect 7970 890 8022 899
rect 7970 856 7979 890
rect 7979 856 8013 890
rect 8013 856 8022 890
rect 7970 847 8022 856
rect 8174 890 8226 899
rect 8174 856 8183 890
rect 8183 856 8217 890
rect 8217 856 8226 890
rect 8174 847 8226 856
rect 8378 890 8430 899
rect 8378 856 8387 890
rect 8387 856 8421 890
rect 8421 856 8430 890
rect 8378 847 8430 856
rect 8582 890 8634 899
rect 8582 856 8591 890
rect 8591 856 8625 890
rect 8625 856 8634 890
rect 8582 847 8634 856
rect 8786 890 8838 899
rect 8786 856 8795 890
rect 8795 856 8829 890
rect 8829 856 8838 890
rect 8786 847 8838 856
rect 8990 890 9042 899
rect 8990 856 8999 890
rect 8999 856 9033 890
rect 9033 856 9042 890
rect 8990 847 9042 856
rect 9194 890 9246 899
rect 9194 856 9203 890
rect 9203 856 9237 890
rect 9237 856 9246 890
rect 9194 847 9246 856
rect 9398 890 9450 899
rect 9398 856 9407 890
rect 9407 856 9441 890
rect 9441 856 9450 890
rect 9398 847 9450 856
rect 9602 890 9654 899
rect 9602 856 9611 890
rect 9611 856 9645 890
rect 9645 856 9654 890
rect 9602 847 9654 856
rect 9806 890 9858 899
rect 9806 856 9815 890
rect 9815 856 9849 890
rect 9849 856 9858 890
rect 9806 847 9858 856
rect 10010 890 10062 899
rect 10010 856 10019 890
rect 10019 856 10053 890
rect 10053 856 10062 890
rect 10010 847 10062 856
rect 10214 890 10266 899
rect 10214 856 10223 890
rect 10223 856 10257 890
rect 10257 856 10266 890
rect 10214 847 10266 856
rect 10418 890 10470 899
rect 10418 856 10427 890
rect 10427 856 10461 890
rect 10461 856 10470 890
rect 10418 847 10470 856
rect 10622 890 10674 899
rect 10622 856 10631 890
rect 10631 856 10665 890
rect 10665 856 10674 890
rect 10622 847 10674 856
rect 10826 890 10878 899
rect 10826 856 10835 890
rect 10835 856 10869 890
rect 10869 856 10878 890
rect 10826 847 10878 856
rect 11030 890 11082 899
rect 11030 856 11039 890
rect 11039 856 11073 890
rect 11073 856 11082 890
rect 11030 847 11082 856
rect 11234 890 11286 899
rect 11234 856 11243 890
rect 11243 856 11277 890
rect 11277 856 11286 890
rect 11234 847 11286 856
rect 11438 890 11490 899
rect 11438 856 11447 890
rect 11447 856 11481 890
rect 11481 856 11490 890
rect 11438 847 11490 856
rect 11642 890 11694 899
rect 11642 856 11651 890
rect 11651 856 11685 890
rect 11685 856 11694 890
rect 11642 847 11694 856
rect 11846 890 11898 899
rect 11846 856 11855 890
rect 11855 856 11889 890
rect 11889 856 11898 890
rect 11846 847 11898 856
rect 12050 890 12102 899
rect 12050 856 12059 890
rect 12059 856 12093 890
rect 12093 856 12102 890
rect 12050 847 12102 856
rect 12254 890 12306 899
rect 12254 856 12263 890
rect 12263 856 12297 890
rect 12297 856 12306 890
rect 12254 847 12306 856
rect 12458 890 12510 899
rect 12458 856 12467 890
rect 12467 856 12501 890
rect 12501 856 12510 890
rect 12458 847 12510 856
rect 12662 890 12714 899
rect 12662 856 12671 890
rect 12671 856 12705 890
rect 12705 856 12714 890
rect 12662 847 12714 856
rect 12866 890 12918 899
rect 12866 856 12875 890
rect 12875 856 12909 890
rect 12909 856 12918 890
rect 12866 847 12918 856
rect 13084 890 13136 899
rect 13084 856 13093 890
rect 13093 856 13127 890
rect 13127 856 13136 890
rect 13084 847 13136 856
<< metal2 >>
rect 7 7893 59 7899
rect 1 7846 7 7889
rect 1639 7893 1691 7899
rect 59 7881 65 7889
rect 1633 7881 1639 7889
rect 59 7853 1639 7881
rect 59 7846 65 7853
rect 1633 7846 1639 7853
rect 7 7835 59 7841
rect 3271 7893 3323 7899
rect 1691 7881 1697 7889
rect 3265 7881 3271 7889
rect 1691 7853 3271 7881
rect 1691 7846 1697 7853
rect 3265 7846 3271 7853
rect 1639 7835 1691 7841
rect 4903 7893 4955 7899
rect 3323 7881 3329 7889
rect 4897 7881 4903 7889
rect 3323 7853 4903 7881
rect 3323 7846 3329 7853
rect 4897 7846 4903 7853
rect 3271 7835 3323 7841
rect 6535 7893 6587 7899
rect 4955 7881 4961 7889
rect 6529 7881 6535 7889
rect 4955 7853 6535 7881
rect 4955 7846 4961 7853
rect 6529 7846 6535 7853
rect 4903 7835 4955 7841
rect 8167 7893 8219 7899
rect 6587 7881 6593 7889
rect 8161 7881 8167 7889
rect 6587 7853 8167 7881
rect 6587 7846 6593 7853
rect 8161 7846 8167 7853
rect 6535 7835 6587 7841
rect 9799 7893 9851 7899
rect 8219 7881 8225 7889
rect 9793 7881 9799 7889
rect 8219 7853 9799 7881
rect 8219 7846 8225 7853
rect 9793 7846 9799 7853
rect 8167 7835 8219 7841
rect 11431 7893 11483 7899
rect 9851 7881 9857 7889
rect 11425 7881 11431 7889
rect 9851 7853 11431 7881
rect 9851 7846 9857 7853
rect 11425 7846 11431 7853
rect 9799 7835 9851 7841
rect 13063 7893 13115 7899
rect 11483 7881 11489 7889
rect 13057 7881 13063 7889
rect 11483 7853 13063 7881
rect 11483 7846 11489 7853
rect 13057 7846 13063 7853
rect 11431 7835 11483 7841
rect 13115 7846 13121 7889
rect 13063 7835 13115 7841
rect 7 7689 59 7695
rect 1 7642 7 7685
rect 1639 7689 1691 7695
rect 59 7677 65 7685
rect 1633 7677 1639 7685
rect 59 7649 1639 7677
rect 59 7642 65 7649
rect 1633 7642 1639 7649
rect 7 7631 59 7637
rect 3271 7689 3323 7695
rect 1691 7677 1697 7685
rect 3265 7677 3271 7685
rect 1691 7649 3271 7677
rect 1691 7642 1697 7649
rect 3265 7642 3271 7649
rect 1639 7631 1691 7637
rect 4903 7689 4955 7695
rect 3323 7677 3329 7685
rect 4897 7677 4903 7685
rect 3323 7649 4903 7677
rect 3323 7642 3329 7649
rect 4897 7642 4903 7649
rect 3271 7631 3323 7637
rect 6535 7689 6587 7695
rect 4955 7677 4961 7685
rect 6529 7677 6535 7685
rect 4955 7649 6535 7677
rect 4955 7642 4961 7649
rect 6529 7642 6535 7649
rect 4903 7631 4955 7637
rect 8167 7689 8219 7695
rect 6587 7677 6593 7685
rect 8161 7677 8167 7685
rect 6587 7649 8167 7677
rect 6587 7642 6593 7649
rect 8161 7642 8167 7649
rect 6535 7631 6587 7637
rect 9799 7689 9851 7695
rect 8219 7677 8225 7685
rect 9793 7677 9799 7685
rect 8219 7649 9799 7677
rect 8219 7642 8225 7649
rect 9793 7642 9799 7649
rect 8167 7631 8219 7637
rect 11431 7689 11483 7695
rect 9851 7677 9857 7685
rect 11425 7677 11431 7685
rect 9851 7649 11431 7677
rect 9851 7642 9857 7649
rect 11425 7642 11431 7649
rect 9799 7631 9851 7637
rect 13063 7689 13115 7695
rect 11483 7677 11489 7685
rect 13057 7677 13063 7685
rect 11483 7649 13063 7677
rect 11483 7642 11489 7649
rect 13057 7642 13063 7649
rect 11431 7631 11483 7637
rect 13115 7642 13121 7685
rect 13063 7631 13115 7637
rect 7 7485 59 7491
rect 1 7438 7 7481
rect 1639 7485 1691 7491
rect 59 7473 65 7481
rect 1633 7473 1639 7481
rect 59 7445 1639 7473
rect 59 7438 65 7445
rect 1633 7438 1639 7445
rect 7 7427 59 7433
rect 3271 7485 3323 7491
rect 1691 7473 1697 7481
rect 3265 7473 3271 7481
rect 1691 7445 3271 7473
rect 1691 7438 1697 7445
rect 3265 7438 3271 7445
rect 1639 7427 1691 7433
rect 4903 7485 4955 7491
rect 3323 7473 3329 7481
rect 4897 7473 4903 7481
rect 3323 7445 4903 7473
rect 3323 7438 3329 7445
rect 4897 7438 4903 7445
rect 3271 7427 3323 7433
rect 6535 7485 6587 7491
rect 4955 7473 4961 7481
rect 6529 7473 6535 7481
rect 4955 7445 6535 7473
rect 4955 7438 4961 7445
rect 6529 7438 6535 7445
rect 4903 7427 4955 7433
rect 8167 7485 8219 7491
rect 6587 7473 6593 7481
rect 8161 7473 8167 7481
rect 6587 7445 8167 7473
rect 6587 7438 6593 7445
rect 8161 7438 8167 7445
rect 6535 7427 6587 7433
rect 9799 7485 9851 7491
rect 8219 7473 8225 7481
rect 9793 7473 9799 7481
rect 8219 7445 9799 7473
rect 8219 7438 8225 7445
rect 9793 7438 9799 7445
rect 8167 7427 8219 7433
rect 11431 7485 11483 7491
rect 9851 7473 9857 7481
rect 11425 7473 11431 7481
rect 9851 7445 11431 7473
rect 9851 7438 9857 7445
rect 11425 7438 11431 7445
rect 9799 7427 9851 7433
rect 13063 7485 13115 7491
rect 11483 7473 11489 7481
rect 13057 7473 13063 7481
rect 11483 7445 13063 7473
rect 11483 7438 11489 7445
rect 13057 7438 13063 7445
rect 11431 7427 11483 7433
rect 13115 7438 13121 7481
rect 13063 7427 13115 7433
rect 7 7281 59 7287
rect 1 7234 7 7277
rect 1639 7281 1691 7287
rect 59 7269 65 7277
rect 1633 7269 1639 7277
rect 59 7241 1639 7269
rect 59 7234 65 7241
rect 1633 7234 1639 7241
rect 7 7223 59 7229
rect 3271 7281 3323 7287
rect 1691 7269 1697 7277
rect 3265 7269 3271 7277
rect 1691 7241 3271 7269
rect 1691 7234 1697 7241
rect 3265 7234 3271 7241
rect 1639 7223 1691 7229
rect 4903 7281 4955 7287
rect 3323 7269 3329 7277
rect 4897 7269 4903 7277
rect 3323 7241 4903 7269
rect 3323 7234 3329 7241
rect 4897 7234 4903 7241
rect 3271 7223 3323 7229
rect 6535 7281 6587 7287
rect 4955 7269 4961 7277
rect 6529 7269 6535 7277
rect 4955 7241 6535 7269
rect 4955 7234 4961 7241
rect 6529 7234 6535 7241
rect 4903 7223 4955 7229
rect 8167 7281 8219 7287
rect 6587 7269 6593 7277
rect 8161 7269 8167 7277
rect 6587 7241 8167 7269
rect 6587 7234 6593 7241
rect 8161 7234 8167 7241
rect 6535 7223 6587 7229
rect 9799 7281 9851 7287
rect 8219 7269 8225 7277
rect 9793 7269 9799 7277
rect 8219 7241 9799 7269
rect 8219 7234 8225 7241
rect 9793 7234 9799 7241
rect 8167 7223 8219 7229
rect 11431 7281 11483 7287
rect 9851 7269 9857 7277
rect 11425 7269 11431 7277
rect 9851 7241 11431 7269
rect 9851 7234 9857 7241
rect 11425 7234 11431 7241
rect 9799 7223 9851 7229
rect 13063 7281 13115 7287
rect 11483 7269 11489 7277
rect 13057 7269 13063 7277
rect 11483 7241 13063 7269
rect 11483 7234 11489 7241
rect 13057 7234 13063 7241
rect 11431 7223 11483 7229
rect 13115 7234 13121 7277
rect 13063 7223 13115 7229
rect 7 7077 59 7083
rect 1 7030 7 7073
rect 1639 7077 1691 7083
rect 59 7065 65 7073
rect 1633 7065 1639 7073
rect 59 7037 1639 7065
rect 59 7030 65 7037
rect 1633 7030 1639 7037
rect 7 7019 59 7025
rect 3271 7077 3323 7083
rect 1691 7065 1697 7073
rect 3265 7065 3271 7073
rect 1691 7037 3271 7065
rect 1691 7030 1697 7037
rect 3265 7030 3271 7037
rect 1639 7019 1691 7025
rect 4903 7077 4955 7083
rect 3323 7065 3329 7073
rect 4897 7065 4903 7073
rect 3323 7037 4903 7065
rect 3323 7030 3329 7037
rect 4897 7030 4903 7037
rect 3271 7019 3323 7025
rect 6535 7077 6587 7083
rect 4955 7065 4961 7073
rect 6529 7065 6535 7073
rect 4955 7037 6535 7065
rect 4955 7030 4961 7037
rect 6529 7030 6535 7037
rect 4903 7019 4955 7025
rect 8167 7077 8219 7083
rect 6587 7065 6593 7073
rect 8161 7065 8167 7073
rect 6587 7037 8167 7065
rect 6587 7030 6593 7037
rect 8161 7030 8167 7037
rect 6535 7019 6587 7025
rect 9799 7077 9851 7083
rect 8219 7065 8225 7073
rect 9793 7065 9799 7073
rect 8219 7037 9799 7065
rect 8219 7030 8225 7037
rect 9793 7030 9799 7037
rect 8167 7019 8219 7025
rect 11431 7077 11483 7083
rect 9851 7065 9857 7073
rect 11425 7065 11431 7073
rect 9851 7037 11431 7065
rect 9851 7030 9857 7037
rect 11425 7030 11431 7037
rect 9799 7019 9851 7025
rect 13063 7077 13115 7083
rect 11483 7065 11489 7073
rect 13057 7065 13063 7073
rect 11483 7037 13063 7065
rect 11483 7030 11489 7037
rect 13057 7030 13063 7037
rect 11431 7019 11483 7025
rect 13115 7030 13121 7073
rect 13063 7019 13115 7025
rect 7 6873 59 6879
rect 1 6826 7 6869
rect 1639 6873 1691 6879
rect 59 6861 65 6869
rect 1633 6861 1639 6869
rect 59 6833 1639 6861
rect 59 6826 65 6833
rect 1633 6826 1639 6833
rect 7 6815 59 6821
rect 3271 6873 3323 6879
rect 1691 6861 1697 6869
rect 3265 6861 3271 6869
rect 1691 6833 3271 6861
rect 1691 6826 1697 6833
rect 3265 6826 3271 6833
rect 1639 6815 1691 6821
rect 4903 6873 4955 6879
rect 3323 6861 3329 6869
rect 4897 6861 4903 6869
rect 3323 6833 4903 6861
rect 3323 6826 3329 6833
rect 4897 6826 4903 6833
rect 3271 6815 3323 6821
rect 6535 6873 6587 6879
rect 4955 6861 4961 6869
rect 6529 6861 6535 6869
rect 4955 6833 6535 6861
rect 4955 6826 4961 6833
rect 6529 6826 6535 6833
rect 4903 6815 4955 6821
rect 8167 6873 8219 6879
rect 6587 6861 6593 6869
rect 8161 6861 8167 6869
rect 6587 6833 8167 6861
rect 6587 6826 6593 6833
rect 8161 6826 8167 6833
rect 6535 6815 6587 6821
rect 9799 6873 9851 6879
rect 8219 6861 8225 6869
rect 9793 6861 9799 6869
rect 8219 6833 9799 6861
rect 8219 6826 8225 6833
rect 9793 6826 9799 6833
rect 8167 6815 8219 6821
rect 11431 6873 11483 6879
rect 9851 6861 9857 6869
rect 11425 6861 11431 6869
rect 9851 6833 11431 6861
rect 9851 6826 9857 6833
rect 11425 6826 11431 6833
rect 9799 6815 9851 6821
rect 13063 6873 13115 6879
rect 11483 6861 11489 6869
rect 13057 6861 13063 6869
rect 11483 6833 13063 6861
rect 11483 6826 11489 6833
rect 13057 6826 13063 6833
rect 11431 6815 11483 6821
rect 13115 6826 13121 6869
rect 13063 6815 13115 6821
rect 7 6669 59 6675
rect 1 6622 7 6665
rect 1639 6669 1691 6675
rect 59 6657 65 6665
rect 1633 6657 1639 6665
rect 59 6629 1639 6657
rect 59 6622 65 6629
rect 1633 6622 1639 6629
rect 7 6611 59 6617
rect 3271 6669 3323 6675
rect 1691 6657 1697 6665
rect 3265 6657 3271 6665
rect 1691 6629 3271 6657
rect 1691 6622 1697 6629
rect 3265 6622 3271 6629
rect 1639 6611 1691 6617
rect 4903 6669 4955 6675
rect 3323 6657 3329 6665
rect 4897 6657 4903 6665
rect 3323 6629 4903 6657
rect 3323 6622 3329 6629
rect 4897 6622 4903 6629
rect 3271 6611 3323 6617
rect 6535 6669 6587 6675
rect 4955 6657 4961 6665
rect 6529 6657 6535 6665
rect 4955 6629 6535 6657
rect 4955 6622 4961 6629
rect 6529 6622 6535 6629
rect 4903 6611 4955 6617
rect 8167 6669 8219 6675
rect 6587 6657 6593 6665
rect 8161 6657 8167 6665
rect 6587 6629 8167 6657
rect 6587 6622 6593 6629
rect 8161 6622 8167 6629
rect 6535 6611 6587 6617
rect 9799 6669 9851 6675
rect 8219 6657 8225 6665
rect 9793 6657 9799 6665
rect 8219 6629 9799 6657
rect 8219 6622 8225 6629
rect 9793 6622 9799 6629
rect 8167 6611 8219 6617
rect 11431 6669 11483 6675
rect 9851 6657 9857 6665
rect 11425 6657 11431 6665
rect 9851 6629 11431 6657
rect 9851 6622 9857 6629
rect 11425 6622 11431 6629
rect 9799 6611 9851 6617
rect 13063 6669 13115 6675
rect 11483 6657 11489 6665
rect 13057 6657 13063 6665
rect 11483 6629 13063 6657
rect 11483 6622 11489 6629
rect 13057 6622 13063 6629
rect 11431 6611 11483 6617
rect 13115 6622 13121 6665
rect 13063 6611 13115 6617
rect 7 6465 59 6471
rect 1 6418 7 6461
rect 1639 6465 1691 6471
rect 59 6453 65 6461
rect 1633 6453 1639 6461
rect 59 6425 1639 6453
rect 59 6418 65 6425
rect 1633 6418 1639 6425
rect 7 6407 59 6413
rect 3271 6465 3323 6471
rect 1691 6453 1697 6461
rect 3265 6453 3271 6461
rect 1691 6425 3271 6453
rect 1691 6418 1697 6425
rect 3265 6418 3271 6425
rect 1639 6407 1691 6413
rect 4903 6465 4955 6471
rect 3323 6453 3329 6461
rect 4897 6453 4903 6461
rect 3323 6425 4903 6453
rect 3323 6418 3329 6425
rect 4897 6418 4903 6425
rect 3271 6407 3323 6413
rect 6535 6465 6587 6471
rect 4955 6453 4961 6461
rect 6529 6453 6535 6461
rect 4955 6425 6535 6453
rect 4955 6418 4961 6425
rect 6529 6418 6535 6425
rect 4903 6407 4955 6413
rect 8167 6465 8219 6471
rect 6587 6453 6593 6461
rect 8161 6453 8167 6461
rect 6587 6425 8167 6453
rect 6587 6418 6593 6425
rect 8161 6418 8167 6425
rect 6535 6407 6587 6413
rect 9799 6465 9851 6471
rect 8219 6453 8225 6461
rect 9793 6453 9799 6461
rect 8219 6425 9799 6453
rect 8219 6418 8225 6425
rect 9793 6418 9799 6425
rect 8167 6407 8219 6413
rect 11431 6465 11483 6471
rect 9851 6453 9857 6461
rect 11425 6453 11431 6461
rect 9851 6425 11431 6453
rect 9851 6418 9857 6425
rect 11425 6418 11431 6425
rect 9799 6407 9851 6413
rect 13063 6465 13115 6471
rect 11483 6453 11489 6461
rect 13057 6453 13063 6461
rect 11483 6425 13063 6453
rect 11483 6418 11489 6425
rect 13057 6418 13063 6425
rect 11431 6407 11483 6413
rect 13115 6418 13121 6461
rect 13063 6407 13115 6413
rect 7 6261 59 6267
rect 1 6214 7 6257
rect 1639 6261 1691 6267
rect 59 6249 65 6257
rect 1633 6249 1639 6257
rect 59 6221 1639 6249
rect 59 6214 65 6221
rect 1633 6214 1639 6221
rect 7 6203 59 6209
rect 3271 6261 3323 6267
rect 1691 6249 1697 6257
rect 3265 6249 3271 6257
rect 1691 6221 3271 6249
rect 1691 6214 1697 6221
rect 3265 6214 3271 6221
rect 1639 6203 1691 6209
rect 4903 6261 4955 6267
rect 3323 6249 3329 6257
rect 4897 6249 4903 6257
rect 3323 6221 4903 6249
rect 3323 6214 3329 6221
rect 4897 6214 4903 6221
rect 3271 6203 3323 6209
rect 6535 6261 6587 6267
rect 4955 6249 4961 6257
rect 6529 6249 6535 6257
rect 4955 6221 6535 6249
rect 4955 6214 4961 6221
rect 6529 6214 6535 6221
rect 4903 6203 4955 6209
rect 8167 6261 8219 6267
rect 6587 6249 6593 6257
rect 8161 6249 8167 6257
rect 6587 6221 8167 6249
rect 6587 6214 6593 6221
rect 8161 6214 8167 6221
rect 6535 6203 6587 6209
rect 9799 6261 9851 6267
rect 8219 6249 8225 6257
rect 9793 6249 9799 6257
rect 8219 6221 9799 6249
rect 8219 6214 8225 6221
rect 9793 6214 9799 6221
rect 8167 6203 8219 6209
rect 11431 6261 11483 6267
rect 9851 6249 9857 6257
rect 11425 6249 11431 6257
rect 9851 6221 11431 6249
rect 9851 6214 9857 6221
rect 11425 6214 11431 6221
rect 9799 6203 9851 6209
rect 13063 6261 13115 6267
rect 11483 6249 11489 6257
rect 13057 6249 13063 6257
rect 11483 6221 13063 6249
rect 11483 6214 11489 6221
rect 13057 6214 13063 6221
rect 11431 6203 11483 6209
rect 13115 6214 13121 6257
rect 13063 6203 13115 6209
rect 212 6055 218 6107
rect 270 6095 276 6107
rect 416 6095 422 6107
rect 270 6067 422 6095
rect 270 6055 276 6067
rect 416 6055 422 6067
rect 474 6095 480 6107
rect 620 6095 626 6107
rect 474 6067 626 6095
rect 474 6055 480 6067
rect 620 6055 626 6067
rect 678 6095 684 6107
rect 824 6095 830 6107
rect 678 6067 830 6095
rect 678 6055 684 6067
rect 824 6055 830 6067
rect 882 6095 888 6107
rect 1028 6095 1034 6107
rect 882 6067 1034 6095
rect 882 6055 888 6067
rect 1028 6055 1034 6067
rect 1086 6095 1092 6107
rect 1232 6095 1238 6107
rect 1086 6067 1238 6095
rect 1086 6055 1092 6067
rect 1232 6055 1238 6067
rect 1290 6095 1296 6107
rect 1436 6095 1442 6107
rect 1290 6067 1442 6095
rect 1290 6055 1296 6067
rect 1436 6055 1442 6067
rect 1494 6095 1500 6107
rect 1640 6095 1646 6107
rect 1494 6067 1646 6095
rect 1494 6055 1500 6067
rect 1640 6055 1646 6067
rect 1698 6095 1704 6107
rect 1844 6095 1850 6107
rect 1698 6067 1850 6095
rect 1698 6055 1704 6067
rect 1844 6055 1850 6067
rect 1902 6095 1908 6107
rect 2048 6095 2054 6107
rect 1902 6067 2054 6095
rect 1902 6055 1908 6067
rect 2048 6055 2054 6067
rect 2106 6095 2112 6107
rect 2252 6095 2258 6107
rect 2106 6067 2258 6095
rect 2106 6055 2112 6067
rect 2252 6055 2258 6067
rect 2310 6095 2316 6107
rect 2456 6095 2462 6107
rect 2310 6067 2462 6095
rect 2310 6055 2316 6067
rect 2456 6055 2462 6067
rect 2514 6095 2520 6107
rect 2660 6095 2666 6107
rect 2514 6067 2666 6095
rect 2514 6055 2520 6067
rect 2660 6055 2666 6067
rect 2718 6095 2724 6107
rect 2864 6095 2870 6107
rect 2718 6067 2870 6095
rect 2718 6055 2724 6067
rect 2864 6055 2870 6067
rect 2922 6095 2928 6107
rect 3068 6095 3074 6107
rect 2922 6067 3074 6095
rect 2922 6055 2928 6067
rect 3068 6055 3074 6067
rect 3126 6095 3132 6107
rect 3272 6095 3278 6107
rect 3126 6067 3278 6095
rect 3126 6055 3132 6067
rect 3272 6055 3278 6067
rect 3330 6095 3336 6107
rect 3476 6095 3482 6107
rect 3330 6067 3482 6095
rect 3330 6055 3336 6067
rect 3476 6055 3482 6067
rect 3534 6095 3540 6107
rect 3680 6095 3686 6107
rect 3534 6067 3686 6095
rect 3534 6055 3540 6067
rect 3680 6055 3686 6067
rect 3738 6095 3744 6107
rect 3884 6095 3890 6107
rect 3738 6067 3890 6095
rect 3738 6055 3744 6067
rect 3884 6055 3890 6067
rect 3942 6095 3948 6107
rect 4088 6095 4094 6107
rect 3942 6067 4094 6095
rect 3942 6055 3948 6067
rect 4088 6055 4094 6067
rect 4146 6095 4152 6107
rect 4292 6095 4298 6107
rect 4146 6067 4298 6095
rect 4146 6055 4152 6067
rect 4292 6055 4298 6067
rect 4350 6095 4356 6107
rect 4496 6095 4502 6107
rect 4350 6067 4502 6095
rect 4350 6055 4356 6067
rect 4496 6055 4502 6067
rect 4554 6095 4560 6107
rect 4700 6095 4706 6107
rect 4554 6067 4706 6095
rect 4554 6055 4560 6067
rect 4700 6055 4706 6067
rect 4758 6095 4764 6107
rect 4904 6095 4910 6107
rect 4758 6067 4910 6095
rect 4758 6055 4764 6067
rect 4904 6055 4910 6067
rect 4962 6095 4968 6107
rect 5108 6095 5114 6107
rect 4962 6067 5114 6095
rect 4962 6055 4968 6067
rect 5108 6055 5114 6067
rect 5166 6095 5172 6107
rect 5312 6095 5318 6107
rect 5166 6067 5318 6095
rect 5166 6055 5172 6067
rect 5312 6055 5318 6067
rect 5370 6095 5376 6107
rect 5516 6095 5522 6107
rect 5370 6067 5522 6095
rect 5370 6055 5376 6067
rect 5516 6055 5522 6067
rect 5574 6095 5580 6107
rect 5720 6095 5726 6107
rect 5574 6067 5726 6095
rect 5574 6055 5580 6067
rect 5720 6055 5726 6067
rect 5778 6095 5784 6107
rect 5924 6095 5930 6107
rect 5778 6067 5930 6095
rect 5778 6055 5784 6067
rect 5924 6055 5930 6067
rect 5982 6095 5988 6107
rect 6128 6095 6134 6107
rect 5982 6067 6134 6095
rect 5982 6055 5988 6067
rect 6128 6055 6134 6067
rect 6186 6095 6192 6107
rect 6332 6095 6338 6107
rect 6186 6067 6338 6095
rect 6186 6055 6192 6067
rect 6332 6055 6338 6067
rect 6390 6095 6396 6107
rect 6536 6095 6542 6107
rect 6390 6067 6542 6095
rect 6390 6055 6396 6067
rect 6536 6055 6542 6067
rect 6594 6095 6600 6107
rect 6740 6095 6746 6107
rect 6594 6067 6746 6095
rect 6594 6055 6600 6067
rect 6740 6055 6746 6067
rect 6798 6095 6804 6107
rect 6944 6095 6950 6107
rect 6798 6067 6950 6095
rect 6798 6055 6804 6067
rect 6944 6055 6950 6067
rect 7002 6095 7008 6107
rect 7148 6095 7154 6107
rect 7002 6067 7154 6095
rect 7002 6055 7008 6067
rect 7148 6055 7154 6067
rect 7206 6095 7212 6107
rect 7352 6095 7358 6107
rect 7206 6067 7358 6095
rect 7206 6055 7212 6067
rect 7352 6055 7358 6067
rect 7410 6095 7416 6107
rect 7556 6095 7562 6107
rect 7410 6067 7562 6095
rect 7410 6055 7416 6067
rect 7556 6055 7562 6067
rect 7614 6095 7620 6107
rect 7760 6095 7766 6107
rect 7614 6067 7766 6095
rect 7614 6055 7620 6067
rect 7760 6055 7766 6067
rect 7818 6095 7824 6107
rect 7964 6095 7970 6107
rect 7818 6067 7970 6095
rect 7818 6055 7824 6067
rect 7964 6055 7970 6067
rect 8022 6095 8028 6107
rect 8168 6095 8174 6107
rect 8022 6067 8174 6095
rect 8022 6055 8028 6067
rect 8168 6055 8174 6067
rect 8226 6095 8232 6107
rect 8372 6095 8378 6107
rect 8226 6067 8378 6095
rect 8226 6055 8232 6067
rect 8372 6055 8378 6067
rect 8430 6095 8436 6107
rect 8576 6095 8582 6107
rect 8430 6067 8582 6095
rect 8430 6055 8436 6067
rect 8576 6055 8582 6067
rect 8634 6095 8640 6107
rect 8780 6095 8786 6107
rect 8634 6067 8786 6095
rect 8634 6055 8640 6067
rect 8780 6055 8786 6067
rect 8838 6095 8844 6107
rect 8984 6095 8990 6107
rect 8838 6067 8990 6095
rect 8838 6055 8844 6067
rect 8984 6055 8990 6067
rect 9042 6095 9048 6107
rect 9188 6095 9194 6107
rect 9042 6067 9194 6095
rect 9042 6055 9048 6067
rect 9188 6055 9194 6067
rect 9246 6095 9252 6107
rect 9392 6095 9398 6107
rect 9246 6067 9398 6095
rect 9246 6055 9252 6067
rect 9392 6055 9398 6067
rect 9450 6095 9456 6107
rect 9596 6095 9602 6107
rect 9450 6067 9602 6095
rect 9450 6055 9456 6067
rect 9596 6055 9602 6067
rect 9654 6095 9660 6107
rect 9800 6095 9806 6107
rect 9654 6067 9806 6095
rect 9654 6055 9660 6067
rect 9800 6055 9806 6067
rect 9858 6095 9864 6107
rect 10004 6095 10010 6107
rect 9858 6067 10010 6095
rect 9858 6055 9864 6067
rect 10004 6055 10010 6067
rect 10062 6095 10068 6107
rect 10208 6095 10214 6107
rect 10062 6067 10214 6095
rect 10062 6055 10068 6067
rect 10208 6055 10214 6067
rect 10266 6095 10272 6107
rect 10412 6095 10418 6107
rect 10266 6067 10418 6095
rect 10266 6055 10272 6067
rect 10412 6055 10418 6067
rect 10470 6095 10476 6107
rect 10616 6095 10622 6107
rect 10470 6067 10622 6095
rect 10470 6055 10476 6067
rect 10616 6055 10622 6067
rect 10674 6095 10680 6107
rect 10820 6095 10826 6107
rect 10674 6067 10826 6095
rect 10674 6055 10680 6067
rect 10820 6055 10826 6067
rect 10878 6095 10884 6107
rect 11024 6095 11030 6107
rect 10878 6067 11030 6095
rect 10878 6055 10884 6067
rect 11024 6055 11030 6067
rect 11082 6095 11088 6107
rect 11228 6095 11234 6107
rect 11082 6067 11234 6095
rect 11082 6055 11088 6067
rect 11228 6055 11234 6067
rect 11286 6095 11292 6107
rect 11432 6095 11438 6107
rect 11286 6067 11438 6095
rect 11286 6055 11292 6067
rect 11432 6055 11438 6067
rect 11490 6095 11496 6107
rect 11636 6095 11642 6107
rect 11490 6067 11642 6095
rect 11490 6055 11496 6067
rect 11636 6055 11642 6067
rect 11694 6095 11700 6107
rect 11840 6095 11846 6107
rect 11694 6067 11846 6095
rect 11694 6055 11700 6067
rect 11840 6055 11846 6067
rect 11898 6095 11904 6107
rect 12044 6095 12050 6107
rect 11898 6067 12050 6095
rect 11898 6055 11904 6067
rect 12044 6055 12050 6067
rect 12102 6095 12108 6107
rect 12248 6095 12254 6107
rect 12102 6067 12254 6095
rect 12102 6055 12108 6067
rect 12248 6055 12254 6067
rect 12306 6095 12312 6107
rect 12452 6095 12458 6107
rect 12306 6067 12458 6095
rect 12306 6055 12312 6067
rect 12452 6055 12458 6067
rect 12510 6095 12516 6107
rect 12656 6095 12662 6107
rect 12510 6067 12662 6095
rect 12510 6055 12516 6067
rect 12656 6055 12662 6067
rect 12714 6095 12720 6107
rect 12860 6095 12866 6107
rect 12714 6067 12866 6095
rect 12714 6055 12720 6067
rect 12860 6055 12866 6067
rect 12918 6095 12924 6107
rect 13078 6095 13084 6107
rect 12918 6067 13084 6095
rect 12918 6055 12924 6067
rect 13078 6055 13084 6067
rect 13136 6055 13142 6107
rect 7 5953 59 5959
rect 1 5906 7 5949
rect 1639 5953 1691 5959
rect 59 5941 65 5949
rect 1633 5941 1639 5949
rect 59 5913 1639 5941
rect 59 5906 65 5913
rect 1633 5906 1639 5913
rect 7 5895 59 5901
rect 3271 5953 3323 5959
rect 1691 5941 1697 5949
rect 3265 5941 3271 5949
rect 1691 5913 3271 5941
rect 1691 5906 1697 5913
rect 3265 5906 3271 5913
rect 1639 5895 1691 5901
rect 4903 5953 4955 5959
rect 3323 5941 3329 5949
rect 4897 5941 4903 5949
rect 3323 5913 4903 5941
rect 3323 5906 3329 5913
rect 4897 5906 4903 5913
rect 3271 5895 3323 5901
rect 6535 5953 6587 5959
rect 4955 5941 4961 5949
rect 6529 5941 6535 5949
rect 4955 5913 6535 5941
rect 4955 5906 4961 5913
rect 6529 5906 6535 5913
rect 4903 5895 4955 5901
rect 8167 5953 8219 5959
rect 6587 5941 6593 5949
rect 8161 5941 8167 5949
rect 6587 5913 8167 5941
rect 6587 5906 6593 5913
rect 8161 5906 8167 5913
rect 6535 5895 6587 5901
rect 9799 5953 9851 5959
rect 8219 5941 8225 5949
rect 9793 5941 9799 5949
rect 8219 5913 9799 5941
rect 8219 5906 8225 5913
rect 9793 5906 9799 5913
rect 8167 5895 8219 5901
rect 11431 5953 11483 5959
rect 9851 5941 9857 5949
rect 11425 5941 11431 5949
rect 9851 5913 11431 5941
rect 9851 5906 9857 5913
rect 11425 5906 11431 5913
rect 9799 5895 9851 5901
rect 13063 5953 13115 5959
rect 11483 5941 11489 5949
rect 13057 5941 13063 5949
rect 11483 5913 13063 5941
rect 11483 5906 11489 5913
rect 13057 5906 13063 5913
rect 11431 5895 11483 5901
rect 13115 5906 13121 5949
rect 13063 5895 13115 5901
rect 7 5749 59 5755
rect 1 5702 7 5745
rect 1639 5749 1691 5755
rect 59 5737 65 5745
rect 1633 5737 1639 5745
rect 59 5709 1639 5737
rect 59 5702 65 5709
rect 1633 5702 1639 5709
rect 7 5691 59 5697
rect 3271 5749 3323 5755
rect 1691 5737 1697 5745
rect 3265 5737 3271 5745
rect 1691 5709 3271 5737
rect 1691 5702 1697 5709
rect 3265 5702 3271 5709
rect 1639 5691 1691 5697
rect 4903 5749 4955 5755
rect 3323 5737 3329 5745
rect 4897 5737 4903 5745
rect 3323 5709 4903 5737
rect 3323 5702 3329 5709
rect 4897 5702 4903 5709
rect 3271 5691 3323 5697
rect 6535 5749 6587 5755
rect 4955 5737 4961 5745
rect 6529 5737 6535 5745
rect 4955 5709 6535 5737
rect 4955 5702 4961 5709
rect 6529 5702 6535 5709
rect 4903 5691 4955 5697
rect 8167 5749 8219 5755
rect 6587 5737 6593 5745
rect 8161 5737 8167 5745
rect 6587 5709 8167 5737
rect 6587 5702 6593 5709
rect 8161 5702 8167 5709
rect 6535 5691 6587 5697
rect 9799 5749 9851 5755
rect 8219 5737 8225 5745
rect 9793 5737 9799 5745
rect 8219 5709 9799 5737
rect 8219 5702 8225 5709
rect 9793 5702 9799 5709
rect 8167 5691 8219 5697
rect 11431 5749 11483 5755
rect 9851 5737 9857 5745
rect 11425 5737 11431 5745
rect 9851 5709 11431 5737
rect 9851 5702 9857 5709
rect 11425 5702 11431 5709
rect 9799 5691 9851 5697
rect 13063 5749 13115 5755
rect 11483 5737 11489 5745
rect 13057 5737 13063 5745
rect 11483 5709 13063 5737
rect 11483 5702 11489 5709
rect 13057 5702 13063 5709
rect 11431 5691 11483 5697
rect 13115 5702 13121 5745
rect 13063 5691 13115 5697
rect 7 5545 59 5551
rect 1 5498 7 5541
rect 1639 5545 1691 5551
rect 59 5533 65 5541
rect 1633 5533 1639 5541
rect 59 5505 1639 5533
rect 59 5498 65 5505
rect 1633 5498 1639 5505
rect 7 5487 59 5493
rect 3271 5545 3323 5551
rect 1691 5533 1697 5541
rect 3265 5533 3271 5541
rect 1691 5505 3271 5533
rect 1691 5498 1697 5505
rect 3265 5498 3271 5505
rect 1639 5487 1691 5493
rect 4903 5545 4955 5551
rect 3323 5533 3329 5541
rect 4897 5533 4903 5541
rect 3323 5505 4903 5533
rect 3323 5498 3329 5505
rect 4897 5498 4903 5505
rect 3271 5487 3323 5493
rect 6535 5545 6587 5551
rect 4955 5533 4961 5541
rect 6529 5533 6535 5541
rect 4955 5505 6535 5533
rect 4955 5498 4961 5505
rect 6529 5498 6535 5505
rect 4903 5487 4955 5493
rect 8167 5545 8219 5551
rect 6587 5533 6593 5541
rect 8161 5533 8167 5541
rect 6587 5505 8167 5533
rect 6587 5498 6593 5505
rect 8161 5498 8167 5505
rect 6535 5487 6587 5493
rect 9799 5545 9851 5551
rect 8219 5533 8225 5541
rect 9793 5533 9799 5541
rect 8219 5505 9799 5533
rect 8219 5498 8225 5505
rect 9793 5498 9799 5505
rect 8167 5487 8219 5493
rect 11431 5545 11483 5551
rect 9851 5533 9857 5541
rect 11425 5533 11431 5541
rect 9851 5505 11431 5533
rect 9851 5498 9857 5505
rect 11425 5498 11431 5505
rect 9799 5487 9851 5493
rect 13063 5545 13115 5551
rect 11483 5533 11489 5541
rect 13057 5533 13063 5541
rect 11483 5505 13063 5533
rect 11483 5498 11489 5505
rect 13057 5498 13063 5505
rect 11431 5487 11483 5493
rect 13115 5498 13121 5541
rect 13063 5487 13115 5493
rect 7 5341 59 5347
rect 1 5294 7 5337
rect 1639 5341 1691 5347
rect 59 5329 65 5337
rect 1633 5329 1639 5337
rect 59 5301 1639 5329
rect 59 5294 65 5301
rect 1633 5294 1639 5301
rect 7 5283 59 5289
rect 3271 5341 3323 5347
rect 1691 5329 1697 5337
rect 3265 5329 3271 5337
rect 1691 5301 3271 5329
rect 1691 5294 1697 5301
rect 3265 5294 3271 5301
rect 1639 5283 1691 5289
rect 4903 5341 4955 5347
rect 3323 5329 3329 5337
rect 4897 5329 4903 5337
rect 3323 5301 4903 5329
rect 3323 5294 3329 5301
rect 4897 5294 4903 5301
rect 3271 5283 3323 5289
rect 6535 5341 6587 5347
rect 4955 5329 4961 5337
rect 6529 5329 6535 5337
rect 4955 5301 6535 5329
rect 4955 5294 4961 5301
rect 6529 5294 6535 5301
rect 4903 5283 4955 5289
rect 8167 5341 8219 5347
rect 6587 5329 6593 5337
rect 8161 5329 8167 5337
rect 6587 5301 8167 5329
rect 6587 5294 6593 5301
rect 8161 5294 8167 5301
rect 6535 5283 6587 5289
rect 9799 5341 9851 5347
rect 8219 5329 8225 5337
rect 9793 5329 9799 5337
rect 8219 5301 9799 5329
rect 8219 5294 8225 5301
rect 9793 5294 9799 5301
rect 8167 5283 8219 5289
rect 11431 5341 11483 5347
rect 9851 5329 9857 5337
rect 11425 5329 11431 5337
rect 9851 5301 11431 5329
rect 9851 5294 9857 5301
rect 11425 5294 11431 5301
rect 9799 5283 9851 5289
rect 13063 5341 13115 5347
rect 11483 5329 11489 5337
rect 13057 5329 13063 5337
rect 11483 5301 13063 5329
rect 11483 5294 11489 5301
rect 13057 5294 13063 5301
rect 11431 5283 11483 5289
rect 13115 5294 13121 5337
rect 13063 5283 13115 5289
rect 7 5137 59 5143
rect 1 5090 7 5133
rect 1639 5137 1691 5143
rect 59 5125 65 5133
rect 1633 5125 1639 5133
rect 59 5097 1639 5125
rect 59 5090 65 5097
rect 1633 5090 1639 5097
rect 7 5079 59 5085
rect 3271 5137 3323 5143
rect 1691 5125 1697 5133
rect 3265 5125 3271 5133
rect 1691 5097 3271 5125
rect 1691 5090 1697 5097
rect 3265 5090 3271 5097
rect 1639 5079 1691 5085
rect 4903 5137 4955 5143
rect 3323 5125 3329 5133
rect 4897 5125 4903 5133
rect 3323 5097 4903 5125
rect 3323 5090 3329 5097
rect 4897 5090 4903 5097
rect 3271 5079 3323 5085
rect 6535 5137 6587 5143
rect 4955 5125 4961 5133
rect 6529 5125 6535 5133
rect 4955 5097 6535 5125
rect 4955 5090 4961 5097
rect 6529 5090 6535 5097
rect 4903 5079 4955 5085
rect 8167 5137 8219 5143
rect 6587 5125 6593 5133
rect 8161 5125 8167 5133
rect 6587 5097 8167 5125
rect 6587 5090 6593 5097
rect 8161 5090 8167 5097
rect 6535 5079 6587 5085
rect 9799 5137 9851 5143
rect 8219 5125 8225 5133
rect 9793 5125 9799 5133
rect 8219 5097 9799 5125
rect 8219 5090 8225 5097
rect 9793 5090 9799 5097
rect 8167 5079 8219 5085
rect 11431 5137 11483 5143
rect 9851 5125 9857 5133
rect 11425 5125 11431 5133
rect 9851 5097 11431 5125
rect 9851 5090 9857 5097
rect 11425 5090 11431 5097
rect 9799 5079 9851 5085
rect 13063 5137 13115 5143
rect 11483 5125 11489 5133
rect 13057 5125 13063 5133
rect 11483 5097 13063 5125
rect 11483 5090 11489 5097
rect 13057 5090 13063 5097
rect 11431 5079 11483 5085
rect 13115 5090 13121 5133
rect 13063 5079 13115 5085
rect 7 4933 59 4939
rect 1 4886 7 4929
rect 1639 4933 1691 4939
rect 59 4921 65 4929
rect 1633 4921 1639 4929
rect 59 4893 1639 4921
rect 59 4886 65 4893
rect 1633 4886 1639 4893
rect 7 4875 59 4881
rect 3271 4933 3323 4939
rect 1691 4921 1697 4929
rect 3265 4921 3271 4929
rect 1691 4893 3271 4921
rect 1691 4886 1697 4893
rect 3265 4886 3271 4893
rect 1639 4875 1691 4881
rect 4903 4933 4955 4939
rect 3323 4921 3329 4929
rect 4897 4921 4903 4929
rect 3323 4893 4903 4921
rect 3323 4886 3329 4893
rect 4897 4886 4903 4893
rect 3271 4875 3323 4881
rect 6535 4933 6587 4939
rect 4955 4921 4961 4929
rect 6529 4921 6535 4929
rect 4955 4893 6535 4921
rect 4955 4886 4961 4893
rect 6529 4886 6535 4893
rect 4903 4875 4955 4881
rect 8167 4933 8219 4939
rect 6587 4921 6593 4929
rect 8161 4921 8167 4929
rect 6587 4893 8167 4921
rect 6587 4886 6593 4893
rect 8161 4886 8167 4893
rect 6535 4875 6587 4881
rect 9799 4933 9851 4939
rect 8219 4921 8225 4929
rect 9793 4921 9799 4929
rect 8219 4893 9799 4921
rect 8219 4886 8225 4893
rect 9793 4886 9799 4893
rect 8167 4875 8219 4881
rect 11431 4933 11483 4939
rect 9851 4921 9857 4929
rect 11425 4921 11431 4929
rect 9851 4893 11431 4921
rect 9851 4886 9857 4893
rect 11425 4886 11431 4893
rect 9799 4875 9851 4881
rect 13063 4933 13115 4939
rect 11483 4921 11489 4929
rect 13057 4921 13063 4929
rect 11483 4893 13063 4921
rect 11483 4886 11489 4893
rect 13057 4886 13063 4893
rect 11431 4875 11483 4881
rect 13115 4886 13121 4929
rect 13063 4875 13115 4881
rect 7 4729 59 4735
rect 1 4682 7 4725
rect 1639 4729 1691 4735
rect 59 4717 65 4725
rect 1633 4717 1639 4725
rect 59 4689 1639 4717
rect 59 4682 65 4689
rect 1633 4682 1639 4689
rect 7 4671 59 4677
rect 3271 4729 3323 4735
rect 1691 4717 1697 4725
rect 3265 4717 3271 4725
rect 1691 4689 3271 4717
rect 1691 4682 1697 4689
rect 3265 4682 3271 4689
rect 1639 4671 1691 4677
rect 4903 4729 4955 4735
rect 3323 4717 3329 4725
rect 4897 4717 4903 4725
rect 3323 4689 4903 4717
rect 3323 4682 3329 4689
rect 4897 4682 4903 4689
rect 3271 4671 3323 4677
rect 6535 4729 6587 4735
rect 4955 4717 4961 4725
rect 6529 4717 6535 4725
rect 4955 4689 6535 4717
rect 4955 4682 4961 4689
rect 6529 4682 6535 4689
rect 4903 4671 4955 4677
rect 8167 4729 8219 4735
rect 6587 4717 6593 4725
rect 8161 4717 8167 4725
rect 6587 4689 8167 4717
rect 6587 4682 6593 4689
rect 8161 4682 8167 4689
rect 6535 4671 6587 4677
rect 9799 4729 9851 4735
rect 8219 4717 8225 4725
rect 9793 4717 9799 4725
rect 8219 4689 9799 4717
rect 8219 4682 8225 4689
rect 9793 4682 9799 4689
rect 8167 4671 8219 4677
rect 11431 4729 11483 4735
rect 9851 4717 9857 4725
rect 11425 4717 11431 4725
rect 9851 4689 11431 4717
rect 9851 4682 9857 4689
rect 11425 4682 11431 4689
rect 9799 4671 9851 4677
rect 13063 4729 13115 4735
rect 11483 4717 11489 4725
rect 13057 4717 13063 4725
rect 11483 4689 13063 4717
rect 11483 4682 11489 4689
rect 13057 4682 13063 4689
rect 11431 4671 11483 4677
rect 13115 4682 13121 4725
rect 13063 4671 13115 4677
rect 7 4525 59 4531
rect 1 4478 7 4521
rect 1639 4525 1691 4531
rect 59 4513 65 4521
rect 1633 4513 1639 4521
rect 59 4485 1639 4513
rect 59 4478 65 4485
rect 1633 4478 1639 4485
rect 7 4467 59 4473
rect 3271 4525 3323 4531
rect 1691 4513 1697 4521
rect 3265 4513 3271 4521
rect 1691 4485 3271 4513
rect 1691 4478 1697 4485
rect 3265 4478 3271 4485
rect 1639 4467 1691 4473
rect 4903 4525 4955 4531
rect 3323 4513 3329 4521
rect 4897 4513 4903 4521
rect 3323 4485 4903 4513
rect 3323 4478 3329 4485
rect 4897 4478 4903 4485
rect 3271 4467 3323 4473
rect 6535 4525 6587 4531
rect 4955 4513 4961 4521
rect 6529 4513 6535 4521
rect 4955 4485 6535 4513
rect 4955 4478 4961 4485
rect 6529 4478 6535 4485
rect 4903 4467 4955 4473
rect 8167 4525 8219 4531
rect 6587 4513 6593 4521
rect 8161 4513 8167 4521
rect 6587 4485 8167 4513
rect 6587 4478 6593 4485
rect 8161 4478 8167 4485
rect 6535 4467 6587 4473
rect 9799 4525 9851 4531
rect 8219 4513 8225 4521
rect 9793 4513 9799 4521
rect 8219 4485 9799 4513
rect 8219 4478 8225 4485
rect 9793 4478 9799 4485
rect 8167 4467 8219 4473
rect 11431 4525 11483 4531
rect 9851 4513 9857 4521
rect 11425 4513 11431 4521
rect 9851 4485 11431 4513
rect 9851 4478 9857 4485
rect 11425 4478 11431 4485
rect 9799 4467 9851 4473
rect 13063 4525 13115 4531
rect 11483 4513 11489 4521
rect 13057 4513 13063 4521
rect 11483 4485 13063 4513
rect 11483 4478 11489 4485
rect 13057 4478 13063 4485
rect 11431 4467 11483 4473
rect 13115 4478 13121 4521
rect 13063 4467 13115 4473
rect 212 4319 218 4371
rect 270 4359 276 4371
rect 416 4359 422 4371
rect 270 4331 422 4359
rect 270 4319 276 4331
rect 416 4319 422 4331
rect 474 4359 480 4371
rect 620 4359 626 4371
rect 474 4331 626 4359
rect 474 4319 480 4331
rect 620 4319 626 4331
rect 678 4359 684 4371
rect 824 4359 830 4371
rect 678 4331 830 4359
rect 678 4319 684 4331
rect 824 4319 830 4331
rect 882 4359 888 4371
rect 1028 4359 1034 4371
rect 882 4331 1034 4359
rect 882 4319 888 4331
rect 1028 4319 1034 4331
rect 1086 4359 1092 4371
rect 1232 4359 1238 4371
rect 1086 4331 1238 4359
rect 1086 4319 1092 4331
rect 1232 4319 1238 4331
rect 1290 4359 1296 4371
rect 1436 4359 1442 4371
rect 1290 4331 1442 4359
rect 1290 4319 1296 4331
rect 1436 4319 1442 4331
rect 1494 4359 1500 4371
rect 1640 4359 1646 4371
rect 1494 4331 1646 4359
rect 1494 4319 1500 4331
rect 1640 4319 1646 4331
rect 1698 4359 1704 4371
rect 1844 4359 1850 4371
rect 1698 4331 1850 4359
rect 1698 4319 1704 4331
rect 1844 4319 1850 4331
rect 1902 4359 1908 4371
rect 2048 4359 2054 4371
rect 1902 4331 2054 4359
rect 1902 4319 1908 4331
rect 2048 4319 2054 4331
rect 2106 4359 2112 4371
rect 2252 4359 2258 4371
rect 2106 4331 2258 4359
rect 2106 4319 2112 4331
rect 2252 4319 2258 4331
rect 2310 4359 2316 4371
rect 2456 4359 2462 4371
rect 2310 4331 2462 4359
rect 2310 4319 2316 4331
rect 2456 4319 2462 4331
rect 2514 4359 2520 4371
rect 2660 4359 2666 4371
rect 2514 4331 2666 4359
rect 2514 4319 2520 4331
rect 2660 4319 2666 4331
rect 2718 4359 2724 4371
rect 2864 4359 2870 4371
rect 2718 4331 2870 4359
rect 2718 4319 2724 4331
rect 2864 4319 2870 4331
rect 2922 4359 2928 4371
rect 3068 4359 3074 4371
rect 2922 4331 3074 4359
rect 2922 4319 2928 4331
rect 3068 4319 3074 4331
rect 3126 4359 3132 4371
rect 3272 4359 3278 4371
rect 3126 4331 3278 4359
rect 3126 4319 3132 4331
rect 3272 4319 3278 4331
rect 3330 4359 3336 4371
rect 3476 4359 3482 4371
rect 3330 4331 3482 4359
rect 3330 4319 3336 4331
rect 3476 4319 3482 4331
rect 3534 4359 3540 4371
rect 3680 4359 3686 4371
rect 3534 4331 3686 4359
rect 3534 4319 3540 4331
rect 3680 4319 3686 4331
rect 3738 4359 3744 4371
rect 3884 4359 3890 4371
rect 3738 4331 3890 4359
rect 3738 4319 3744 4331
rect 3884 4319 3890 4331
rect 3942 4359 3948 4371
rect 4088 4359 4094 4371
rect 3942 4331 4094 4359
rect 3942 4319 3948 4331
rect 4088 4319 4094 4331
rect 4146 4359 4152 4371
rect 4292 4359 4298 4371
rect 4146 4331 4298 4359
rect 4146 4319 4152 4331
rect 4292 4319 4298 4331
rect 4350 4359 4356 4371
rect 4496 4359 4502 4371
rect 4350 4331 4502 4359
rect 4350 4319 4356 4331
rect 4496 4319 4502 4331
rect 4554 4359 4560 4371
rect 4700 4359 4706 4371
rect 4554 4331 4706 4359
rect 4554 4319 4560 4331
rect 4700 4319 4706 4331
rect 4758 4359 4764 4371
rect 4904 4359 4910 4371
rect 4758 4331 4910 4359
rect 4758 4319 4764 4331
rect 4904 4319 4910 4331
rect 4962 4359 4968 4371
rect 5108 4359 5114 4371
rect 4962 4331 5114 4359
rect 4962 4319 4968 4331
rect 5108 4319 5114 4331
rect 5166 4359 5172 4371
rect 5312 4359 5318 4371
rect 5166 4331 5318 4359
rect 5166 4319 5172 4331
rect 5312 4319 5318 4331
rect 5370 4359 5376 4371
rect 5516 4359 5522 4371
rect 5370 4331 5522 4359
rect 5370 4319 5376 4331
rect 5516 4319 5522 4331
rect 5574 4359 5580 4371
rect 5720 4359 5726 4371
rect 5574 4331 5726 4359
rect 5574 4319 5580 4331
rect 5720 4319 5726 4331
rect 5778 4359 5784 4371
rect 5924 4359 5930 4371
rect 5778 4331 5930 4359
rect 5778 4319 5784 4331
rect 5924 4319 5930 4331
rect 5982 4359 5988 4371
rect 6128 4359 6134 4371
rect 5982 4331 6134 4359
rect 5982 4319 5988 4331
rect 6128 4319 6134 4331
rect 6186 4359 6192 4371
rect 6332 4359 6338 4371
rect 6186 4331 6338 4359
rect 6186 4319 6192 4331
rect 6332 4319 6338 4331
rect 6390 4359 6396 4371
rect 6536 4359 6542 4371
rect 6390 4331 6542 4359
rect 6390 4319 6396 4331
rect 6536 4319 6542 4331
rect 6594 4359 6600 4371
rect 6740 4359 6746 4371
rect 6594 4331 6746 4359
rect 6594 4319 6600 4331
rect 6740 4319 6746 4331
rect 6798 4359 6804 4371
rect 6944 4359 6950 4371
rect 6798 4331 6950 4359
rect 6798 4319 6804 4331
rect 6944 4319 6950 4331
rect 7002 4359 7008 4371
rect 7148 4359 7154 4371
rect 7002 4331 7154 4359
rect 7002 4319 7008 4331
rect 7148 4319 7154 4331
rect 7206 4359 7212 4371
rect 7352 4359 7358 4371
rect 7206 4331 7358 4359
rect 7206 4319 7212 4331
rect 7352 4319 7358 4331
rect 7410 4359 7416 4371
rect 7556 4359 7562 4371
rect 7410 4331 7562 4359
rect 7410 4319 7416 4331
rect 7556 4319 7562 4331
rect 7614 4359 7620 4371
rect 7760 4359 7766 4371
rect 7614 4331 7766 4359
rect 7614 4319 7620 4331
rect 7760 4319 7766 4331
rect 7818 4359 7824 4371
rect 7964 4359 7970 4371
rect 7818 4331 7970 4359
rect 7818 4319 7824 4331
rect 7964 4319 7970 4331
rect 8022 4359 8028 4371
rect 8168 4359 8174 4371
rect 8022 4331 8174 4359
rect 8022 4319 8028 4331
rect 8168 4319 8174 4331
rect 8226 4359 8232 4371
rect 8372 4359 8378 4371
rect 8226 4331 8378 4359
rect 8226 4319 8232 4331
rect 8372 4319 8378 4331
rect 8430 4359 8436 4371
rect 8576 4359 8582 4371
rect 8430 4331 8582 4359
rect 8430 4319 8436 4331
rect 8576 4319 8582 4331
rect 8634 4359 8640 4371
rect 8780 4359 8786 4371
rect 8634 4331 8786 4359
rect 8634 4319 8640 4331
rect 8780 4319 8786 4331
rect 8838 4359 8844 4371
rect 8984 4359 8990 4371
rect 8838 4331 8990 4359
rect 8838 4319 8844 4331
rect 8984 4319 8990 4331
rect 9042 4359 9048 4371
rect 9188 4359 9194 4371
rect 9042 4331 9194 4359
rect 9042 4319 9048 4331
rect 9188 4319 9194 4331
rect 9246 4359 9252 4371
rect 9392 4359 9398 4371
rect 9246 4331 9398 4359
rect 9246 4319 9252 4331
rect 9392 4319 9398 4331
rect 9450 4359 9456 4371
rect 9596 4359 9602 4371
rect 9450 4331 9602 4359
rect 9450 4319 9456 4331
rect 9596 4319 9602 4331
rect 9654 4359 9660 4371
rect 9800 4359 9806 4371
rect 9654 4331 9806 4359
rect 9654 4319 9660 4331
rect 9800 4319 9806 4331
rect 9858 4359 9864 4371
rect 10004 4359 10010 4371
rect 9858 4331 10010 4359
rect 9858 4319 9864 4331
rect 10004 4319 10010 4331
rect 10062 4359 10068 4371
rect 10208 4359 10214 4371
rect 10062 4331 10214 4359
rect 10062 4319 10068 4331
rect 10208 4319 10214 4331
rect 10266 4359 10272 4371
rect 10412 4359 10418 4371
rect 10266 4331 10418 4359
rect 10266 4319 10272 4331
rect 10412 4319 10418 4331
rect 10470 4359 10476 4371
rect 10616 4359 10622 4371
rect 10470 4331 10622 4359
rect 10470 4319 10476 4331
rect 10616 4319 10622 4331
rect 10674 4359 10680 4371
rect 10820 4359 10826 4371
rect 10674 4331 10826 4359
rect 10674 4319 10680 4331
rect 10820 4319 10826 4331
rect 10878 4359 10884 4371
rect 11024 4359 11030 4371
rect 10878 4331 11030 4359
rect 10878 4319 10884 4331
rect 11024 4319 11030 4331
rect 11082 4359 11088 4371
rect 11228 4359 11234 4371
rect 11082 4331 11234 4359
rect 11082 4319 11088 4331
rect 11228 4319 11234 4331
rect 11286 4359 11292 4371
rect 11432 4359 11438 4371
rect 11286 4331 11438 4359
rect 11286 4319 11292 4331
rect 11432 4319 11438 4331
rect 11490 4359 11496 4371
rect 11636 4359 11642 4371
rect 11490 4331 11642 4359
rect 11490 4319 11496 4331
rect 11636 4319 11642 4331
rect 11694 4359 11700 4371
rect 11840 4359 11846 4371
rect 11694 4331 11846 4359
rect 11694 4319 11700 4331
rect 11840 4319 11846 4331
rect 11898 4359 11904 4371
rect 12044 4359 12050 4371
rect 11898 4331 12050 4359
rect 11898 4319 11904 4331
rect 12044 4319 12050 4331
rect 12102 4359 12108 4371
rect 12248 4359 12254 4371
rect 12102 4331 12254 4359
rect 12102 4319 12108 4331
rect 12248 4319 12254 4331
rect 12306 4359 12312 4371
rect 12452 4359 12458 4371
rect 12306 4331 12458 4359
rect 12306 4319 12312 4331
rect 12452 4319 12458 4331
rect 12510 4359 12516 4371
rect 12656 4359 12662 4371
rect 12510 4331 12662 4359
rect 12510 4319 12516 4331
rect 12656 4319 12662 4331
rect 12714 4359 12720 4371
rect 12860 4359 12866 4371
rect 12714 4331 12866 4359
rect 12714 4319 12720 4331
rect 12860 4319 12866 4331
rect 12918 4359 12924 4371
rect 13078 4359 13084 4371
rect 12918 4331 13084 4359
rect 12918 4319 12924 4331
rect 13078 4319 13084 4331
rect 13136 4319 13142 4371
rect 7 4217 59 4223
rect 1 4170 7 4213
rect 1639 4217 1691 4223
rect 59 4205 65 4213
rect 1633 4205 1639 4213
rect 59 4177 1639 4205
rect 59 4170 65 4177
rect 1633 4170 1639 4177
rect 7 4159 59 4165
rect 3271 4217 3323 4223
rect 1691 4205 1697 4213
rect 3265 4205 3271 4213
rect 1691 4177 3271 4205
rect 1691 4170 1697 4177
rect 3265 4170 3271 4177
rect 1639 4159 1691 4165
rect 4903 4217 4955 4223
rect 3323 4205 3329 4213
rect 4897 4205 4903 4213
rect 3323 4177 4903 4205
rect 3323 4170 3329 4177
rect 4897 4170 4903 4177
rect 3271 4159 3323 4165
rect 6535 4217 6587 4223
rect 4955 4205 4961 4213
rect 6529 4205 6535 4213
rect 4955 4177 6535 4205
rect 4955 4170 4961 4177
rect 6529 4170 6535 4177
rect 4903 4159 4955 4165
rect 8167 4217 8219 4223
rect 6587 4205 6593 4213
rect 8161 4205 8167 4213
rect 6587 4177 8167 4205
rect 6587 4170 6593 4177
rect 8161 4170 8167 4177
rect 6535 4159 6587 4165
rect 9799 4217 9851 4223
rect 8219 4205 8225 4213
rect 9793 4205 9799 4213
rect 8219 4177 9799 4205
rect 8219 4170 8225 4177
rect 9793 4170 9799 4177
rect 8167 4159 8219 4165
rect 11431 4217 11483 4223
rect 9851 4205 9857 4213
rect 11425 4205 11431 4213
rect 9851 4177 11431 4205
rect 9851 4170 9857 4177
rect 11425 4170 11431 4177
rect 9799 4159 9851 4165
rect 13063 4217 13115 4223
rect 11483 4205 11489 4213
rect 13057 4205 13063 4213
rect 11483 4177 13063 4205
rect 11483 4170 11489 4177
rect 13057 4170 13063 4177
rect 11431 4159 11483 4165
rect 13115 4170 13121 4213
rect 13063 4159 13115 4165
rect 7 4013 59 4019
rect 1 3966 7 4009
rect 1639 4013 1691 4019
rect 59 4001 65 4009
rect 1633 4001 1639 4009
rect 59 3973 1639 4001
rect 59 3966 65 3973
rect 1633 3966 1639 3973
rect 7 3955 59 3961
rect 3271 4013 3323 4019
rect 1691 4001 1697 4009
rect 3265 4001 3271 4009
rect 1691 3973 3271 4001
rect 1691 3966 1697 3973
rect 3265 3966 3271 3973
rect 1639 3955 1691 3961
rect 4903 4013 4955 4019
rect 3323 4001 3329 4009
rect 4897 4001 4903 4009
rect 3323 3973 4903 4001
rect 3323 3966 3329 3973
rect 4897 3966 4903 3973
rect 3271 3955 3323 3961
rect 6535 4013 6587 4019
rect 4955 4001 4961 4009
rect 6529 4001 6535 4009
rect 4955 3973 6535 4001
rect 4955 3966 4961 3973
rect 6529 3966 6535 3973
rect 4903 3955 4955 3961
rect 8167 4013 8219 4019
rect 6587 4001 6593 4009
rect 8161 4001 8167 4009
rect 6587 3973 8167 4001
rect 6587 3966 6593 3973
rect 8161 3966 8167 3973
rect 6535 3955 6587 3961
rect 9799 4013 9851 4019
rect 8219 4001 8225 4009
rect 9793 4001 9799 4009
rect 8219 3973 9799 4001
rect 8219 3966 8225 3973
rect 9793 3966 9799 3973
rect 8167 3955 8219 3961
rect 11431 4013 11483 4019
rect 9851 4001 9857 4009
rect 11425 4001 11431 4009
rect 9851 3973 11431 4001
rect 9851 3966 9857 3973
rect 11425 3966 11431 3973
rect 9799 3955 9851 3961
rect 13063 4013 13115 4019
rect 11483 4001 11489 4009
rect 13057 4001 13063 4009
rect 11483 3973 13063 4001
rect 11483 3966 11489 3973
rect 13057 3966 13063 3973
rect 11431 3955 11483 3961
rect 13115 3966 13121 4009
rect 13063 3955 13115 3961
rect 7 3809 59 3815
rect 1 3762 7 3805
rect 1639 3809 1691 3815
rect 59 3797 65 3805
rect 1633 3797 1639 3805
rect 59 3769 1639 3797
rect 59 3762 65 3769
rect 1633 3762 1639 3769
rect 7 3751 59 3757
rect 3271 3809 3323 3815
rect 1691 3797 1697 3805
rect 3265 3797 3271 3805
rect 1691 3769 3271 3797
rect 1691 3762 1697 3769
rect 3265 3762 3271 3769
rect 1639 3751 1691 3757
rect 4903 3809 4955 3815
rect 3323 3797 3329 3805
rect 4897 3797 4903 3805
rect 3323 3769 4903 3797
rect 3323 3762 3329 3769
rect 4897 3762 4903 3769
rect 3271 3751 3323 3757
rect 6535 3809 6587 3815
rect 4955 3797 4961 3805
rect 6529 3797 6535 3805
rect 4955 3769 6535 3797
rect 4955 3762 4961 3769
rect 6529 3762 6535 3769
rect 4903 3751 4955 3757
rect 8167 3809 8219 3815
rect 6587 3797 6593 3805
rect 8161 3797 8167 3805
rect 6587 3769 8167 3797
rect 6587 3762 6593 3769
rect 8161 3762 8167 3769
rect 6535 3751 6587 3757
rect 9799 3809 9851 3815
rect 8219 3797 8225 3805
rect 9793 3797 9799 3805
rect 8219 3769 9799 3797
rect 8219 3762 8225 3769
rect 9793 3762 9799 3769
rect 8167 3751 8219 3757
rect 11431 3809 11483 3815
rect 9851 3797 9857 3805
rect 11425 3797 11431 3805
rect 9851 3769 11431 3797
rect 9851 3762 9857 3769
rect 11425 3762 11431 3769
rect 9799 3751 9851 3757
rect 13063 3809 13115 3815
rect 11483 3797 11489 3805
rect 13057 3797 13063 3805
rect 11483 3769 13063 3797
rect 11483 3762 11489 3769
rect 13057 3762 13063 3769
rect 11431 3751 11483 3757
rect 13115 3762 13121 3805
rect 13063 3751 13115 3757
rect 7 3605 59 3611
rect 1 3558 7 3601
rect 1639 3605 1691 3611
rect 59 3593 65 3601
rect 1633 3593 1639 3601
rect 59 3565 1639 3593
rect 59 3558 65 3565
rect 1633 3558 1639 3565
rect 7 3547 59 3553
rect 3271 3605 3323 3611
rect 1691 3593 1697 3601
rect 3265 3593 3271 3601
rect 1691 3565 3271 3593
rect 1691 3558 1697 3565
rect 3265 3558 3271 3565
rect 1639 3547 1691 3553
rect 4903 3605 4955 3611
rect 3323 3593 3329 3601
rect 4897 3593 4903 3601
rect 3323 3565 4903 3593
rect 3323 3558 3329 3565
rect 4897 3558 4903 3565
rect 3271 3547 3323 3553
rect 6535 3605 6587 3611
rect 4955 3593 4961 3601
rect 6529 3593 6535 3601
rect 4955 3565 6535 3593
rect 4955 3558 4961 3565
rect 6529 3558 6535 3565
rect 4903 3547 4955 3553
rect 8167 3605 8219 3611
rect 6587 3593 6593 3601
rect 8161 3593 8167 3601
rect 6587 3565 8167 3593
rect 6587 3558 6593 3565
rect 8161 3558 8167 3565
rect 6535 3547 6587 3553
rect 9799 3605 9851 3611
rect 8219 3593 8225 3601
rect 9793 3593 9799 3601
rect 8219 3565 9799 3593
rect 8219 3558 8225 3565
rect 9793 3558 9799 3565
rect 8167 3547 8219 3553
rect 11431 3605 11483 3611
rect 9851 3593 9857 3601
rect 11425 3593 11431 3601
rect 9851 3565 11431 3593
rect 9851 3558 9857 3565
rect 11425 3558 11431 3565
rect 9799 3547 9851 3553
rect 13063 3605 13115 3611
rect 11483 3593 11489 3601
rect 13057 3593 13063 3601
rect 11483 3565 13063 3593
rect 11483 3558 11489 3565
rect 13057 3558 13063 3565
rect 11431 3547 11483 3553
rect 13115 3558 13121 3601
rect 13063 3547 13115 3553
rect 7 3401 59 3407
rect 1 3354 7 3397
rect 1639 3401 1691 3407
rect 59 3389 65 3397
rect 1633 3389 1639 3397
rect 59 3361 1639 3389
rect 59 3354 65 3361
rect 1633 3354 1639 3361
rect 7 3343 59 3349
rect 3271 3401 3323 3407
rect 1691 3389 1697 3397
rect 3265 3389 3271 3397
rect 1691 3361 3271 3389
rect 1691 3354 1697 3361
rect 3265 3354 3271 3361
rect 1639 3343 1691 3349
rect 4903 3401 4955 3407
rect 3323 3389 3329 3397
rect 4897 3389 4903 3397
rect 3323 3361 4903 3389
rect 3323 3354 3329 3361
rect 4897 3354 4903 3361
rect 3271 3343 3323 3349
rect 6535 3401 6587 3407
rect 4955 3389 4961 3397
rect 6529 3389 6535 3397
rect 4955 3361 6535 3389
rect 4955 3354 4961 3361
rect 6529 3354 6535 3361
rect 4903 3343 4955 3349
rect 8167 3401 8219 3407
rect 6587 3389 6593 3397
rect 8161 3389 8167 3397
rect 6587 3361 8167 3389
rect 6587 3354 6593 3361
rect 8161 3354 8167 3361
rect 6535 3343 6587 3349
rect 9799 3401 9851 3407
rect 8219 3389 8225 3397
rect 9793 3389 9799 3397
rect 8219 3361 9799 3389
rect 8219 3354 8225 3361
rect 9793 3354 9799 3361
rect 8167 3343 8219 3349
rect 11431 3401 11483 3407
rect 9851 3389 9857 3397
rect 11425 3389 11431 3397
rect 9851 3361 11431 3389
rect 9851 3354 9857 3361
rect 11425 3354 11431 3361
rect 9799 3343 9851 3349
rect 13063 3401 13115 3407
rect 11483 3389 11489 3397
rect 13057 3389 13063 3397
rect 11483 3361 13063 3389
rect 11483 3354 11489 3361
rect 13057 3354 13063 3361
rect 11431 3343 11483 3349
rect 13115 3354 13121 3397
rect 13063 3343 13115 3349
rect 7 3197 59 3203
rect 1 3150 7 3193
rect 1639 3197 1691 3203
rect 59 3185 65 3193
rect 1633 3185 1639 3193
rect 59 3157 1639 3185
rect 59 3150 65 3157
rect 1633 3150 1639 3157
rect 7 3139 59 3145
rect 3271 3197 3323 3203
rect 1691 3185 1697 3193
rect 3265 3185 3271 3193
rect 1691 3157 3271 3185
rect 1691 3150 1697 3157
rect 3265 3150 3271 3157
rect 1639 3139 1691 3145
rect 4903 3197 4955 3203
rect 3323 3185 3329 3193
rect 4897 3185 4903 3193
rect 3323 3157 4903 3185
rect 3323 3150 3329 3157
rect 4897 3150 4903 3157
rect 3271 3139 3323 3145
rect 6535 3197 6587 3203
rect 4955 3185 4961 3193
rect 6529 3185 6535 3193
rect 4955 3157 6535 3185
rect 4955 3150 4961 3157
rect 6529 3150 6535 3157
rect 4903 3139 4955 3145
rect 8167 3197 8219 3203
rect 6587 3185 6593 3193
rect 8161 3185 8167 3193
rect 6587 3157 8167 3185
rect 6587 3150 6593 3157
rect 8161 3150 8167 3157
rect 6535 3139 6587 3145
rect 9799 3197 9851 3203
rect 8219 3185 8225 3193
rect 9793 3185 9799 3193
rect 8219 3157 9799 3185
rect 8219 3150 8225 3157
rect 9793 3150 9799 3157
rect 8167 3139 8219 3145
rect 11431 3197 11483 3203
rect 9851 3185 9857 3193
rect 11425 3185 11431 3193
rect 9851 3157 11431 3185
rect 9851 3150 9857 3157
rect 11425 3150 11431 3157
rect 9799 3139 9851 3145
rect 13063 3197 13115 3203
rect 11483 3185 11489 3193
rect 13057 3185 13063 3193
rect 11483 3157 13063 3185
rect 11483 3150 11489 3157
rect 13057 3150 13063 3157
rect 11431 3139 11483 3145
rect 13115 3150 13121 3193
rect 13063 3139 13115 3145
rect 7 2993 59 2999
rect 1 2946 7 2989
rect 1639 2993 1691 2999
rect 59 2981 65 2989
rect 1633 2981 1639 2989
rect 59 2953 1639 2981
rect 59 2946 65 2953
rect 1633 2946 1639 2953
rect 7 2935 59 2941
rect 3271 2993 3323 2999
rect 1691 2981 1697 2989
rect 3265 2981 3271 2989
rect 1691 2953 3271 2981
rect 1691 2946 1697 2953
rect 3265 2946 3271 2953
rect 1639 2935 1691 2941
rect 4903 2993 4955 2999
rect 3323 2981 3329 2989
rect 4897 2981 4903 2989
rect 3323 2953 4903 2981
rect 3323 2946 3329 2953
rect 4897 2946 4903 2953
rect 3271 2935 3323 2941
rect 6535 2993 6587 2999
rect 4955 2981 4961 2989
rect 6529 2981 6535 2989
rect 4955 2953 6535 2981
rect 4955 2946 4961 2953
rect 6529 2946 6535 2953
rect 4903 2935 4955 2941
rect 8167 2993 8219 2999
rect 6587 2981 6593 2989
rect 8161 2981 8167 2989
rect 6587 2953 8167 2981
rect 6587 2946 6593 2953
rect 8161 2946 8167 2953
rect 6535 2935 6587 2941
rect 9799 2993 9851 2999
rect 8219 2981 8225 2989
rect 9793 2981 9799 2989
rect 8219 2953 9799 2981
rect 8219 2946 8225 2953
rect 9793 2946 9799 2953
rect 8167 2935 8219 2941
rect 11431 2993 11483 2999
rect 9851 2981 9857 2989
rect 11425 2981 11431 2989
rect 9851 2953 11431 2981
rect 9851 2946 9857 2953
rect 11425 2946 11431 2953
rect 9799 2935 9851 2941
rect 13063 2993 13115 2999
rect 11483 2981 11489 2989
rect 13057 2981 13063 2989
rect 11483 2953 13063 2981
rect 11483 2946 11489 2953
rect 13057 2946 13063 2953
rect 11431 2935 11483 2941
rect 13115 2946 13121 2989
rect 13063 2935 13115 2941
rect 7 2789 59 2795
rect 1 2742 7 2785
rect 1639 2789 1691 2795
rect 59 2777 65 2785
rect 1633 2777 1639 2785
rect 59 2749 1639 2777
rect 59 2742 65 2749
rect 1633 2742 1639 2749
rect 7 2731 59 2737
rect 3271 2789 3323 2795
rect 1691 2777 1697 2785
rect 3265 2777 3271 2785
rect 1691 2749 3271 2777
rect 1691 2742 1697 2749
rect 3265 2742 3271 2749
rect 1639 2731 1691 2737
rect 4903 2789 4955 2795
rect 3323 2777 3329 2785
rect 4897 2777 4903 2785
rect 3323 2749 4903 2777
rect 3323 2742 3329 2749
rect 4897 2742 4903 2749
rect 3271 2731 3323 2737
rect 6535 2789 6587 2795
rect 4955 2777 4961 2785
rect 6529 2777 6535 2785
rect 4955 2749 6535 2777
rect 4955 2742 4961 2749
rect 6529 2742 6535 2749
rect 4903 2731 4955 2737
rect 8167 2789 8219 2795
rect 6587 2777 6593 2785
rect 8161 2777 8167 2785
rect 6587 2749 8167 2777
rect 6587 2742 6593 2749
rect 8161 2742 8167 2749
rect 6535 2731 6587 2737
rect 9799 2789 9851 2795
rect 8219 2777 8225 2785
rect 9793 2777 9799 2785
rect 8219 2749 9799 2777
rect 8219 2742 8225 2749
rect 9793 2742 9799 2749
rect 8167 2731 8219 2737
rect 11431 2789 11483 2795
rect 9851 2777 9857 2785
rect 11425 2777 11431 2785
rect 9851 2749 11431 2777
rect 9851 2742 9857 2749
rect 11425 2742 11431 2749
rect 9799 2731 9851 2737
rect 13063 2789 13115 2795
rect 11483 2777 11489 2785
rect 13057 2777 13063 2785
rect 11483 2749 13063 2777
rect 11483 2742 11489 2749
rect 13057 2742 13063 2749
rect 11431 2731 11483 2737
rect 13115 2742 13121 2785
rect 13063 2731 13115 2737
rect 212 2583 218 2635
rect 270 2623 276 2635
rect 416 2623 422 2635
rect 270 2595 422 2623
rect 270 2583 276 2595
rect 416 2583 422 2595
rect 474 2623 480 2635
rect 620 2623 626 2635
rect 474 2595 626 2623
rect 474 2583 480 2595
rect 620 2583 626 2595
rect 678 2623 684 2635
rect 824 2623 830 2635
rect 678 2595 830 2623
rect 678 2583 684 2595
rect 824 2583 830 2595
rect 882 2623 888 2635
rect 1028 2623 1034 2635
rect 882 2595 1034 2623
rect 882 2583 888 2595
rect 1028 2583 1034 2595
rect 1086 2623 1092 2635
rect 1232 2623 1238 2635
rect 1086 2595 1238 2623
rect 1086 2583 1092 2595
rect 1232 2583 1238 2595
rect 1290 2623 1296 2635
rect 1436 2623 1442 2635
rect 1290 2595 1442 2623
rect 1290 2583 1296 2595
rect 1436 2583 1442 2595
rect 1494 2623 1500 2635
rect 1640 2623 1646 2635
rect 1494 2595 1646 2623
rect 1494 2583 1500 2595
rect 1640 2583 1646 2595
rect 1698 2623 1704 2635
rect 1844 2623 1850 2635
rect 1698 2595 1850 2623
rect 1698 2583 1704 2595
rect 1844 2583 1850 2595
rect 1902 2623 1908 2635
rect 2048 2623 2054 2635
rect 1902 2595 2054 2623
rect 1902 2583 1908 2595
rect 2048 2583 2054 2595
rect 2106 2623 2112 2635
rect 2252 2623 2258 2635
rect 2106 2595 2258 2623
rect 2106 2583 2112 2595
rect 2252 2583 2258 2595
rect 2310 2623 2316 2635
rect 2456 2623 2462 2635
rect 2310 2595 2462 2623
rect 2310 2583 2316 2595
rect 2456 2583 2462 2595
rect 2514 2623 2520 2635
rect 2660 2623 2666 2635
rect 2514 2595 2666 2623
rect 2514 2583 2520 2595
rect 2660 2583 2666 2595
rect 2718 2623 2724 2635
rect 2864 2623 2870 2635
rect 2718 2595 2870 2623
rect 2718 2583 2724 2595
rect 2864 2583 2870 2595
rect 2922 2623 2928 2635
rect 3068 2623 3074 2635
rect 2922 2595 3074 2623
rect 2922 2583 2928 2595
rect 3068 2583 3074 2595
rect 3126 2623 3132 2635
rect 3272 2623 3278 2635
rect 3126 2595 3278 2623
rect 3126 2583 3132 2595
rect 3272 2583 3278 2595
rect 3330 2623 3336 2635
rect 3476 2623 3482 2635
rect 3330 2595 3482 2623
rect 3330 2583 3336 2595
rect 3476 2583 3482 2595
rect 3534 2623 3540 2635
rect 3680 2623 3686 2635
rect 3534 2595 3686 2623
rect 3534 2583 3540 2595
rect 3680 2583 3686 2595
rect 3738 2623 3744 2635
rect 3884 2623 3890 2635
rect 3738 2595 3890 2623
rect 3738 2583 3744 2595
rect 3884 2583 3890 2595
rect 3942 2623 3948 2635
rect 4088 2623 4094 2635
rect 3942 2595 4094 2623
rect 3942 2583 3948 2595
rect 4088 2583 4094 2595
rect 4146 2623 4152 2635
rect 4292 2623 4298 2635
rect 4146 2595 4298 2623
rect 4146 2583 4152 2595
rect 4292 2583 4298 2595
rect 4350 2623 4356 2635
rect 4496 2623 4502 2635
rect 4350 2595 4502 2623
rect 4350 2583 4356 2595
rect 4496 2583 4502 2595
rect 4554 2623 4560 2635
rect 4700 2623 4706 2635
rect 4554 2595 4706 2623
rect 4554 2583 4560 2595
rect 4700 2583 4706 2595
rect 4758 2623 4764 2635
rect 4904 2623 4910 2635
rect 4758 2595 4910 2623
rect 4758 2583 4764 2595
rect 4904 2583 4910 2595
rect 4962 2623 4968 2635
rect 5108 2623 5114 2635
rect 4962 2595 5114 2623
rect 4962 2583 4968 2595
rect 5108 2583 5114 2595
rect 5166 2623 5172 2635
rect 5312 2623 5318 2635
rect 5166 2595 5318 2623
rect 5166 2583 5172 2595
rect 5312 2583 5318 2595
rect 5370 2623 5376 2635
rect 5516 2623 5522 2635
rect 5370 2595 5522 2623
rect 5370 2583 5376 2595
rect 5516 2583 5522 2595
rect 5574 2623 5580 2635
rect 5720 2623 5726 2635
rect 5574 2595 5726 2623
rect 5574 2583 5580 2595
rect 5720 2583 5726 2595
rect 5778 2623 5784 2635
rect 5924 2623 5930 2635
rect 5778 2595 5930 2623
rect 5778 2583 5784 2595
rect 5924 2583 5930 2595
rect 5982 2623 5988 2635
rect 6128 2623 6134 2635
rect 5982 2595 6134 2623
rect 5982 2583 5988 2595
rect 6128 2583 6134 2595
rect 6186 2623 6192 2635
rect 6332 2623 6338 2635
rect 6186 2595 6338 2623
rect 6186 2583 6192 2595
rect 6332 2583 6338 2595
rect 6390 2623 6396 2635
rect 6536 2623 6542 2635
rect 6390 2595 6542 2623
rect 6390 2583 6396 2595
rect 6536 2583 6542 2595
rect 6594 2623 6600 2635
rect 6740 2623 6746 2635
rect 6594 2595 6746 2623
rect 6594 2583 6600 2595
rect 6740 2583 6746 2595
rect 6798 2623 6804 2635
rect 6944 2623 6950 2635
rect 6798 2595 6950 2623
rect 6798 2583 6804 2595
rect 6944 2583 6950 2595
rect 7002 2623 7008 2635
rect 7148 2623 7154 2635
rect 7002 2595 7154 2623
rect 7002 2583 7008 2595
rect 7148 2583 7154 2595
rect 7206 2623 7212 2635
rect 7352 2623 7358 2635
rect 7206 2595 7358 2623
rect 7206 2583 7212 2595
rect 7352 2583 7358 2595
rect 7410 2623 7416 2635
rect 7556 2623 7562 2635
rect 7410 2595 7562 2623
rect 7410 2583 7416 2595
rect 7556 2583 7562 2595
rect 7614 2623 7620 2635
rect 7760 2623 7766 2635
rect 7614 2595 7766 2623
rect 7614 2583 7620 2595
rect 7760 2583 7766 2595
rect 7818 2623 7824 2635
rect 7964 2623 7970 2635
rect 7818 2595 7970 2623
rect 7818 2583 7824 2595
rect 7964 2583 7970 2595
rect 8022 2623 8028 2635
rect 8168 2623 8174 2635
rect 8022 2595 8174 2623
rect 8022 2583 8028 2595
rect 8168 2583 8174 2595
rect 8226 2623 8232 2635
rect 8372 2623 8378 2635
rect 8226 2595 8378 2623
rect 8226 2583 8232 2595
rect 8372 2583 8378 2595
rect 8430 2623 8436 2635
rect 8576 2623 8582 2635
rect 8430 2595 8582 2623
rect 8430 2583 8436 2595
rect 8576 2583 8582 2595
rect 8634 2623 8640 2635
rect 8780 2623 8786 2635
rect 8634 2595 8786 2623
rect 8634 2583 8640 2595
rect 8780 2583 8786 2595
rect 8838 2623 8844 2635
rect 8984 2623 8990 2635
rect 8838 2595 8990 2623
rect 8838 2583 8844 2595
rect 8984 2583 8990 2595
rect 9042 2623 9048 2635
rect 9188 2623 9194 2635
rect 9042 2595 9194 2623
rect 9042 2583 9048 2595
rect 9188 2583 9194 2595
rect 9246 2623 9252 2635
rect 9392 2623 9398 2635
rect 9246 2595 9398 2623
rect 9246 2583 9252 2595
rect 9392 2583 9398 2595
rect 9450 2623 9456 2635
rect 9596 2623 9602 2635
rect 9450 2595 9602 2623
rect 9450 2583 9456 2595
rect 9596 2583 9602 2595
rect 9654 2623 9660 2635
rect 9800 2623 9806 2635
rect 9654 2595 9806 2623
rect 9654 2583 9660 2595
rect 9800 2583 9806 2595
rect 9858 2623 9864 2635
rect 10004 2623 10010 2635
rect 9858 2595 10010 2623
rect 9858 2583 9864 2595
rect 10004 2583 10010 2595
rect 10062 2623 10068 2635
rect 10208 2623 10214 2635
rect 10062 2595 10214 2623
rect 10062 2583 10068 2595
rect 10208 2583 10214 2595
rect 10266 2623 10272 2635
rect 10412 2623 10418 2635
rect 10266 2595 10418 2623
rect 10266 2583 10272 2595
rect 10412 2583 10418 2595
rect 10470 2623 10476 2635
rect 10616 2623 10622 2635
rect 10470 2595 10622 2623
rect 10470 2583 10476 2595
rect 10616 2583 10622 2595
rect 10674 2623 10680 2635
rect 10820 2623 10826 2635
rect 10674 2595 10826 2623
rect 10674 2583 10680 2595
rect 10820 2583 10826 2595
rect 10878 2623 10884 2635
rect 11024 2623 11030 2635
rect 10878 2595 11030 2623
rect 10878 2583 10884 2595
rect 11024 2583 11030 2595
rect 11082 2623 11088 2635
rect 11228 2623 11234 2635
rect 11082 2595 11234 2623
rect 11082 2583 11088 2595
rect 11228 2583 11234 2595
rect 11286 2623 11292 2635
rect 11432 2623 11438 2635
rect 11286 2595 11438 2623
rect 11286 2583 11292 2595
rect 11432 2583 11438 2595
rect 11490 2623 11496 2635
rect 11636 2623 11642 2635
rect 11490 2595 11642 2623
rect 11490 2583 11496 2595
rect 11636 2583 11642 2595
rect 11694 2623 11700 2635
rect 11840 2623 11846 2635
rect 11694 2595 11846 2623
rect 11694 2583 11700 2595
rect 11840 2583 11846 2595
rect 11898 2623 11904 2635
rect 12044 2623 12050 2635
rect 11898 2595 12050 2623
rect 11898 2583 11904 2595
rect 12044 2583 12050 2595
rect 12102 2623 12108 2635
rect 12248 2623 12254 2635
rect 12102 2595 12254 2623
rect 12102 2583 12108 2595
rect 12248 2583 12254 2595
rect 12306 2623 12312 2635
rect 12452 2623 12458 2635
rect 12306 2595 12458 2623
rect 12306 2583 12312 2595
rect 12452 2583 12458 2595
rect 12510 2623 12516 2635
rect 12656 2623 12662 2635
rect 12510 2595 12662 2623
rect 12510 2583 12516 2595
rect 12656 2583 12662 2595
rect 12714 2623 12720 2635
rect 12860 2623 12866 2635
rect 12714 2595 12866 2623
rect 12714 2583 12720 2595
rect 12860 2583 12866 2595
rect 12918 2623 12924 2635
rect 13078 2623 13084 2635
rect 12918 2595 13084 2623
rect 12918 2583 12924 2595
rect 13078 2583 13084 2595
rect 13136 2583 13142 2635
rect 7 2481 59 2487
rect 1 2434 7 2477
rect 1639 2481 1691 2487
rect 59 2469 65 2477
rect 1633 2469 1639 2477
rect 59 2441 1639 2469
rect 59 2434 65 2441
rect 1633 2434 1639 2441
rect 7 2423 59 2429
rect 3271 2481 3323 2487
rect 1691 2469 1697 2477
rect 3265 2469 3271 2477
rect 1691 2441 3271 2469
rect 1691 2434 1697 2441
rect 3265 2434 3271 2441
rect 1639 2423 1691 2429
rect 4903 2481 4955 2487
rect 3323 2469 3329 2477
rect 4897 2469 4903 2477
rect 3323 2441 4903 2469
rect 3323 2434 3329 2441
rect 4897 2434 4903 2441
rect 3271 2423 3323 2429
rect 6535 2481 6587 2487
rect 4955 2469 4961 2477
rect 6529 2469 6535 2477
rect 4955 2441 6535 2469
rect 4955 2434 4961 2441
rect 6529 2434 6535 2441
rect 4903 2423 4955 2429
rect 8167 2481 8219 2487
rect 6587 2469 6593 2477
rect 8161 2469 8167 2477
rect 6587 2441 8167 2469
rect 6587 2434 6593 2441
rect 8161 2434 8167 2441
rect 6535 2423 6587 2429
rect 9799 2481 9851 2487
rect 8219 2469 8225 2477
rect 9793 2469 9799 2477
rect 8219 2441 9799 2469
rect 8219 2434 8225 2441
rect 9793 2434 9799 2441
rect 8167 2423 8219 2429
rect 11431 2481 11483 2487
rect 9851 2469 9857 2477
rect 11425 2469 11431 2477
rect 9851 2441 11431 2469
rect 9851 2434 9857 2441
rect 11425 2434 11431 2441
rect 9799 2423 9851 2429
rect 13063 2481 13115 2487
rect 11483 2469 11489 2477
rect 13057 2469 13063 2477
rect 11483 2441 13063 2469
rect 11483 2434 11489 2441
rect 13057 2434 13063 2441
rect 11431 2423 11483 2429
rect 13115 2434 13121 2477
rect 13063 2423 13115 2429
rect 7 2277 59 2283
rect 1 2230 7 2273
rect 1639 2277 1691 2283
rect 59 2265 65 2273
rect 1633 2265 1639 2273
rect 59 2237 1639 2265
rect 59 2230 65 2237
rect 1633 2230 1639 2237
rect 7 2219 59 2225
rect 3271 2277 3323 2283
rect 1691 2265 1697 2273
rect 3265 2265 3271 2273
rect 1691 2237 3271 2265
rect 1691 2230 1697 2237
rect 3265 2230 3271 2237
rect 1639 2219 1691 2225
rect 4903 2277 4955 2283
rect 3323 2265 3329 2273
rect 4897 2265 4903 2273
rect 3323 2237 4903 2265
rect 3323 2230 3329 2237
rect 4897 2230 4903 2237
rect 3271 2219 3323 2225
rect 6535 2277 6587 2283
rect 4955 2265 4961 2273
rect 6529 2265 6535 2273
rect 4955 2237 6535 2265
rect 4955 2230 4961 2237
rect 6529 2230 6535 2237
rect 4903 2219 4955 2225
rect 8167 2277 8219 2283
rect 6587 2265 6593 2273
rect 8161 2265 8167 2273
rect 6587 2237 8167 2265
rect 6587 2230 6593 2237
rect 8161 2230 8167 2237
rect 6535 2219 6587 2225
rect 9799 2277 9851 2283
rect 8219 2265 8225 2273
rect 9793 2265 9799 2273
rect 8219 2237 9799 2265
rect 8219 2230 8225 2237
rect 9793 2230 9799 2237
rect 8167 2219 8219 2225
rect 11431 2277 11483 2283
rect 9851 2265 9857 2273
rect 11425 2265 11431 2273
rect 9851 2237 11431 2265
rect 9851 2230 9857 2237
rect 11425 2230 11431 2237
rect 9799 2219 9851 2225
rect 13063 2277 13115 2283
rect 11483 2265 11489 2273
rect 13057 2265 13063 2273
rect 11483 2237 13063 2265
rect 11483 2230 11489 2237
rect 13057 2230 13063 2237
rect 11431 2219 11483 2225
rect 13115 2230 13121 2273
rect 13063 2219 13115 2225
rect 7 2073 59 2079
rect 1 2026 7 2069
rect 1639 2073 1691 2079
rect 59 2061 65 2069
rect 1633 2061 1639 2069
rect 59 2033 1639 2061
rect 59 2026 65 2033
rect 1633 2026 1639 2033
rect 7 2015 59 2021
rect 3271 2073 3323 2079
rect 1691 2061 1697 2069
rect 3265 2061 3271 2069
rect 1691 2033 3271 2061
rect 1691 2026 1697 2033
rect 3265 2026 3271 2033
rect 1639 2015 1691 2021
rect 4903 2073 4955 2079
rect 3323 2061 3329 2069
rect 4897 2061 4903 2069
rect 3323 2033 4903 2061
rect 3323 2026 3329 2033
rect 4897 2026 4903 2033
rect 3271 2015 3323 2021
rect 6535 2073 6587 2079
rect 4955 2061 4961 2069
rect 6529 2061 6535 2069
rect 4955 2033 6535 2061
rect 4955 2026 4961 2033
rect 6529 2026 6535 2033
rect 4903 2015 4955 2021
rect 8167 2073 8219 2079
rect 6587 2061 6593 2069
rect 8161 2061 8167 2069
rect 6587 2033 8167 2061
rect 6587 2026 6593 2033
rect 8161 2026 8167 2033
rect 6535 2015 6587 2021
rect 9799 2073 9851 2079
rect 8219 2061 8225 2069
rect 9793 2061 9799 2069
rect 8219 2033 9799 2061
rect 8219 2026 8225 2033
rect 9793 2026 9799 2033
rect 8167 2015 8219 2021
rect 11431 2073 11483 2079
rect 9851 2061 9857 2069
rect 11425 2061 11431 2069
rect 9851 2033 11431 2061
rect 9851 2026 9857 2033
rect 11425 2026 11431 2033
rect 9799 2015 9851 2021
rect 13063 2073 13115 2079
rect 11483 2061 11489 2069
rect 13057 2061 13063 2069
rect 11483 2033 13063 2061
rect 11483 2026 11489 2033
rect 13057 2026 13063 2033
rect 11431 2015 11483 2021
rect 13115 2026 13121 2069
rect 13063 2015 13115 2021
rect 7 1869 59 1875
rect 1 1822 7 1865
rect 1639 1869 1691 1875
rect 59 1857 65 1865
rect 1633 1857 1639 1865
rect 59 1829 1639 1857
rect 59 1822 65 1829
rect 1633 1822 1639 1829
rect 7 1811 59 1817
rect 3271 1869 3323 1875
rect 1691 1857 1697 1865
rect 3265 1857 3271 1865
rect 1691 1829 3271 1857
rect 1691 1822 1697 1829
rect 3265 1822 3271 1829
rect 1639 1811 1691 1817
rect 4903 1869 4955 1875
rect 3323 1857 3329 1865
rect 4897 1857 4903 1865
rect 3323 1829 4903 1857
rect 3323 1822 3329 1829
rect 4897 1822 4903 1829
rect 3271 1811 3323 1817
rect 6535 1869 6587 1875
rect 4955 1857 4961 1865
rect 6529 1857 6535 1865
rect 4955 1829 6535 1857
rect 4955 1822 4961 1829
rect 6529 1822 6535 1829
rect 4903 1811 4955 1817
rect 8167 1869 8219 1875
rect 6587 1857 6593 1865
rect 8161 1857 8167 1865
rect 6587 1829 8167 1857
rect 6587 1822 6593 1829
rect 8161 1822 8167 1829
rect 6535 1811 6587 1817
rect 9799 1869 9851 1875
rect 8219 1857 8225 1865
rect 9793 1857 9799 1865
rect 8219 1829 9799 1857
rect 8219 1822 8225 1829
rect 9793 1822 9799 1829
rect 8167 1811 8219 1817
rect 11431 1869 11483 1875
rect 9851 1857 9857 1865
rect 11425 1857 11431 1865
rect 9851 1829 11431 1857
rect 9851 1822 9857 1829
rect 11425 1822 11431 1829
rect 9799 1811 9851 1817
rect 13063 1869 13115 1875
rect 11483 1857 11489 1865
rect 13057 1857 13063 1865
rect 11483 1829 13063 1857
rect 11483 1822 11489 1829
rect 13057 1822 13063 1829
rect 11431 1811 11483 1817
rect 13115 1822 13121 1865
rect 13063 1811 13115 1817
rect 7 1665 59 1671
rect 1 1618 7 1661
rect 1639 1665 1691 1671
rect 59 1653 65 1661
rect 1633 1653 1639 1661
rect 59 1625 1639 1653
rect 59 1618 65 1625
rect 1633 1618 1639 1625
rect 7 1607 59 1613
rect 3271 1665 3323 1671
rect 1691 1653 1697 1661
rect 3265 1653 3271 1661
rect 1691 1625 3271 1653
rect 1691 1618 1697 1625
rect 3265 1618 3271 1625
rect 1639 1607 1691 1613
rect 4903 1665 4955 1671
rect 3323 1653 3329 1661
rect 4897 1653 4903 1661
rect 3323 1625 4903 1653
rect 3323 1618 3329 1625
rect 4897 1618 4903 1625
rect 3271 1607 3323 1613
rect 6535 1665 6587 1671
rect 4955 1653 4961 1661
rect 6529 1653 6535 1661
rect 4955 1625 6535 1653
rect 4955 1618 4961 1625
rect 6529 1618 6535 1625
rect 4903 1607 4955 1613
rect 8167 1665 8219 1671
rect 6587 1653 6593 1661
rect 8161 1653 8167 1661
rect 6587 1625 8167 1653
rect 6587 1618 6593 1625
rect 8161 1618 8167 1625
rect 6535 1607 6587 1613
rect 9799 1665 9851 1671
rect 8219 1653 8225 1661
rect 9793 1653 9799 1661
rect 8219 1625 9799 1653
rect 8219 1618 8225 1625
rect 9793 1618 9799 1625
rect 8167 1607 8219 1613
rect 11431 1665 11483 1671
rect 9851 1653 9857 1661
rect 11425 1653 11431 1661
rect 9851 1625 11431 1653
rect 9851 1618 9857 1625
rect 11425 1618 11431 1625
rect 9799 1607 9851 1613
rect 13063 1665 13115 1671
rect 11483 1653 11489 1661
rect 13057 1653 13063 1661
rect 11483 1625 13063 1653
rect 11483 1618 11489 1625
rect 13057 1618 13063 1625
rect 11431 1607 11483 1613
rect 13115 1618 13121 1661
rect 13063 1607 13115 1613
rect 7 1461 59 1467
rect 1 1414 7 1457
rect 1639 1461 1691 1467
rect 59 1449 65 1457
rect 1633 1449 1639 1457
rect 59 1421 1639 1449
rect 59 1414 65 1421
rect 1633 1414 1639 1421
rect 7 1403 59 1409
rect 3271 1461 3323 1467
rect 1691 1449 1697 1457
rect 3265 1449 3271 1457
rect 1691 1421 3271 1449
rect 1691 1414 1697 1421
rect 3265 1414 3271 1421
rect 1639 1403 1691 1409
rect 4903 1461 4955 1467
rect 3323 1449 3329 1457
rect 4897 1449 4903 1457
rect 3323 1421 4903 1449
rect 3323 1414 3329 1421
rect 4897 1414 4903 1421
rect 3271 1403 3323 1409
rect 6535 1461 6587 1467
rect 4955 1449 4961 1457
rect 6529 1449 6535 1457
rect 4955 1421 6535 1449
rect 4955 1414 4961 1421
rect 6529 1414 6535 1421
rect 4903 1403 4955 1409
rect 8167 1461 8219 1467
rect 6587 1449 6593 1457
rect 8161 1449 8167 1457
rect 6587 1421 8167 1449
rect 6587 1414 6593 1421
rect 8161 1414 8167 1421
rect 6535 1403 6587 1409
rect 9799 1461 9851 1467
rect 8219 1449 8225 1457
rect 9793 1449 9799 1457
rect 8219 1421 9799 1449
rect 8219 1414 8225 1421
rect 9793 1414 9799 1421
rect 8167 1403 8219 1409
rect 11431 1461 11483 1467
rect 9851 1449 9857 1457
rect 11425 1449 11431 1457
rect 9851 1421 11431 1449
rect 9851 1414 9857 1421
rect 11425 1414 11431 1421
rect 9799 1403 9851 1409
rect 13063 1461 13115 1467
rect 11483 1449 11489 1457
rect 13057 1449 13063 1457
rect 11483 1421 13063 1449
rect 11483 1414 11489 1421
rect 13057 1414 13063 1421
rect 11431 1403 11483 1409
rect 13115 1414 13121 1457
rect 13063 1403 13115 1409
rect 7 1257 59 1263
rect 1 1210 7 1253
rect 1639 1257 1691 1263
rect 59 1245 65 1253
rect 1633 1245 1639 1253
rect 59 1217 1639 1245
rect 59 1210 65 1217
rect 1633 1210 1639 1217
rect 7 1199 59 1205
rect 3271 1257 3323 1263
rect 1691 1245 1697 1253
rect 3265 1245 3271 1253
rect 1691 1217 3271 1245
rect 1691 1210 1697 1217
rect 3265 1210 3271 1217
rect 1639 1199 1691 1205
rect 4903 1257 4955 1263
rect 3323 1245 3329 1253
rect 4897 1245 4903 1253
rect 3323 1217 4903 1245
rect 3323 1210 3329 1217
rect 4897 1210 4903 1217
rect 3271 1199 3323 1205
rect 6535 1257 6587 1263
rect 4955 1245 4961 1253
rect 6529 1245 6535 1253
rect 4955 1217 6535 1245
rect 4955 1210 4961 1217
rect 6529 1210 6535 1217
rect 4903 1199 4955 1205
rect 8167 1257 8219 1263
rect 6587 1245 6593 1253
rect 8161 1245 8167 1253
rect 6587 1217 8167 1245
rect 6587 1210 6593 1217
rect 8161 1210 8167 1217
rect 6535 1199 6587 1205
rect 9799 1257 9851 1263
rect 8219 1245 8225 1253
rect 9793 1245 9799 1253
rect 8219 1217 9799 1245
rect 8219 1210 8225 1217
rect 9793 1210 9799 1217
rect 8167 1199 8219 1205
rect 11431 1257 11483 1263
rect 9851 1245 9857 1253
rect 11425 1245 11431 1253
rect 9851 1217 11431 1245
rect 9851 1210 9857 1217
rect 11425 1210 11431 1217
rect 9799 1199 9851 1205
rect 13063 1257 13115 1263
rect 11483 1245 11489 1253
rect 13057 1245 13063 1253
rect 11483 1217 13063 1245
rect 11483 1210 11489 1217
rect 13057 1210 13063 1217
rect 11431 1199 11483 1205
rect 13115 1210 13121 1253
rect 13063 1199 13115 1205
rect 7 1053 59 1059
rect 1 1006 7 1049
rect 1639 1053 1691 1059
rect 59 1041 65 1049
rect 1633 1041 1639 1049
rect 59 1013 1639 1041
rect 59 1006 65 1013
rect 1633 1006 1639 1013
rect 7 995 59 1001
rect 3271 1053 3323 1059
rect 1691 1041 1697 1049
rect 3265 1041 3271 1049
rect 1691 1013 3271 1041
rect 1691 1006 1697 1013
rect 3265 1006 3271 1013
rect 1639 995 1691 1001
rect 4903 1053 4955 1059
rect 3323 1041 3329 1049
rect 4897 1041 4903 1049
rect 3323 1013 4903 1041
rect 3323 1006 3329 1013
rect 4897 1006 4903 1013
rect 3271 995 3323 1001
rect 6535 1053 6587 1059
rect 4955 1041 4961 1049
rect 6529 1041 6535 1049
rect 4955 1013 6535 1041
rect 4955 1006 4961 1013
rect 6529 1006 6535 1013
rect 4903 995 4955 1001
rect 8167 1053 8219 1059
rect 6587 1041 6593 1049
rect 8161 1041 8167 1049
rect 6587 1013 8167 1041
rect 6587 1006 6593 1013
rect 8161 1006 8167 1013
rect 6535 995 6587 1001
rect 9799 1053 9851 1059
rect 8219 1041 8225 1049
rect 9793 1041 9799 1049
rect 8219 1013 9799 1041
rect 8219 1006 8225 1013
rect 9793 1006 9799 1013
rect 8167 995 8219 1001
rect 11431 1053 11483 1059
rect 9851 1041 9857 1049
rect 11425 1041 11431 1049
rect 9851 1013 11431 1041
rect 9851 1006 9857 1013
rect 11425 1006 11431 1013
rect 9799 995 9851 1001
rect 13063 1053 13115 1059
rect 11483 1041 11489 1049
rect 13057 1041 13063 1049
rect 11483 1013 13063 1041
rect 11483 1006 11489 1013
rect 13057 1006 13063 1013
rect 11431 995 11483 1001
rect 13115 1006 13121 1049
rect 13063 995 13115 1001
rect 212 847 218 899
rect 270 887 276 899
rect 416 887 422 899
rect 270 859 422 887
rect 270 847 276 859
rect 416 847 422 859
rect 474 887 480 899
rect 620 887 626 899
rect 474 859 626 887
rect 474 847 480 859
rect 620 847 626 859
rect 678 887 684 899
rect 824 887 830 899
rect 678 859 830 887
rect 678 847 684 859
rect 824 847 830 859
rect 882 887 888 899
rect 1028 887 1034 899
rect 882 859 1034 887
rect 882 847 888 859
rect 1028 847 1034 859
rect 1086 887 1092 899
rect 1232 887 1238 899
rect 1086 859 1238 887
rect 1086 847 1092 859
rect 1232 847 1238 859
rect 1290 887 1296 899
rect 1436 887 1442 899
rect 1290 859 1442 887
rect 1290 847 1296 859
rect 1436 847 1442 859
rect 1494 887 1500 899
rect 1640 887 1646 899
rect 1494 859 1646 887
rect 1494 847 1500 859
rect 1640 847 1646 859
rect 1698 887 1704 899
rect 1844 887 1850 899
rect 1698 859 1850 887
rect 1698 847 1704 859
rect 1844 847 1850 859
rect 1902 887 1908 899
rect 2048 887 2054 899
rect 1902 859 2054 887
rect 1902 847 1908 859
rect 2048 847 2054 859
rect 2106 887 2112 899
rect 2252 887 2258 899
rect 2106 859 2258 887
rect 2106 847 2112 859
rect 2252 847 2258 859
rect 2310 887 2316 899
rect 2456 887 2462 899
rect 2310 859 2462 887
rect 2310 847 2316 859
rect 2456 847 2462 859
rect 2514 887 2520 899
rect 2660 887 2666 899
rect 2514 859 2666 887
rect 2514 847 2520 859
rect 2660 847 2666 859
rect 2718 887 2724 899
rect 2864 887 2870 899
rect 2718 859 2870 887
rect 2718 847 2724 859
rect 2864 847 2870 859
rect 2922 887 2928 899
rect 3068 887 3074 899
rect 2922 859 3074 887
rect 2922 847 2928 859
rect 3068 847 3074 859
rect 3126 887 3132 899
rect 3272 887 3278 899
rect 3126 859 3278 887
rect 3126 847 3132 859
rect 3272 847 3278 859
rect 3330 887 3336 899
rect 3476 887 3482 899
rect 3330 859 3482 887
rect 3330 847 3336 859
rect 3476 847 3482 859
rect 3534 887 3540 899
rect 3680 887 3686 899
rect 3534 859 3686 887
rect 3534 847 3540 859
rect 3680 847 3686 859
rect 3738 887 3744 899
rect 3884 887 3890 899
rect 3738 859 3890 887
rect 3738 847 3744 859
rect 3884 847 3890 859
rect 3942 887 3948 899
rect 4088 887 4094 899
rect 3942 859 4094 887
rect 3942 847 3948 859
rect 4088 847 4094 859
rect 4146 887 4152 899
rect 4292 887 4298 899
rect 4146 859 4298 887
rect 4146 847 4152 859
rect 4292 847 4298 859
rect 4350 887 4356 899
rect 4496 887 4502 899
rect 4350 859 4502 887
rect 4350 847 4356 859
rect 4496 847 4502 859
rect 4554 887 4560 899
rect 4700 887 4706 899
rect 4554 859 4706 887
rect 4554 847 4560 859
rect 4700 847 4706 859
rect 4758 887 4764 899
rect 4904 887 4910 899
rect 4758 859 4910 887
rect 4758 847 4764 859
rect 4904 847 4910 859
rect 4962 887 4968 899
rect 5108 887 5114 899
rect 4962 859 5114 887
rect 4962 847 4968 859
rect 5108 847 5114 859
rect 5166 887 5172 899
rect 5312 887 5318 899
rect 5166 859 5318 887
rect 5166 847 5172 859
rect 5312 847 5318 859
rect 5370 887 5376 899
rect 5516 887 5522 899
rect 5370 859 5522 887
rect 5370 847 5376 859
rect 5516 847 5522 859
rect 5574 887 5580 899
rect 5720 887 5726 899
rect 5574 859 5726 887
rect 5574 847 5580 859
rect 5720 847 5726 859
rect 5778 887 5784 899
rect 5924 887 5930 899
rect 5778 859 5930 887
rect 5778 847 5784 859
rect 5924 847 5930 859
rect 5982 887 5988 899
rect 6128 887 6134 899
rect 5982 859 6134 887
rect 5982 847 5988 859
rect 6128 847 6134 859
rect 6186 887 6192 899
rect 6332 887 6338 899
rect 6186 859 6338 887
rect 6186 847 6192 859
rect 6332 847 6338 859
rect 6390 887 6396 899
rect 6536 887 6542 899
rect 6390 859 6542 887
rect 6390 847 6396 859
rect 6536 847 6542 859
rect 6594 887 6600 899
rect 6740 887 6746 899
rect 6594 859 6746 887
rect 6594 847 6600 859
rect 6740 847 6746 859
rect 6798 887 6804 899
rect 6944 887 6950 899
rect 6798 859 6950 887
rect 6798 847 6804 859
rect 6944 847 6950 859
rect 7002 887 7008 899
rect 7148 887 7154 899
rect 7002 859 7154 887
rect 7002 847 7008 859
rect 7148 847 7154 859
rect 7206 887 7212 899
rect 7352 887 7358 899
rect 7206 859 7358 887
rect 7206 847 7212 859
rect 7352 847 7358 859
rect 7410 887 7416 899
rect 7556 887 7562 899
rect 7410 859 7562 887
rect 7410 847 7416 859
rect 7556 847 7562 859
rect 7614 887 7620 899
rect 7760 887 7766 899
rect 7614 859 7766 887
rect 7614 847 7620 859
rect 7760 847 7766 859
rect 7818 887 7824 899
rect 7964 887 7970 899
rect 7818 859 7970 887
rect 7818 847 7824 859
rect 7964 847 7970 859
rect 8022 887 8028 899
rect 8168 887 8174 899
rect 8022 859 8174 887
rect 8022 847 8028 859
rect 8168 847 8174 859
rect 8226 887 8232 899
rect 8372 887 8378 899
rect 8226 859 8378 887
rect 8226 847 8232 859
rect 8372 847 8378 859
rect 8430 887 8436 899
rect 8576 887 8582 899
rect 8430 859 8582 887
rect 8430 847 8436 859
rect 8576 847 8582 859
rect 8634 887 8640 899
rect 8780 887 8786 899
rect 8634 859 8786 887
rect 8634 847 8640 859
rect 8780 847 8786 859
rect 8838 887 8844 899
rect 8984 887 8990 899
rect 8838 859 8990 887
rect 8838 847 8844 859
rect 8984 847 8990 859
rect 9042 887 9048 899
rect 9188 887 9194 899
rect 9042 859 9194 887
rect 9042 847 9048 859
rect 9188 847 9194 859
rect 9246 887 9252 899
rect 9392 887 9398 899
rect 9246 859 9398 887
rect 9246 847 9252 859
rect 9392 847 9398 859
rect 9450 887 9456 899
rect 9596 887 9602 899
rect 9450 859 9602 887
rect 9450 847 9456 859
rect 9596 847 9602 859
rect 9654 887 9660 899
rect 9800 887 9806 899
rect 9654 859 9806 887
rect 9654 847 9660 859
rect 9800 847 9806 859
rect 9858 887 9864 899
rect 10004 887 10010 899
rect 9858 859 10010 887
rect 9858 847 9864 859
rect 10004 847 10010 859
rect 10062 887 10068 899
rect 10208 887 10214 899
rect 10062 859 10214 887
rect 10062 847 10068 859
rect 10208 847 10214 859
rect 10266 887 10272 899
rect 10412 887 10418 899
rect 10266 859 10418 887
rect 10266 847 10272 859
rect 10412 847 10418 859
rect 10470 887 10476 899
rect 10616 887 10622 899
rect 10470 859 10622 887
rect 10470 847 10476 859
rect 10616 847 10622 859
rect 10674 887 10680 899
rect 10820 887 10826 899
rect 10674 859 10826 887
rect 10674 847 10680 859
rect 10820 847 10826 859
rect 10878 887 10884 899
rect 11024 887 11030 899
rect 10878 859 11030 887
rect 10878 847 10884 859
rect 11024 847 11030 859
rect 11082 887 11088 899
rect 11228 887 11234 899
rect 11082 859 11234 887
rect 11082 847 11088 859
rect 11228 847 11234 859
rect 11286 887 11292 899
rect 11432 887 11438 899
rect 11286 859 11438 887
rect 11286 847 11292 859
rect 11432 847 11438 859
rect 11490 887 11496 899
rect 11636 887 11642 899
rect 11490 859 11642 887
rect 11490 847 11496 859
rect 11636 847 11642 859
rect 11694 887 11700 899
rect 11840 887 11846 899
rect 11694 859 11846 887
rect 11694 847 11700 859
rect 11840 847 11846 859
rect 11898 887 11904 899
rect 12044 887 12050 899
rect 11898 859 12050 887
rect 11898 847 11904 859
rect 12044 847 12050 859
rect 12102 887 12108 899
rect 12248 887 12254 899
rect 12102 859 12254 887
rect 12102 847 12108 859
rect 12248 847 12254 859
rect 12306 887 12312 899
rect 12452 887 12458 899
rect 12306 859 12458 887
rect 12306 847 12312 859
rect 12452 847 12458 859
rect 12510 887 12516 899
rect 12656 887 12662 899
rect 12510 859 12662 887
rect 12510 847 12516 859
rect 12656 847 12662 859
rect 12714 887 12720 899
rect 12860 887 12866 899
rect 12714 859 12866 887
rect 12714 847 12720 859
rect 12860 847 12866 859
rect 12918 887 12924 899
rect 13078 887 13084 899
rect 12918 859 13084 887
rect 12918 847 12924 859
rect 13078 847 13084 859
rect 13136 847 13142 899
rect 61 368 89 396
rect 12 -32 40 32
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_0
timestamp 1581320205
transform 1 0 12852 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1
timestamp 1581320205
transform 1 0 12648 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_2
timestamp 1581320205
transform 1 0 12444 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_3
timestamp 1581320205
transform 1 0 12240 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_4
timestamp 1581320205
transform 1 0 12036 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_5
timestamp 1581320205
transform 1 0 11832 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_6
timestamp 1581320205
transform 1 0 11628 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_7
timestamp 1581320205
transform 1 0 11424 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_8
timestamp 1581320205
transform 1 0 11220 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_9
timestamp 1581320205
transform 1 0 11016 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_10
timestamp 1581320205
transform 1 0 10812 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_11
timestamp 1581320205
transform 1 0 10608 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_12
timestamp 1581320205
transform 1 0 10404 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_13
timestamp 1581320205
transform 1 0 10200 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_14
timestamp 1581320205
transform 1 0 9996 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_15
timestamp 1581320205
transform 1 0 9792 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_16
timestamp 1581320205
transform 1 0 9588 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_17
timestamp 1581320205
transform 1 0 9384 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_18
timestamp 1581320205
transform 1 0 9180 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_19
timestamp 1581320205
transform 1 0 8976 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_20
timestamp 1581320205
transform 1 0 8772 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_21
timestamp 1581320205
transform 1 0 8568 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_22
timestamp 1581320205
transform 1 0 8364 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_23
timestamp 1581320205
transform 1 0 8160 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_24
timestamp 1581320205
transform 1 0 7956 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_25
timestamp 1581320205
transform 1 0 7752 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_26
timestamp 1581320205
transform 1 0 7548 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_27
timestamp 1581320205
transform 1 0 7344 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_28
timestamp 1581320205
transform 1 0 7140 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_29
timestamp 1581320205
transform 1 0 6936 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_30
timestamp 1581320205
transform 1 0 6732 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_31
timestamp 1581320205
transform 1 0 6528 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_32
timestamp 1581320205
transform 1 0 6324 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_33
timestamp 1581320205
transform 1 0 6120 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_34
timestamp 1581320205
transform 1 0 5916 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_35
timestamp 1581320205
transform 1 0 5712 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_36
timestamp 1581320205
transform 1 0 5508 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_37
timestamp 1581320205
transform 1 0 5304 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_38
timestamp 1581320205
transform 1 0 5100 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_39
timestamp 1581320205
transform 1 0 4896 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_40
timestamp 1581320205
transform 1 0 4692 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_41
timestamp 1581320205
transform 1 0 4488 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_42
timestamp 1581320205
transform 1 0 4284 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_43
timestamp 1581320205
transform 1 0 4080 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_44
timestamp 1581320205
transform 1 0 3876 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_45
timestamp 1581320205
transform 1 0 3672 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_46
timestamp 1581320205
transform 1 0 3468 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_47
timestamp 1581320205
transform 1 0 3264 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_48
timestamp 1581320205
transform 1 0 3060 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_49
timestamp 1581320205
transform 1 0 2856 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_50
timestamp 1581320205
transform 1 0 2652 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_51
timestamp 1581320205
transform 1 0 2448 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_52
timestamp 1581320205
transform 1 0 2244 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_53
timestamp 1581320205
transform 1 0 2040 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_54
timestamp 1581320205
transform 1 0 1836 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_55
timestamp 1581320205
transform 1 0 1632 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_56
timestamp 1581320205
transform 1 0 1428 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_57
timestamp 1581320205
transform 1 0 1224 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_58
timestamp 1581320205
transform 1 0 1020 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_59
timestamp 1581320205
transform 1 0 816 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_60
timestamp 1581320205
transform 1 0 612 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_61
timestamp 1581320205
transform 1 0 408 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_62
timestamp 1581320205
transform 1 0 204 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_63
timestamp 1581320205
transform 1 0 0 0 1 7817
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_64
timestamp 1581320205
transform 1 0 12444 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_65
timestamp 1581320205
transform 1 0 12036 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_66
timestamp 1581320205
transform 1 0 11832 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_67
timestamp 1581320205
transform 1 0 11628 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_68
timestamp 1581320205
transform 1 0 11220 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_69
timestamp 1581320205
transform 1 0 10608 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_70
timestamp 1581320205
transform 1 0 10404 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_71
timestamp 1581320205
transform 1 0 10200 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_72
timestamp 1581320205
transform 1 0 9792 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_73
timestamp 1581320205
transform 1 0 8976 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_74
timestamp 1581320205
transform 1 0 8772 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_75
timestamp 1581320205
transform 1 0 8160 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_76
timestamp 1581320205
transform 1 0 7752 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_77
timestamp 1581320205
transform 1 0 6732 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_78
timestamp 1581320205
transform 1 0 6528 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_79
timestamp 1581320205
transform 1 0 6324 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_80
timestamp 1581320205
transform 1 0 6120 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_81
timestamp 1581320205
transform 1 0 5916 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_82
timestamp 1581320205
transform 1 0 5508 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_83
timestamp 1581320205
transform 1 0 5100 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_84
timestamp 1581320205
transform 1 0 4896 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_85
timestamp 1581320205
transform 1 0 4692 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_86
timestamp 1581320205
transform 1 0 4488 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_87
timestamp 1581320205
transform 1 0 4284 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_88
timestamp 1581320205
transform 1 0 3876 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_89
timestamp 1581320205
transform 1 0 3672 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_90
timestamp 1581320205
transform 1 0 3468 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_91
timestamp 1581320205
transform 1 0 3264 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_92
timestamp 1581320205
transform 1 0 3060 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_93
timestamp 1581320205
transform 1 0 2856 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_94
timestamp 1581320205
transform 1 0 2652 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_95
timestamp 1581320205
transform 1 0 2448 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_96
timestamp 1581320205
transform 1 0 2244 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_97
timestamp 1581320205
transform 1 0 1836 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_98
timestamp 1581320205
transform 1 0 1428 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_99
timestamp 1581320205
transform 1 0 816 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_100
timestamp 1581320205
transform 1 0 612 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_101
timestamp 1581320205
transform 1 0 408 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_102
timestamp 1581320205
transform 1 0 204 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_103
timestamp 1581320205
transform 1 0 0 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_104
timestamp 1581320205
transform 1 0 12852 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_105
timestamp 1581320205
transform 1 0 11832 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_106
timestamp 1581320205
transform 1 0 11220 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_107
timestamp 1581320205
transform 1 0 10404 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_108
timestamp 1581320205
transform 1 0 10200 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_109
timestamp 1581320205
transform 1 0 9996 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_110
timestamp 1581320205
transform 1 0 9384 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_111
timestamp 1581320205
transform 1 0 8976 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_112
timestamp 1581320205
transform 1 0 8568 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_113
timestamp 1581320205
transform 1 0 8364 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_114
timestamp 1581320205
transform 1 0 7956 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_115
timestamp 1581320205
transform 1 0 7752 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_116
timestamp 1581320205
transform 1 0 7140 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_117
timestamp 1581320205
transform 1 0 6936 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_118
timestamp 1581320205
transform 1 0 6732 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_119
timestamp 1581320205
transform 1 0 5916 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_120
timestamp 1581320205
transform 1 0 5508 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_121
timestamp 1581320205
transform 1 0 5304 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_122
timestamp 1581320205
transform 1 0 5100 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_123
timestamp 1581320205
transform 1 0 4896 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_124
timestamp 1581320205
transform 1 0 4692 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_125
timestamp 1581320205
transform 1 0 4488 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_126
timestamp 1581320205
transform 1 0 4080 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_127
timestamp 1581320205
transform 1 0 3876 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_128
timestamp 1581320205
transform 1 0 3672 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_129
timestamp 1581320205
transform 1 0 3468 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_130
timestamp 1581320205
transform 1 0 3060 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_131
timestamp 1581320205
transform 1 0 2856 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_132
timestamp 1581320205
transform 1 0 2652 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_133
timestamp 1581320205
transform 1 0 2244 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_134
timestamp 1581320205
transform 1 0 2040 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_135
timestamp 1581320205
transform 1 0 1428 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_136
timestamp 1581320205
transform 1 0 816 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_137
timestamp 1581320205
transform 1 0 612 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_138
timestamp 1581320205
transform 1 0 408 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_139
timestamp 1581320205
transform 1 0 204 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_140
timestamp 1581320205
transform 1 0 0 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_141
timestamp 1581320205
transform 1 0 12444 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_142
timestamp 1581320205
transform 1 0 11016 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_143
timestamp 1581320205
transform 1 0 10812 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_144
timestamp 1581320205
transform 1 0 9180 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_145
timestamp 1581320205
transform 1 0 8976 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_146
timestamp 1581320205
transform 1 0 8772 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_147
timestamp 1581320205
transform 1 0 8160 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_148
timestamp 1581320205
transform 1 0 7956 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_149
timestamp 1581320205
transform 1 0 7344 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_150
timestamp 1581320205
transform 1 0 6936 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_151
timestamp 1581320205
transform 1 0 6732 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_152
timestamp 1581320205
transform 1 0 5508 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_153
timestamp 1581320205
transform 1 0 5304 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_154
timestamp 1581320205
transform 1 0 3672 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_155
timestamp 1581320205
transform 1 0 2652 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_156
timestamp 1581320205
transform 1 0 2040 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_157
timestamp 1581320205
transform 1 0 1836 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_158
timestamp 1581320205
transform 1 0 1020 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_159
timestamp 1581320205
transform 1 0 816 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_160
timestamp 1581320205
transform 1 0 204 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_161
timestamp 1581320205
transform 1 0 0 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_162
timestamp 1581320205
transform 1 0 12852 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_163
timestamp 1581320205
transform 1 0 12648 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_164
timestamp 1581320205
transform 1 0 12444 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_165
timestamp 1581320205
transform 1 0 11628 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_166
timestamp 1581320205
transform 1 0 11220 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_167
timestamp 1581320205
transform 1 0 11016 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_168
timestamp 1581320205
transform 1 0 10404 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_169
timestamp 1581320205
transform 1 0 10200 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_170
timestamp 1581320205
transform 1 0 9996 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_171
timestamp 1581320205
transform 1 0 9588 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_172
timestamp 1581320205
transform 1 0 9180 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_173
timestamp 1581320205
transform 1 0 8772 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_174
timestamp 1581320205
transform 1 0 8364 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_175
timestamp 1581320205
transform 1 0 8160 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_176
timestamp 1581320205
transform 1 0 7956 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_177
timestamp 1581320205
transform 1 0 7344 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_178
timestamp 1581320205
transform 1 0 7140 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_179
timestamp 1581320205
transform 1 0 6732 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_180
timestamp 1581320205
transform 1 0 5712 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_181
timestamp 1581320205
transform 1 0 4896 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_182
timestamp 1581320205
transform 1 0 4692 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_183
timestamp 1581320205
transform 1 0 4488 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_184
timestamp 1581320205
transform 1 0 4284 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_185
timestamp 1581320205
transform 1 0 4080 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_186
timestamp 1581320205
transform 1 0 3876 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_187
timestamp 1581320205
transform 1 0 3264 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_188
timestamp 1581320205
transform 1 0 3060 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_189
timestamp 1581320205
transform 1 0 2856 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_190
timestamp 1581320205
transform 1 0 2448 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_191
timestamp 1581320205
transform 1 0 2244 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_192
timestamp 1581320205
transform 1 0 1632 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_193
timestamp 1581320205
transform 1 0 1020 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_194
timestamp 1581320205
transform 1 0 612 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_195
timestamp 1581320205
transform 1 0 408 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_196
timestamp 1581320205
transform 1 0 204 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_197
timestamp 1581320205
transform 1 0 12852 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_198
timestamp 1581320205
transform 1 0 12648 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_199
timestamp 1581320205
transform 1 0 12036 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_200
timestamp 1581320205
transform 1 0 11424 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_201
timestamp 1581320205
transform 1 0 11220 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_202
timestamp 1581320205
transform 1 0 11016 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_203
timestamp 1581320205
transform 1 0 10812 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_204
timestamp 1581320205
transform 1 0 10404 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_205
timestamp 1581320205
transform 1 0 10200 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_206
timestamp 1581320205
transform 1 0 9792 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_207
timestamp 1581320205
transform 1 0 9384 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_208
timestamp 1581320205
transform 1 0 9180 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_209
timestamp 1581320205
transform 1 0 8772 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_210
timestamp 1581320205
transform 1 0 8364 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_211
timestamp 1581320205
transform 1 0 7752 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_212
timestamp 1581320205
transform 1 0 7548 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_213
timestamp 1581320205
transform 1 0 7344 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_214
timestamp 1581320205
transform 1 0 7140 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_215
timestamp 1581320205
transform 1 0 6936 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_216
timestamp 1581320205
transform 1 0 6732 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_217
timestamp 1581320205
transform 1 0 6528 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_218
timestamp 1581320205
transform 1 0 6324 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_219
timestamp 1581320205
transform 1 0 5100 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_220
timestamp 1581320205
transform 1 0 4896 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_221
timestamp 1581320205
transform 1 0 4692 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_222
timestamp 1581320205
transform 1 0 4488 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_223
timestamp 1581320205
transform 1 0 4284 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_224
timestamp 1581320205
transform 1 0 4080 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_225
timestamp 1581320205
transform 1 0 3060 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_226
timestamp 1581320205
transform 1 0 2856 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_227
timestamp 1581320205
transform 1 0 2448 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_228
timestamp 1581320205
transform 1 0 2244 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_229
timestamp 1581320205
transform 1 0 2040 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_230
timestamp 1581320205
transform 1 0 1632 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_231
timestamp 1581320205
transform 1 0 1428 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_232
timestamp 1581320205
transform 1 0 408 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_233
timestamp 1581320205
transform 1 0 204 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_234
timestamp 1581320205
transform 1 0 12036 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_235
timestamp 1581320205
transform 1 0 11424 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_236
timestamp 1581320205
transform 1 0 11220 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_237
timestamp 1581320205
transform 1 0 11016 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_238
timestamp 1581320205
transform 1 0 10608 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_239
timestamp 1581320205
transform 1 0 10404 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_240
timestamp 1581320205
transform 1 0 8976 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_241
timestamp 1581320205
transform 1 0 8568 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_242
timestamp 1581320205
transform 1 0 8364 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_243
timestamp 1581320205
transform 1 0 7956 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_244
timestamp 1581320205
transform 1 0 7752 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_245
timestamp 1581320205
transform 1 0 7548 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_246
timestamp 1581320205
transform 1 0 7344 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_247
timestamp 1581320205
transform 1 0 6936 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_248
timestamp 1581320205
transform 1 0 6732 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_249
timestamp 1581320205
transform 1 0 6528 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_250
timestamp 1581320205
transform 1 0 5916 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_251
timestamp 1581320205
transform 1 0 5508 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_252
timestamp 1581320205
transform 1 0 5100 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_253
timestamp 1581320205
transform 1 0 4896 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_254
timestamp 1581320205
transform 1 0 4488 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_255
timestamp 1581320205
transform 1 0 3876 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_256
timestamp 1581320205
transform 1 0 3264 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_257
timestamp 1581320205
transform 1 0 3060 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_258
timestamp 1581320205
transform 1 0 2652 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_259
timestamp 1581320205
transform 1 0 2448 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_260
timestamp 1581320205
transform 1 0 1224 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_261
timestamp 1581320205
transform 1 0 1020 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_262
timestamp 1581320205
transform 1 0 612 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_263
timestamp 1581320205
transform 1 0 12852 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_264
timestamp 1581320205
transform 1 0 11832 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_265
timestamp 1581320205
transform 1 0 11424 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_266
timestamp 1581320205
transform 1 0 10200 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_267
timestamp 1581320205
transform 1 0 9792 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_268
timestamp 1581320205
transform 1 0 9588 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_269
timestamp 1581320205
transform 1 0 9384 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_270
timestamp 1581320205
transform 1 0 8976 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_271
timestamp 1581320205
transform 1 0 8772 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_272
timestamp 1581320205
transform 1 0 8568 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_273
timestamp 1581320205
transform 1 0 8160 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_274
timestamp 1581320205
transform 1 0 7752 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_275
timestamp 1581320205
transform 1 0 7140 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_276
timestamp 1581320205
transform 1 0 6732 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_277
timestamp 1581320205
transform 1 0 6324 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_278
timestamp 1581320205
transform 1 0 6120 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_279
timestamp 1581320205
transform 1 0 5916 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_280
timestamp 1581320205
transform 1 0 5712 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_281
timestamp 1581320205
transform 1 0 5304 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_282
timestamp 1581320205
transform 1 0 4692 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_283
timestamp 1581320205
transform 1 0 4488 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_284
timestamp 1581320205
transform 1 0 4284 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_285
timestamp 1581320205
transform 1 0 4080 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_286
timestamp 1581320205
transform 1 0 3672 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_287
timestamp 1581320205
transform 1 0 3264 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_288
timestamp 1581320205
transform 1 0 2244 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_289
timestamp 1581320205
transform 1 0 2040 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_290
timestamp 1581320205
transform 1 0 1836 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_291
timestamp 1581320205
transform 1 0 1428 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_292
timestamp 1581320205
transform 1 0 1224 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_293
timestamp 1581320205
transform 1 0 1020 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_294
timestamp 1581320205
transform 1 0 12444 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_295
timestamp 1581320205
transform 1 0 11832 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_296
timestamp 1581320205
transform 1 0 11424 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_297
timestamp 1581320205
transform 1 0 10812 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_298
timestamp 1581320205
transform 1 0 10608 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_299
timestamp 1581320205
transform 1 0 10404 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_300
timestamp 1581320205
transform 1 0 9384 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_301
timestamp 1581320205
transform 1 0 9180 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_302
timestamp 1581320205
transform 1 0 8976 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_303
timestamp 1581320205
transform 1 0 8772 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_304
timestamp 1581320205
transform 1 0 8364 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_305
timestamp 1581320205
transform 1 0 7956 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_306
timestamp 1581320205
transform 1 0 7752 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_307
timestamp 1581320205
transform 1 0 7344 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_308
timestamp 1581320205
transform 1 0 6528 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_309
timestamp 1581320205
transform 1 0 5916 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_310
timestamp 1581320205
transform 1 0 5712 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_311
timestamp 1581320205
transform 1 0 5508 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_312
timestamp 1581320205
transform 1 0 4896 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_313
timestamp 1581320205
transform 1 0 4488 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_314
timestamp 1581320205
transform 1 0 4284 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_315
timestamp 1581320205
transform 1 0 3468 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_316
timestamp 1581320205
transform 1 0 2856 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_317
timestamp 1581320205
transform 1 0 2040 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_318
timestamp 1581320205
transform 1 0 408 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_319
timestamp 1581320205
transform 1 0 204 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_320
timestamp 1581320205
transform 1 0 12036 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_321
timestamp 1581320205
transform 1 0 11832 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_322
timestamp 1581320205
transform 1 0 10812 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_323
timestamp 1581320205
transform 1 0 9996 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_324
timestamp 1581320205
transform 1 0 8772 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_325
timestamp 1581320205
transform 1 0 8568 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_326
timestamp 1581320205
transform 1 0 8364 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_327
timestamp 1581320205
transform 1 0 8160 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_328
timestamp 1581320205
transform 1 0 7548 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_329
timestamp 1581320205
transform 1 0 6732 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_330
timestamp 1581320205
transform 1 0 6324 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_331
timestamp 1581320205
transform 1 0 5712 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_332
timestamp 1581320205
transform 1 0 5304 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_333
timestamp 1581320205
transform 1 0 4896 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_334
timestamp 1581320205
transform 1 0 4692 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_335
timestamp 1581320205
transform 1 0 4488 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_336
timestamp 1581320205
transform 1 0 4284 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_337
timestamp 1581320205
transform 1 0 3672 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_338
timestamp 1581320205
transform 1 0 3264 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_339
timestamp 1581320205
transform 1 0 3060 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_340
timestamp 1581320205
transform 1 0 2652 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_341
timestamp 1581320205
transform 1 0 1632 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_342
timestamp 1581320205
transform 1 0 1224 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_343
timestamp 1581320205
transform 1 0 612 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_344
timestamp 1581320205
transform 1 0 0 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_345
timestamp 1581320205
transform 1 0 12444 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_346
timestamp 1581320205
transform 1 0 12036 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_347
timestamp 1581320205
transform 1 0 11424 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_348
timestamp 1581320205
transform 1 0 11016 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_349
timestamp 1581320205
transform 1 0 10608 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_350
timestamp 1581320205
transform 1 0 9996 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_351
timestamp 1581320205
transform 1 0 9588 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_352
timestamp 1581320205
transform 1 0 9384 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_353
timestamp 1581320205
transform 1 0 8976 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_354
timestamp 1581320205
transform 1 0 7548 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_355
timestamp 1581320205
transform 1 0 7140 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_356
timestamp 1581320205
transform 1 0 6936 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_357
timestamp 1581320205
transform 1 0 5916 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_358
timestamp 1581320205
transform 1 0 5712 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_359
timestamp 1581320205
transform 1 0 5508 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_360
timestamp 1581320205
transform 1 0 5100 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_361
timestamp 1581320205
transform 1 0 4896 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_362
timestamp 1581320205
transform 1 0 4692 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_363
timestamp 1581320205
transform 1 0 3672 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_364
timestamp 1581320205
transform 1 0 2448 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_365
timestamp 1581320205
transform 1 0 2040 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_366
timestamp 1581320205
transform 1 0 1632 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_367
timestamp 1581320205
transform 1 0 1020 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_368
timestamp 1581320205
transform 1 0 816 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_369
timestamp 1581320205
transform 1 0 408 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_370
timestamp 1581320205
transform 1 0 204 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_371
timestamp 1581320205
transform 1 0 0 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_372
timestamp 1581320205
transform 1 0 12852 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_373
timestamp 1581320205
transform 1 0 12648 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_374
timestamp 1581320205
transform 1 0 12240 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_375
timestamp 1581320205
transform 1 0 11832 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_376
timestamp 1581320205
transform 1 0 11628 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_377
timestamp 1581320205
transform 1 0 11220 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_378
timestamp 1581320205
transform 1 0 10608 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_379
timestamp 1581320205
transform 1 0 10200 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_380
timestamp 1581320205
transform 1 0 9996 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_381
timestamp 1581320205
transform 1 0 9792 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_382
timestamp 1581320205
transform 1 0 9180 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_383
timestamp 1581320205
transform 1 0 8976 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_384
timestamp 1581320205
transform 1 0 7548 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_385
timestamp 1581320205
transform 1 0 6936 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_386
timestamp 1581320205
transform 1 0 6732 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_387
timestamp 1581320205
transform 1 0 6120 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_388
timestamp 1581320205
transform 1 0 5508 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_389
timestamp 1581320205
transform 1 0 4692 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_390
timestamp 1581320205
transform 1 0 4284 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_391
timestamp 1581320205
transform 1 0 3876 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_392
timestamp 1581320205
transform 1 0 2856 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_393
timestamp 1581320205
transform 1 0 2652 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_394
timestamp 1581320205
transform 1 0 2448 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_395
timestamp 1581320205
transform 1 0 2244 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_396
timestamp 1581320205
transform 1 0 1836 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_397
timestamp 1581320205
transform 1 0 1632 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_398
timestamp 1581320205
transform 1 0 1428 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_399
timestamp 1581320205
transform 1 0 816 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_400
timestamp 1581320205
transform 1 0 408 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_401
timestamp 1581320205
transform 1 0 0 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_402
timestamp 1581320205
transform 1 0 12852 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_403
timestamp 1581320205
transform 1 0 12036 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_404
timestamp 1581320205
transform 1 0 11628 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_405
timestamp 1581320205
transform 1 0 11220 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_406
timestamp 1581320205
transform 1 0 11016 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_407
timestamp 1581320205
transform 1 0 10812 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_408
timestamp 1581320205
transform 1 0 9996 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_409
timestamp 1581320205
transform 1 0 9792 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_410
timestamp 1581320205
transform 1 0 9384 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_411
timestamp 1581320205
transform 1 0 8364 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_412
timestamp 1581320205
transform 1 0 7956 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_413
timestamp 1581320205
transform 1 0 7548 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_414
timestamp 1581320205
transform 1 0 7344 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_415
timestamp 1581320205
transform 1 0 6936 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_416
timestamp 1581320205
transform 1 0 6732 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_417
timestamp 1581320205
transform 1 0 5916 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_418
timestamp 1581320205
transform 1 0 5100 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_419
timestamp 1581320205
transform 1 0 4488 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_420
timestamp 1581320205
transform 1 0 4080 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_421
timestamp 1581320205
transform 1 0 3876 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_422
timestamp 1581320205
transform 1 0 3672 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_423
timestamp 1581320205
transform 1 0 3468 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_424
timestamp 1581320205
transform 1 0 3264 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_425
timestamp 1581320205
transform 1 0 3060 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_426
timestamp 1581320205
transform 1 0 2856 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_427
timestamp 1581320205
transform 1 0 2040 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_428
timestamp 1581320205
transform 1 0 816 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_429
timestamp 1581320205
transform 1 0 612 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_430
timestamp 1581320205
transform 1 0 408 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_431
timestamp 1581320205
transform 1 0 204 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_432
timestamp 1581320205
transform 1 0 0 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_433
timestamp 1581320205
transform 1 0 12852 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_434
timestamp 1581320205
transform 1 0 11832 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_435
timestamp 1581320205
transform 1 0 11424 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_436
timestamp 1581320205
transform 1 0 10812 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_437
timestamp 1581320205
transform 1 0 10608 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_438
timestamp 1581320205
transform 1 0 10404 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_439
timestamp 1581320205
transform 1 0 9996 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_440
timestamp 1581320205
transform 1 0 9588 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_441
timestamp 1581320205
transform 1 0 9384 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_442
timestamp 1581320205
transform 1 0 8772 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_443
timestamp 1581320205
transform 1 0 7752 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_444
timestamp 1581320205
transform 1 0 7140 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_445
timestamp 1581320205
transform 1 0 6936 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_446
timestamp 1581320205
transform 1 0 5916 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_447
timestamp 1581320205
transform 1 0 5712 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_448
timestamp 1581320205
transform 1 0 4488 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_449
timestamp 1581320205
transform 1 0 4284 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_450
timestamp 1581320205
transform 1 0 3876 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_451
timestamp 1581320205
transform 1 0 2652 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_452
timestamp 1581320205
transform 1 0 2040 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_453
timestamp 1581320205
transform 1 0 1836 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_454
timestamp 1581320205
transform 1 0 1428 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_455
timestamp 1581320205
transform 1 0 816 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_456
timestamp 1581320205
transform 1 0 408 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_457
timestamp 1581320205
transform 1 0 204 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_458
timestamp 1581320205
transform 1 0 0 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_459
timestamp 1581320205
transform 1 0 12852 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_460
timestamp 1581320205
transform 1 0 11832 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_461
timestamp 1581320205
transform 1 0 11424 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_462
timestamp 1581320205
transform 1 0 11220 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_463
timestamp 1581320205
transform 1 0 11016 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_464
timestamp 1581320205
transform 1 0 10812 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_465
timestamp 1581320205
transform 1 0 10608 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_466
timestamp 1581320205
transform 1 0 10200 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_467
timestamp 1581320205
transform 1 0 9996 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_468
timestamp 1581320205
transform 1 0 8976 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_469
timestamp 1581320205
transform 1 0 8772 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_470
timestamp 1581320205
transform 1 0 8160 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_471
timestamp 1581320205
transform 1 0 7956 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_472
timestamp 1581320205
transform 1 0 7752 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_473
timestamp 1581320205
transform 1 0 7548 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_474
timestamp 1581320205
transform 1 0 6732 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_475
timestamp 1581320205
transform 1 0 6324 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_476
timestamp 1581320205
transform 1 0 5712 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_477
timestamp 1581320205
transform 1 0 5508 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_478
timestamp 1581320205
transform 1 0 5304 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_479
timestamp 1581320205
transform 1 0 4692 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_480
timestamp 1581320205
transform 1 0 4284 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_481
timestamp 1581320205
transform 1 0 4080 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_482
timestamp 1581320205
transform 1 0 3672 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_483
timestamp 1581320205
transform 1 0 3264 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_484
timestamp 1581320205
transform 1 0 2652 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_485
timestamp 1581320205
transform 1 0 2448 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_486
timestamp 1581320205
transform 1 0 2244 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_487
timestamp 1581320205
transform 1 0 2040 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_488
timestamp 1581320205
transform 1 0 1632 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_489
timestamp 1581320205
transform 1 0 1428 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_490
timestamp 1581320205
transform 1 0 12852 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_491
timestamp 1581320205
transform 1 0 12648 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_492
timestamp 1581320205
transform 1 0 12240 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_493
timestamp 1581320205
transform 1 0 11832 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_494
timestamp 1581320205
transform 1 0 11424 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_495
timestamp 1581320205
transform 1 0 11220 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_496
timestamp 1581320205
transform 1 0 10608 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_497
timestamp 1581320205
transform 1 0 9384 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_498
timestamp 1581320205
transform 1 0 8772 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_499
timestamp 1581320205
transform 1 0 8568 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_500
timestamp 1581320205
transform 1 0 8364 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_501
timestamp 1581320205
transform 1 0 8160 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_502
timestamp 1581320205
transform 1 0 7752 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_503
timestamp 1581320205
transform 1 0 7548 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_504
timestamp 1581320205
transform 1 0 7140 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_505
timestamp 1581320205
transform 1 0 6936 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_506
timestamp 1581320205
transform 1 0 6732 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_507
timestamp 1581320205
transform 1 0 6528 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_508
timestamp 1581320205
transform 1 0 6324 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_509
timestamp 1581320205
transform 1 0 5916 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_510
timestamp 1581320205
transform 1 0 5712 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_511
timestamp 1581320205
transform 1 0 5508 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_512
timestamp 1581320205
transform 1 0 4284 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_513
timestamp 1581320205
transform 1 0 3876 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_514
timestamp 1581320205
transform 1 0 3672 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_515
timestamp 1581320205
transform 1 0 3468 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_516
timestamp 1581320205
transform 1 0 2448 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_517
timestamp 1581320205
transform 1 0 2244 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_518
timestamp 1581320205
transform 1 0 2040 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_519
timestamp 1581320205
transform 1 0 1632 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_520
timestamp 1581320205
transform 1 0 612 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_521
timestamp 1581320205
transform 1 0 12648 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_522
timestamp 1581320205
transform 1 0 12444 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_523
timestamp 1581320205
transform 1 0 12036 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_524
timestamp 1581320205
transform 1 0 11628 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_525
timestamp 1581320205
transform 1 0 11424 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_526
timestamp 1581320205
transform 1 0 10812 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_527
timestamp 1581320205
transform 1 0 10608 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_528
timestamp 1581320205
transform 1 0 10200 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_529
timestamp 1581320205
transform 1 0 9996 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_530
timestamp 1581320205
transform 1 0 9792 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_531
timestamp 1581320205
transform 1 0 8976 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_532
timestamp 1581320205
transform 1 0 8772 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_533
timestamp 1581320205
transform 1 0 8364 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_534
timestamp 1581320205
transform 1 0 8160 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_535
timestamp 1581320205
transform 1 0 7956 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_536
timestamp 1581320205
transform 1 0 7548 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_537
timestamp 1581320205
transform 1 0 7344 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_538
timestamp 1581320205
transform 1 0 6936 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_539
timestamp 1581320205
transform 1 0 6324 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_540
timestamp 1581320205
transform 1 0 5916 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_541
timestamp 1581320205
transform 1 0 5100 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_542
timestamp 1581320205
transform 1 0 4692 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_543
timestamp 1581320205
transform 1 0 4488 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_544
timestamp 1581320205
transform 1 0 4080 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_545
timestamp 1581320205
transform 1 0 3468 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_546
timestamp 1581320205
transform 1 0 3264 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_547
timestamp 1581320205
transform 1 0 612 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_548
timestamp 1581320205
transform 1 0 204 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_549
timestamp 1581320205
transform 1 0 12852 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_550
timestamp 1581320205
transform 1 0 12648 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_551
timestamp 1581320205
transform 1 0 12444 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_552
timestamp 1581320205
transform 1 0 12036 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_553
timestamp 1581320205
transform 1 0 11832 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_554
timestamp 1581320205
transform 1 0 11220 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_555
timestamp 1581320205
transform 1 0 10200 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_556
timestamp 1581320205
transform 1 0 9996 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_557
timestamp 1581320205
transform 1 0 9792 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_558
timestamp 1581320205
transform 1 0 9588 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_559
timestamp 1581320205
transform 1 0 8976 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_560
timestamp 1581320205
transform 1 0 8160 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_561
timestamp 1581320205
transform 1 0 7752 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_562
timestamp 1581320205
transform 1 0 7548 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_563
timestamp 1581320205
transform 1 0 6732 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_564
timestamp 1581320205
transform 1 0 5712 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_565
timestamp 1581320205
transform 1 0 5508 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_566
timestamp 1581320205
transform 1 0 4692 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_567
timestamp 1581320205
transform 1 0 4488 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_568
timestamp 1581320205
transform 1 0 4284 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_569
timestamp 1581320205
transform 1 0 3672 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_570
timestamp 1581320205
transform 1 0 3060 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_571
timestamp 1581320205
transform 1 0 2244 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_572
timestamp 1581320205
transform 1 0 2040 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_573
timestamp 1581320205
transform 1 0 1836 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_574
timestamp 1581320205
transform 1 0 204 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_575
timestamp 1581320205
transform 1 0 12852 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_576
timestamp 1581320205
transform 1 0 12648 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_577
timestamp 1581320205
transform 1 0 12444 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_578
timestamp 1581320205
transform 1 0 12240 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_579
timestamp 1581320205
transform 1 0 12036 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_580
timestamp 1581320205
transform 1 0 11832 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_581
timestamp 1581320205
transform 1 0 11220 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_582
timestamp 1581320205
transform 1 0 10812 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_583
timestamp 1581320205
transform 1 0 10404 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_584
timestamp 1581320205
transform 1 0 10200 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_585
timestamp 1581320205
transform 1 0 9792 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_586
timestamp 1581320205
transform 1 0 9588 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_587
timestamp 1581320205
transform 1 0 9180 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_588
timestamp 1581320205
transform 1 0 8976 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_589
timestamp 1581320205
transform 1 0 8160 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_590
timestamp 1581320205
transform 1 0 6936 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_591
timestamp 1581320205
transform 1 0 6120 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_592
timestamp 1581320205
transform 1 0 5712 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_593
timestamp 1581320205
transform 1 0 5508 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_594
timestamp 1581320205
transform 1 0 4284 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_595
timestamp 1581320205
transform 1 0 3876 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_596
timestamp 1581320205
transform 1 0 3468 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_597
timestamp 1581320205
transform 1 0 3060 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_598
timestamp 1581320205
transform 1 0 2448 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_599
timestamp 1581320205
transform 1 0 2244 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_600
timestamp 1581320205
transform 1 0 1836 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_601
timestamp 1581320205
transform 1 0 1632 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_602
timestamp 1581320205
transform 1 0 1224 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_603
timestamp 1581320205
transform 1 0 1020 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_604
timestamp 1581320205
transform 1 0 816 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_605
timestamp 1581320205
transform 1 0 612 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_606
timestamp 1581320205
transform 1 0 204 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_607
timestamp 1581320205
transform 1 0 0 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_608
timestamp 1581320205
transform 1 0 12852 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_609
timestamp 1581320205
transform 1 0 12648 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_610
timestamp 1581320205
transform 1 0 12444 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_611
timestamp 1581320205
transform 1 0 12240 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_612
timestamp 1581320205
transform 1 0 11832 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_613
timestamp 1581320205
transform 1 0 11628 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_614
timestamp 1581320205
transform 1 0 11220 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_615
timestamp 1581320205
transform 1 0 11016 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_616
timestamp 1581320205
transform 1 0 10608 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_617
timestamp 1581320205
transform 1 0 10200 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_618
timestamp 1581320205
transform 1 0 9996 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_619
timestamp 1581320205
transform 1 0 9588 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_620
timestamp 1581320205
transform 1 0 9384 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_621
timestamp 1581320205
transform 1 0 8976 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_622
timestamp 1581320205
transform 1 0 8568 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_623
timestamp 1581320205
transform 1 0 7752 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_624
timestamp 1581320205
transform 1 0 7548 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_625
timestamp 1581320205
transform 1 0 7344 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_626
timestamp 1581320205
transform 1 0 7140 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_627
timestamp 1581320205
transform 1 0 6120 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_628
timestamp 1581320205
transform 1 0 5916 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_629
timestamp 1581320205
transform 1 0 5712 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_630
timestamp 1581320205
transform 1 0 4896 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_631
timestamp 1581320205
transform 1 0 4488 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_632
timestamp 1581320205
transform 1 0 4080 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_633
timestamp 1581320205
transform 1 0 3672 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_634
timestamp 1581320205
transform 1 0 3264 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_635
timestamp 1581320205
transform 1 0 3060 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_636
timestamp 1581320205
transform 1 0 2856 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_637
timestamp 1581320205
transform 1 0 2652 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_638
timestamp 1581320205
transform 1 0 2244 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_639
timestamp 1581320205
transform 1 0 1428 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_640
timestamp 1581320205
transform 1 0 816 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_641
timestamp 1581320205
transform 1 0 612 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_642
timestamp 1581320205
transform 1 0 0 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_643
timestamp 1581320205
transform 1 0 12852 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_644
timestamp 1581320205
transform 1 0 12444 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_645
timestamp 1581320205
transform 1 0 11832 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_646
timestamp 1581320205
transform 1 0 11016 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_647
timestamp 1581320205
transform 1 0 10404 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_648
timestamp 1581320205
transform 1 0 9996 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_649
timestamp 1581320205
transform 1 0 9588 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_650
timestamp 1581320205
transform 1 0 9384 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_651
timestamp 1581320205
transform 1 0 8364 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_652
timestamp 1581320205
transform 1 0 7956 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_653
timestamp 1581320205
transform 1 0 7344 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_654
timestamp 1581320205
transform 1 0 6732 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_655
timestamp 1581320205
transform 1 0 6528 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_656
timestamp 1581320205
transform 1 0 5916 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_657
timestamp 1581320205
transform 1 0 5508 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_658
timestamp 1581320205
transform 1 0 5304 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_659
timestamp 1581320205
transform 1 0 5100 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_660
timestamp 1581320205
transform 1 0 4896 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_661
timestamp 1581320205
transform 1 0 4692 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_662
timestamp 1581320205
transform 1 0 4284 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_663
timestamp 1581320205
transform 1 0 4080 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_664
timestamp 1581320205
transform 1 0 3468 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_665
timestamp 1581320205
transform 1 0 3060 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_666
timestamp 1581320205
transform 1 0 2856 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_667
timestamp 1581320205
transform 1 0 2244 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_668
timestamp 1581320205
transform 1 0 2040 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_669
timestamp 1581320205
transform 1 0 1224 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_670
timestamp 1581320205
transform 1 0 816 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_671
timestamp 1581320205
transform 1 0 0 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_672
timestamp 1581320205
transform 1 0 12444 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_673
timestamp 1581320205
transform 1 0 11832 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_674
timestamp 1581320205
transform 1 0 11220 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_675
timestamp 1581320205
transform 1 0 10608 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_676
timestamp 1581320205
transform 1 0 8976 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_677
timestamp 1581320205
transform 1 0 8772 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_678
timestamp 1581320205
transform 1 0 8160 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_679
timestamp 1581320205
transform 1 0 7956 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_680
timestamp 1581320205
transform 1 0 7752 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_681
timestamp 1581320205
transform 1 0 7548 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_682
timestamp 1581320205
transform 1 0 7140 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_683
timestamp 1581320205
transform 1 0 6936 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_684
timestamp 1581320205
transform 1 0 6528 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_685
timestamp 1581320205
transform 1 0 6324 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_686
timestamp 1581320205
transform 1 0 5916 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_687
timestamp 1581320205
transform 1 0 5712 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_688
timestamp 1581320205
transform 1 0 5508 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_689
timestamp 1581320205
transform 1 0 5100 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_690
timestamp 1581320205
transform 1 0 4896 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_691
timestamp 1581320205
transform 1 0 4284 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_692
timestamp 1581320205
transform 1 0 4080 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_693
timestamp 1581320205
transform 1 0 3672 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_694
timestamp 1581320205
transform 1 0 3468 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_695
timestamp 1581320205
transform 1 0 3060 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_696
timestamp 1581320205
transform 1 0 2652 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_697
timestamp 1581320205
transform 1 0 2448 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_698
timestamp 1581320205
transform 1 0 2244 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_699
timestamp 1581320205
transform 1 0 1632 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_700
timestamp 1581320205
transform 1 0 1428 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_701
timestamp 1581320205
transform 1 0 1224 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_702
timestamp 1581320205
transform 1 0 1020 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_703
timestamp 1581320205
transform 1 0 612 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_704
timestamp 1581320205
transform 1 0 408 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_705
timestamp 1581320205
transform 1 0 204 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_706
timestamp 1581320205
transform 1 0 12036 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_707
timestamp 1581320205
transform 1 0 11628 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_708
timestamp 1581320205
transform 1 0 11424 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_709
timestamp 1581320205
transform 1 0 11220 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_710
timestamp 1581320205
transform 1 0 10608 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_711
timestamp 1581320205
transform 1 0 10404 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_712
timestamp 1581320205
transform 1 0 9384 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_713
timestamp 1581320205
transform 1 0 9180 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_714
timestamp 1581320205
transform 1 0 8772 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_715
timestamp 1581320205
transform 1 0 8568 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_716
timestamp 1581320205
transform 1 0 8160 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_717
timestamp 1581320205
transform 1 0 7956 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_718
timestamp 1581320205
transform 1 0 7344 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_719
timestamp 1581320205
transform 1 0 7140 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_720
timestamp 1581320205
transform 1 0 6936 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_721
timestamp 1581320205
transform 1 0 6732 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_722
timestamp 1581320205
transform 1 0 6528 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_723
timestamp 1581320205
transform 1 0 5916 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_724
timestamp 1581320205
transform 1 0 4692 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_725
timestamp 1581320205
transform 1 0 4284 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_726
timestamp 1581320205
transform 1 0 3876 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_727
timestamp 1581320205
transform 1 0 3672 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_728
timestamp 1581320205
transform 1 0 3468 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_729
timestamp 1581320205
transform 1 0 3264 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_730
timestamp 1581320205
transform 1 0 2652 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_731
timestamp 1581320205
transform 1 0 2448 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_732
timestamp 1581320205
transform 1 0 2244 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_733
timestamp 1581320205
transform 1 0 1836 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_734
timestamp 1581320205
transform 1 0 1428 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_735
timestamp 1581320205
transform 1 0 1224 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_736
timestamp 1581320205
transform 1 0 204 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_737
timestamp 1581320205
transform 1 0 12648 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_738
timestamp 1581320205
transform 1 0 11832 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_739
timestamp 1581320205
transform 1 0 11628 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_740
timestamp 1581320205
transform 1 0 11424 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_741
timestamp 1581320205
transform 1 0 10404 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_742
timestamp 1581320205
transform 1 0 9792 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_743
timestamp 1581320205
transform 1 0 9588 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_744
timestamp 1581320205
transform 1 0 9180 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_745
timestamp 1581320205
transform 1 0 8976 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_746
timestamp 1581320205
transform 1 0 8772 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_747
timestamp 1581320205
transform 1 0 8568 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_748
timestamp 1581320205
transform 1 0 8160 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_749
timestamp 1581320205
transform 1 0 7956 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_750
timestamp 1581320205
transform 1 0 7548 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_751
timestamp 1581320205
transform 1 0 6936 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_752
timestamp 1581320205
transform 1 0 6528 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_753
timestamp 1581320205
transform 1 0 5304 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_754
timestamp 1581320205
transform 1 0 4488 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_755
timestamp 1581320205
transform 1 0 4080 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_756
timestamp 1581320205
transform 1 0 3060 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_757
timestamp 1581320205
transform 1 0 2244 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_758
timestamp 1581320205
transform 1 0 1836 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_759
timestamp 1581320205
transform 1 0 1428 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_760
timestamp 1581320205
transform 1 0 1224 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_761
timestamp 1581320205
transform 1 0 612 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_762
timestamp 1581320205
transform 1 0 408 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_763
timestamp 1581320205
transform 1 0 204 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_764
timestamp 1581320205
transform 1 0 12648 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_765
timestamp 1581320205
transform 1 0 12240 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_766
timestamp 1581320205
transform 1 0 12036 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_767
timestamp 1581320205
transform 1 0 11832 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_768
timestamp 1581320205
transform 1 0 11628 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_769
timestamp 1581320205
transform 1 0 11220 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_770
timestamp 1581320205
transform 1 0 11016 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_771
timestamp 1581320205
transform 1 0 10812 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_772
timestamp 1581320205
transform 1 0 10608 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_773
timestamp 1581320205
transform 1 0 9996 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_774
timestamp 1581320205
transform 1 0 9588 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_775
timestamp 1581320205
transform 1 0 9384 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_776
timestamp 1581320205
transform 1 0 9180 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_777
timestamp 1581320205
transform 1 0 8976 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_778
timestamp 1581320205
transform 1 0 8160 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_779
timestamp 1581320205
transform 1 0 7548 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_780
timestamp 1581320205
transform 1 0 7344 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_781
timestamp 1581320205
transform 1 0 6936 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_782
timestamp 1581320205
transform 1 0 6732 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_783
timestamp 1581320205
transform 1 0 5916 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_784
timestamp 1581320205
transform 1 0 5100 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_785
timestamp 1581320205
transform 1 0 4284 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_786
timestamp 1581320205
transform 1 0 4080 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_787
timestamp 1581320205
transform 1 0 3672 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_788
timestamp 1581320205
transform 1 0 3264 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_789
timestamp 1581320205
transform 1 0 2856 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_790
timestamp 1581320205
transform 1 0 2448 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_791
timestamp 1581320205
transform 1 0 2244 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_792
timestamp 1581320205
transform 1 0 2040 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_793
timestamp 1581320205
transform 1 0 1632 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_794
timestamp 1581320205
transform 1 0 1428 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_795
timestamp 1581320205
transform 1 0 1020 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_796
timestamp 1581320205
transform 1 0 816 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_797
timestamp 1581320205
transform 1 0 612 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_798
timestamp 1581320205
transform 1 0 204 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_799
timestamp 1581320205
transform 1 0 0 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_800
timestamp 1581320205
transform 1 0 12648 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_801
timestamp 1581320205
transform 1 0 12444 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_802
timestamp 1581320205
transform 1 0 12240 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_803
timestamp 1581320205
transform 1 0 12036 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_804
timestamp 1581320205
transform 1 0 11424 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_805
timestamp 1581320205
transform 1 0 10812 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_806
timestamp 1581320205
transform 1 0 10404 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_807
timestamp 1581320205
transform 1 0 10200 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_808
timestamp 1581320205
transform 1 0 9792 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_809
timestamp 1581320205
transform 1 0 9588 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_810
timestamp 1581320205
transform 1 0 8772 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_811
timestamp 1581320205
transform 1 0 8568 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_812
timestamp 1581320205
transform 1 0 8364 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_813
timestamp 1581320205
transform 1 0 7548 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_814
timestamp 1581320205
transform 1 0 6732 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_815
timestamp 1581320205
transform 1 0 6528 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_816
timestamp 1581320205
transform 1 0 6324 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_817
timestamp 1581320205
transform 1 0 6120 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_818
timestamp 1581320205
transform 1 0 5916 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_819
timestamp 1581320205
transform 1 0 5100 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_820
timestamp 1581320205
transform 1 0 4896 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_821
timestamp 1581320205
transform 1 0 4692 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_822
timestamp 1581320205
transform 1 0 4488 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_823
timestamp 1581320205
transform 1 0 3876 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_824
timestamp 1581320205
transform 1 0 3060 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_825
timestamp 1581320205
transform 1 0 2856 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_826
timestamp 1581320205
transform 1 0 2448 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_827
timestamp 1581320205
transform 1 0 1836 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_828
timestamp 1581320205
transform 1 0 1224 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_829
timestamp 1581320205
transform 1 0 1020 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_830
timestamp 1581320205
transform 1 0 816 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_831
timestamp 1581320205
transform 1 0 612 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_832
timestamp 1581320205
transform 1 0 204 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_833
timestamp 1581320205
transform 1 0 0 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_834
timestamp 1581320205
transform 1 0 12648 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_835
timestamp 1581320205
transform 1 0 11832 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_836
timestamp 1581320205
transform 1 0 11220 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_837
timestamp 1581320205
transform 1 0 10812 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_838
timestamp 1581320205
transform 1 0 9996 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_839
timestamp 1581320205
transform 1 0 9792 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_840
timestamp 1581320205
transform 1 0 9588 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_841
timestamp 1581320205
transform 1 0 9180 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_842
timestamp 1581320205
transform 1 0 8772 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_843
timestamp 1581320205
transform 1 0 8568 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_844
timestamp 1581320205
transform 1 0 8364 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_845
timestamp 1581320205
transform 1 0 7956 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_846
timestamp 1581320205
transform 1 0 7548 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_847
timestamp 1581320205
transform 1 0 6936 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_848
timestamp 1581320205
transform 1 0 6732 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_849
timestamp 1581320205
transform 1 0 6324 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_850
timestamp 1581320205
transform 1 0 6120 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_851
timestamp 1581320205
transform 1 0 5916 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_852
timestamp 1581320205
transform 1 0 5508 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_853
timestamp 1581320205
transform 1 0 5304 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_854
timestamp 1581320205
transform 1 0 5100 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_855
timestamp 1581320205
transform 1 0 4896 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_856
timestamp 1581320205
transform 1 0 4692 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_857
timestamp 1581320205
transform 1 0 4488 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_858
timestamp 1581320205
transform 1 0 3876 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_859
timestamp 1581320205
transform 1 0 3468 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_860
timestamp 1581320205
transform 1 0 3264 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_861
timestamp 1581320205
transform 1 0 3060 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_862
timestamp 1581320205
transform 1 0 2652 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_863
timestamp 1581320205
transform 1 0 2244 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_864
timestamp 1581320205
transform 1 0 2040 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_865
timestamp 1581320205
transform 1 0 1632 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_866
timestamp 1581320205
transform 1 0 1428 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_867
timestamp 1581320205
transform 1 0 1224 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_868
timestamp 1581320205
transform 1 0 1020 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_869
timestamp 1581320205
transform 1 0 816 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_870
timestamp 1581320205
transform 1 0 204 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_871
timestamp 1581320205
transform 1 0 12852 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_872
timestamp 1581320205
transform 1 0 12648 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_873
timestamp 1581320205
transform 1 0 12240 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_874
timestamp 1581320205
transform 1 0 11832 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_875
timestamp 1581320205
transform 1 0 11628 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_876
timestamp 1581320205
transform 1 0 11220 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_877
timestamp 1581320205
transform 1 0 10404 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_878
timestamp 1581320205
transform 1 0 9384 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_879
timestamp 1581320205
transform 1 0 9180 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_880
timestamp 1581320205
transform 1 0 8976 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_881
timestamp 1581320205
transform 1 0 8772 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_882
timestamp 1581320205
transform 1 0 8568 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_883
timestamp 1581320205
transform 1 0 8160 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_884
timestamp 1581320205
transform 1 0 7752 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_885
timestamp 1581320205
transform 1 0 7548 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_886
timestamp 1581320205
transform 1 0 7140 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_887
timestamp 1581320205
transform 1 0 6120 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_888
timestamp 1581320205
transform 1 0 5712 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_889
timestamp 1581320205
transform 1 0 5508 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_890
timestamp 1581320205
transform 1 0 5100 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_891
timestamp 1581320205
transform 1 0 4488 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_892
timestamp 1581320205
transform 1 0 3876 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_893
timestamp 1581320205
transform 1 0 3468 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_894
timestamp 1581320205
transform 1 0 3264 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_895
timestamp 1581320205
transform 1 0 3060 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_896
timestamp 1581320205
transform 1 0 2856 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_897
timestamp 1581320205
transform 1 0 2448 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_898
timestamp 1581320205
transform 1 0 1428 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_899
timestamp 1581320205
transform 1 0 612 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_900
timestamp 1581320205
transform 1 0 408 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_901
timestamp 1581320205
transform 1 0 12852 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_902
timestamp 1581320205
transform 1 0 12648 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_903
timestamp 1581320205
transform 1 0 12444 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_904
timestamp 1581320205
transform 1 0 11628 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_905
timestamp 1581320205
transform 1 0 11016 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_906
timestamp 1581320205
transform 1 0 10812 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_907
timestamp 1581320205
transform 1 0 10608 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_908
timestamp 1581320205
transform 1 0 10200 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_909
timestamp 1581320205
transform 1 0 9996 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_910
timestamp 1581320205
transform 1 0 8364 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_911
timestamp 1581320205
transform 1 0 7752 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_912
timestamp 1581320205
transform 1 0 7140 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_913
timestamp 1581320205
transform 1 0 6936 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_914
timestamp 1581320205
transform 1 0 6528 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_915
timestamp 1581320205
transform 1 0 6120 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_916
timestamp 1581320205
transform 1 0 5712 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_917
timestamp 1581320205
transform 1 0 5508 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_918
timestamp 1581320205
transform 1 0 4896 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_919
timestamp 1581320205
transform 1 0 3672 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_920
timestamp 1581320205
transform 1 0 2856 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_921
timestamp 1581320205
transform 1 0 1632 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_922
timestamp 1581320205
transform 1 0 1020 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_923
timestamp 1581320205
transform 1 0 612 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_924
timestamp 1581320205
transform 1 0 408 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_925
timestamp 1581320205
transform 1 0 0 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_926
timestamp 1581320205
transform 1 0 12852 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_927
timestamp 1581320205
transform 1 0 12240 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_928
timestamp 1581320205
transform 1 0 11628 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_929
timestamp 1581320205
transform 1 0 11016 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_930
timestamp 1581320205
transform 1 0 10608 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_931
timestamp 1581320205
transform 1 0 10200 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_932
timestamp 1581320205
transform 1 0 9996 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_933
timestamp 1581320205
transform 1 0 9792 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_934
timestamp 1581320205
transform 1 0 9588 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_935
timestamp 1581320205
transform 1 0 9384 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_936
timestamp 1581320205
transform 1 0 9180 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_937
timestamp 1581320205
transform 1 0 8772 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_938
timestamp 1581320205
transform 1 0 8364 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_939
timestamp 1581320205
transform 1 0 7752 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_940
timestamp 1581320205
transform 1 0 7548 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_941
timestamp 1581320205
transform 1 0 7344 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_942
timestamp 1581320205
transform 1 0 6732 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_943
timestamp 1581320205
transform 1 0 6324 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_944
timestamp 1581320205
transform 1 0 6120 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_945
timestamp 1581320205
transform 1 0 5916 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_946
timestamp 1581320205
transform 1 0 5100 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_947
timestamp 1581320205
transform 1 0 4896 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_948
timestamp 1581320205
transform 1 0 4080 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_949
timestamp 1581320205
transform 1 0 3876 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_950
timestamp 1581320205
transform 1 0 3468 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_951
timestamp 1581320205
transform 1 0 3060 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_952
timestamp 1581320205
transform 1 0 2856 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_953
timestamp 1581320205
transform 1 0 1428 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_954
timestamp 1581320205
transform 1 0 816 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_955
timestamp 1581320205
transform 1 0 612 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_956
timestamp 1581320205
transform 1 0 408 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_957
timestamp 1581320205
transform 1 0 0 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_958
timestamp 1581320205
transform 1 0 12852 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_959
timestamp 1581320205
transform 1 0 12648 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_960
timestamp 1581320205
transform 1 0 12444 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_961
timestamp 1581320205
transform 1 0 12240 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_962
timestamp 1581320205
transform 1 0 12036 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_963
timestamp 1581320205
transform 1 0 11424 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_964
timestamp 1581320205
transform 1 0 10404 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_965
timestamp 1581320205
transform 1 0 10200 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_966
timestamp 1581320205
transform 1 0 9996 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_967
timestamp 1581320205
transform 1 0 8364 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_968
timestamp 1581320205
transform 1 0 7344 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_969
timestamp 1581320205
transform 1 0 7140 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_970
timestamp 1581320205
transform 1 0 6528 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_971
timestamp 1581320205
transform 1 0 6324 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_972
timestamp 1581320205
transform 1 0 6120 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_973
timestamp 1581320205
transform 1 0 5916 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_974
timestamp 1581320205
transform 1 0 5712 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_975
timestamp 1581320205
transform 1 0 5508 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_976
timestamp 1581320205
transform 1 0 5100 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_977
timestamp 1581320205
transform 1 0 4896 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_978
timestamp 1581320205
transform 1 0 4692 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_979
timestamp 1581320205
transform 1 0 4284 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_980
timestamp 1581320205
transform 1 0 3264 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_981
timestamp 1581320205
transform 1 0 3060 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_982
timestamp 1581320205
transform 1 0 2652 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_983
timestamp 1581320205
transform 1 0 2448 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_984
timestamp 1581320205
transform 1 0 2244 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_985
timestamp 1581320205
transform 1 0 2040 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_986
timestamp 1581320205
transform 1 0 1836 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_987
timestamp 1581320205
transform 1 0 1428 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_988
timestamp 1581320205
transform 1 0 1020 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_989
timestamp 1581320205
transform 1 0 408 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_990
timestamp 1581320205
transform 1 0 12852 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_991
timestamp 1581320205
transform 1 0 12648 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_992
timestamp 1581320205
transform 1 0 12444 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_993
timestamp 1581320205
transform 1 0 12240 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_994
timestamp 1581320205
transform 1 0 12036 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_995
timestamp 1581320205
transform 1 0 11832 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_996
timestamp 1581320205
transform 1 0 11424 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_997
timestamp 1581320205
transform 1 0 11016 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_998
timestamp 1581320205
transform 1 0 10404 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_999
timestamp 1581320205
transform 1 0 10200 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1000
timestamp 1581320205
transform 1 0 9588 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1001
timestamp 1581320205
transform 1 0 9180 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1002
timestamp 1581320205
transform 1 0 8772 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1003
timestamp 1581320205
transform 1 0 8160 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1004
timestamp 1581320205
transform 1 0 7752 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1005
timestamp 1581320205
transform 1 0 7344 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1006
timestamp 1581320205
transform 1 0 7140 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1007
timestamp 1581320205
transform 1 0 6936 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1008
timestamp 1581320205
transform 1 0 6120 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1009
timestamp 1581320205
transform 1 0 5916 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1010
timestamp 1581320205
transform 1 0 5304 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1011
timestamp 1581320205
transform 1 0 4896 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1012
timestamp 1581320205
transform 1 0 4692 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1013
timestamp 1581320205
transform 1 0 4284 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1014
timestamp 1581320205
transform 1 0 4080 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1015
timestamp 1581320205
transform 1 0 3672 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1016
timestamp 1581320205
transform 1 0 3264 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1017
timestamp 1581320205
transform 1 0 2856 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1018
timestamp 1581320205
transform 1 0 2448 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1019
timestamp 1581320205
transform 1 0 2244 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1020
timestamp 1581320205
transform 1 0 2040 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1021
timestamp 1581320205
transform 1 0 1836 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1022
timestamp 1581320205
transform 1 0 1428 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1023
timestamp 1581320205
transform 1 0 1224 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1024
timestamp 1581320205
transform 1 0 1020 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1025
timestamp 1581320205
transform 1 0 816 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1026
timestamp 1581320205
transform 1 0 612 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1027
timestamp 1581320205
transform 1 0 408 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1028
timestamp 1581320205
transform 1 0 204 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1029
timestamp 1581320205
transform 1 0 0 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1030
timestamp 1581320205
transform 1 0 12852 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1031
timestamp 1581320205
transform 1 0 12444 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1032
timestamp 1581320205
transform 1 0 12240 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1033
timestamp 1581320205
transform 1 0 11832 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1034
timestamp 1581320205
transform 1 0 10812 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1035
timestamp 1581320205
transform 1 0 10200 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1036
timestamp 1581320205
transform 1 0 9996 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1037
timestamp 1581320205
transform 1 0 9792 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1038
timestamp 1581320205
transform 1 0 9384 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1039
timestamp 1581320205
transform 1 0 9180 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1040
timestamp 1581320205
transform 1 0 8568 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1041
timestamp 1581320205
transform 1 0 7140 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1042
timestamp 1581320205
transform 1 0 6936 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1043
timestamp 1581320205
transform 1 0 6732 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1044
timestamp 1581320205
transform 1 0 6324 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1045
timestamp 1581320205
transform 1 0 5916 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1046
timestamp 1581320205
transform 1 0 5712 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1047
timestamp 1581320205
transform 1 0 5508 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1048
timestamp 1581320205
transform 1 0 4284 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1049
timestamp 1581320205
transform 1 0 4080 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1050
timestamp 1581320205
transform 1 0 3672 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1051
timestamp 1581320205
transform 1 0 2856 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1052
timestamp 1581320205
transform 1 0 2448 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1053
timestamp 1581320205
transform 1 0 1632 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1054
timestamp 1581320205
transform 1 0 1428 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1055
timestamp 1581320205
transform 1 0 612 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1056
timestamp 1581320205
transform 1 0 204 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_0
timestamp 1581320205
transform 1 0 12852 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1
timestamp 1581320205
transform 1 0 12648 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_2
timestamp 1581320205
transform 1 0 12240 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_3
timestamp 1581320205
transform 1 0 11424 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_4
timestamp 1581320205
transform 1 0 11016 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_5
timestamp 1581320205
transform 1 0 10812 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_6
timestamp 1581320205
transform 1 0 9996 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_7
timestamp 1581320205
transform 1 0 9588 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_8
timestamp 1581320205
transform 1 0 9384 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_9
timestamp 1581320205
transform 1 0 9180 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_10
timestamp 1581320205
transform 1 0 8568 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_11
timestamp 1581320205
transform 1 0 8364 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_12
timestamp 1581320205
transform 1 0 7956 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_13
timestamp 1581320205
transform 1 0 7548 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_14
timestamp 1581320205
transform 1 0 7344 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_15
timestamp 1581320205
transform 1 0 7140 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_16
timestamp 1581320205
transform 1 0 6936 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_17
timestamp 1581320205
transform 1 0 5712 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_18
timestamp 1581320205
transform 1 0 5304 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_19
timestamp 1581320205
transform 1 0 4080 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_20
timestamp 1581320205
transform 1 0 2040 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_21
timestamp 1581320205
transform 1 0 1632 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_22
timestamp 1581320205
transform 1 0 1224 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_23
timestamp 1581320205
transform 1 0 1020 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_24
timestamp 1581320205
transform 1 0 12648 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_25
timestamp 1581320205
transform 1 0 12444 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_26
timestamp 1581320205
transform 1 0 12240 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_27
timestamp 1581320205
transform 1 0 12036 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_28
timestamp 1581320205
transform 1 0 11628 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_29
timestamp 1581320205
transform 1 0 11424 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_30
timestamp 1581320205
transform 1 0 11016 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_31
timestamp 1581320205
transform 1 0 10812 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_32
timestamp 1581320205
transform 1 0 10608 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_33
timestamp 1581320205
transform 1 0 9792 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_34
timestamp 1581320205
transform 1 0 9588 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_35
timestamp 1581320205
transform 1 0 9180 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_36
timestamp 1581320205
transform 1 0 8772 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_37
timestamp 1581320205
transform 1 0 8160 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_38
timestamp 1581320205
transform 1 0 7548 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_39
timestamp 1581320205
transform 1 0 7344 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_40
timestamp 1581320205
transform 1 0 6528 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_41
timestamp 1581320205
transform 1 0 6324 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_42
timestamp 1581320205
transform 1 0 6120 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_43
timestamp 1581320205
transform 1 0 5712 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_44
timestamp 1581320205
transform 1 0 4284 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_45
timestamp 1581320205
transform 1 0 3264 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_46
timestamp 1581320205
transform 1 0 2448 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_47
timestamp 1581320205
transform 1 0 1836 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_48
timestamp 1581320205
transform 1 0 1632 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_49
timestamp 1581320205
transform 1 0 1224 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_50
timestamp 1581320205
transform 1 0 1020 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_51
timestamp 1581320205
transform 1 0 12852 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_52
timestamp 1581320205
transform 1 0 12648 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_53
timestamp 1581320205
transform 1 0 12240 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_54
timestamp 1581320205
transform 1 0 12036 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_55
timestamp 1581320205
transform 1 0 11832 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_56
timestamp 1581320205
transform 1 0 11628 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_57
timestamp 1581320205
transform 1 0 11424 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_58
timestamp 1581320205
transform 1 0 11220 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_59
timestamp 1581320205
transform 1 0 10608 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_60
timestamp 1581320205
transform 1 0 10404 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_61
timestamp 1581320205
transform 1 0 10200 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_62
timestamp 1581320205
transform 1 0 9996 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_63
timestamp 1581320205
transform 1 0 9792 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_64
timestamp 1581320205
transform 1 0 9588 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_65
timestamp 1581320205
transform 1 0 9384 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_66
timestamp 1581320205
transform 1 0 8568 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_67
timestamp 1581320205
transform 1 0 8364 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_68
timestamp 1581320205
transform 1 0 7752 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_69
timestamp 1581320205
transform 1 0 7548 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_70
timestamp 1581320205
transform 1 0 7140 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_71
timestamp 1581320205
transform 1 0 6528 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_72
timestamp 1581320205
transform 1 0 6324 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_73
timestamp 1581320205
transform 1 0 6120 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_74
timestamp 1581320205
transform 1 0 5916 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_75
timestamp 1581320205
transform 1 0 5712 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_76
timestamp 1581320205
transform 1 0 5100 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_77
timestamp 1581320205
transform 1 0 4896 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_78
timestamp 1581320205
transform 1 0 4692 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_79
timestamp 1581320205
transform 1 0 4488 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_80
timestamp 1581320205
transform 1 0 4284 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_81
timestamp 1581320205
transform 1 0 4080 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_82
timestamp 1581320205
transform 1 0 3876 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_83
timestamp 1581320205
transform 1 0 3468 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_84
timestamp 1581320205
transform 1 0 3264 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_85
timestamp 1581320205
transform 1 0 3060 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_86
timestamp 1581320205
transform 1 0 2856 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_87
timestamp 1581320205
transform 1 0 2448 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_88
timestamp 1581320205
transform 1 0 2244 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_89
timestamp 1581320205
transform 1 0 1632 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_90
timestamp 1581320205
transform 1 0 1428 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_91
timestamp 1581320205
transform 1 0 1224 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_92
timestamp 1581320205
transform 1 0 612 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_93
timestamp 1581320205
transform 1 0 408 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_94
timestamp 1581320205
transform 1 0 12240 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_95
timestamp 1581320205
transform 1 0 12036 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_96
timestamp 1581320205
transform 1 0 11832 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_97
timestamp 1581320205
transform 1 0 11424 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_98
timestamp 1581320205
transform 1 0 10812 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_99
timestamp 1581320205
transform 1 0 10608 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_100
timestamp 1581320205
transform 1 0 9792 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_101
timestamp 1581320205
transform 1 0 9384 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_102
timestamp 1581320205
transform 1 0 8976 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_103
timestamp 1581320205
transform 1 0 8568 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_104
timestamp 1581320205
transform 1 0 7752 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_105
timestamp 1581320205
transform 1 0 7548 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_106
timestamp 1581320205
transform 1 0 6936 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_107
timestamp 1581320205
transform 1 0 6528 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_108
timestamp 1581320205
transform 1 0 6324 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_109
timestamp 1581320205
transform 1 0 6120 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_110
timestamp 1581320205
transform 1 0 5916 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_111
timestamp 1581320205
transform 1 0 5508 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_112
timestamp 1581320205
transform 1 0 5304 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_113
timestamp 1581320205
transform 1 0 5100 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_114
timestamp 1581320205
transform 1 0 3672 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_115
timestamp 1581320205
transform 1 0 3468 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_116
timestamp 1581320205
transform 1 0 2652 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_117
timestamp 1581320205
transform 1 0 2040 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_118
timestamp 1581320205
transform 1 0 1836 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_119
timestamp 1581320205
transform 1 0 1428 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_120
timestamp 1581320205
transform 1 0 1224 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_121
timestamp 1581320205
transform 1 0 816 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_122
timestamp 1581320205
transform 1 0 0 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_123
timestamp 1581320205
transform 1 0 12444 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_124
timestamp 1581320205
transform 1 0 12240 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_125
timestamp 1581320205
transform 1 0 11832 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_126
timestamp 1581320205
transform 1 0 11628 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_127
timestamp 1581320205
transform 1 0 10608 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_128
timestamp 1581320205
transform 1 0 9996 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_129
timestamp 1581320205
transform 1 0 9588 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_130
timestamp 1581320205
transform 1 0 8976 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_131
timestamp 1581320205
transform 1 0 8568 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_132
timestamp 1581320205
transform 1 0 8160 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_133
timestamp 1581320205
transform 1 0 7956 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_134
timestamp 1581320205
transform 1 0 6120 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_135
timestamp 1581320205
transform 1 0 5916 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_136
timestamp 1581320205
transform 1 0 5712 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_137
timestamp 1581320205
transform 1 0 5508 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_138
timestamp 1581320205
transform 1 0 5304 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_139
timestamp 1581320205
transform 1 0 3876 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_140
timestamp 1581320205
transform 1 0 3672 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_141
timestamp 1581320205
transform 1 0 3468 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_142
timestamp 1581320205
transform 1 0 3264 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_143
timestamp 1581320205
transform 1 0 2652 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_144
timestamp 1581320205
transform 1 0 1836 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_145
timestamp 1581320205
transform 1 0 1224 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_146
timestamp 1581320205
transform 1 0 1020 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_147
timestamp 1581320205
transform 1 0 816 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_148
timestamp 1581320205
transform 1 0 612 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_149
timestamp 1581320205
transform 1 0 0 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_150
timestamp 1581320205
transform 1 0 12852 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_151
timestamp 1581320205
transform 1 0 12648 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_152
timestamp 1581320205
transform 1 0 12444 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_153
timestamp 1581320205
transform 1 0 12240 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_154
timestamp 1581320205
transform 1 0 11832 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_155
timestamp 1581320205
transform 1 0 11628 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_156
timestamp 1581320205
transform 1 0 10812 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_157
timestamp 1581320205
transform 1 0 10200 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_158
timestamp 1581320205
transform 1 0 9996 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_159
timestamp 1581320205
transform 1 0 9792 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_160
timestamp 1581320205
transform 1 0 9588 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_161
timestamp 1581320205
transform 1 0 9384 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_162
timestamp 1581320205
transform 1 0 9180 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_163
timestamp 1581320205
transform 1 0 8772 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_164
timestamp 1581320205
transform 1 0 8160 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_165
timestamp 1581320205
transform 1 0 7140 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_166
timestamp 1581320205
transform 1 0 6324 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_167
timestamp 1581320205
transform 1 0 6120 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_168
timestamp 1581320205
transform 1 0 5712 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_169
timestamp 1581320205
transform 1 0 5304 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_170
timestamp 1581320205
transform 1 0 4692 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_171
timestamp 1581320205
transform 1 0 4284 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_172
timestamp 1581320205
transform 1 0 4080 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_173
timestamp 1581320205
transform 1 0 3672 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_174
timestamp 1581320205
transform 1 0 3468 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_175
timestamp 1581320205
transform 1 0 2856 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_176
timestamp 1581320205
transform 1 0 2244 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_177
timestamp 1581320205
transform 1 0 2040 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_178
timestamp 1581320205
transform 1 0 1836 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_179
timestamp 1581320205
transform 1 0 1632 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_180
timestamp 1581320205
transform 1 0 1428 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_181
timestamp 1581320205
transform 1 0 816 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_182
timestamp 1581320205
transform 1 0 408 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_183
timestamp 1581320205
transform 1 0 204 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_184
timestamp 1581320205
transform 1 0 0 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_185
timestamp 1581320205
transform 1 0 12648 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_186
timestamp 1581320205
transform 1 0 12444 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_187
timestamp 1581320205
transform 1 0 12240 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_188
timestamp 1581320205
transform 1 0 12036 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_189
timestamp 1581320205
transform 1 0 11628 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_190
timestamp 1581320205
transform 1 0 11220 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_191
timestamp 1581320205
transform 1 0 11016 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_192
timestamp 1581320205
transform 1 0 10812 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_193
timestamp 1581320205
transform 1 0 10608 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_194
timestamp 1581320205
transform 1 0 10404 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_195
timestamp 1581320205
transform 1 0 9996 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_196
timestamp 1581320205
transform 1 0 9180 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_197
timestamp 1581320205
transform 1 0 8364 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_198
timestamp 1581320205
transform 1 0 7956 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_199
timestamp 1581320205
transform 1 0 7548 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_200
timestamp 1581320205
transform 1 0 7344 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_201
timestamp 1581320205
transform 1 0 6936 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_202
timestamp 1581320205
transform 1 0 6528 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_203
timestamp 1581320205
transform 1 0 5508 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_204
timestamp 1581320205
transform 1 0 5100 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_205
timestamp 1581320205
transform 1 0 4896 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_206
timestamp 1581320205
transform 1 0 3876 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_207
timestamp 1581320205
transform 1 0 3468 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_208
timestamp 1581320205
transform 1 0 3060 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_209
timestamp 1581320205
transform 1 0 2856 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_210
timestamp 1581320205
transform 1 0 2652 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_211
timestamp 1581320205
transform 1 0 2448 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_212
timestamp 1581320205
transform 1 0 1632 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_213
timestamp 1581320205
transform 1 0 816 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_214
timestamp 1581320205
transform 1 0 612 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_215
timestamp 1581320205
transform 1 0 408 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_216
timestamp 1581320205
transform 1 0 204 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_217
timestamp 1581320205
transform 1 0 0 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_218
timestamp 1581320205
transform 1 0 12852 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_219
timestamp 1581320205
transform 1 0 12648 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_220
timestamp 1581320205
transform 1 0 12240 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_221
timestamp 1581320205
transform 1 0 12036 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_222
timestamp 1581320205
transform 1 0 11628 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_223
timestamp 1581320205
transform 1 0 11220 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_224
timestamp 1581320205
transform 1 0 11016 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_225
timestamp 1581320205
transform 1 0 10200 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_226
timestamp 1581320205
transform 1 0 9996 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_227
timestamp 1581320205
transform 1 0 9792 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_228
timestamp 1581320205
transform 1 0 9588 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_229
timestamp 1581320205
transform 1 0 8568 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_230
timestamp 1581320205
transform 1 0 8160 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_231
timestamp 1581320205
transform 1 0 7548 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_232
timestamp 1581320205
transform 1 0 7140 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_233
timestamp 1581320205
transform 1 0 6936 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_234
timestamp 1581320205
transform 1 0 6732 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_235
timestamp 1581320205
transform 1 0 6324 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_236
timestamp 1581320205
transform 1 0 6120 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_237
timestamp 1581320205
transform 1 0 5304 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_238
timestamp 1581320205
transform 1 0 5100 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_239
timestamp 1581320205
transform 1 0 4692 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_240
timestamp 1581320205
transform 1 0 4080 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_241
timestamp 1581320205
transform 1 0 3876 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_242
timestamp 1581320205
transform 1 0 3672 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_243
timestamp 1581320205
transform 1 0 3264 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_244
timestamp 1581320205
transform 1 0 3060 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_245
timestamp 1581320205
transform 1 0 2652 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_246
timestamp 1581320205
transform 1 0 2448 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_247
timestamp 1581320205
transform 1 0 2244 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_248
timestamp 1581320205
transform 1 0 1836 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_249
timestamp 1581320205
transform 1 0 1632 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_250
timestamp 1581320205
transform 1 0 1428 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_251
timestamp 1581320205
transform 1 0 1224 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_252
timestamp 1581320205
transform 1 0 1020 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_253
timestamp 1581320205
transform 1 0 816 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_254
timestamp 1581320205
transform 1 0 612 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_255
timestamp 1581320205
transform 1 0 0 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_256
timestamp 1581320205
transform 1 0 12852 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_257
timestamp 1581320205
transform 1 0 12648 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_258
timestamp 1581320205
transform 1 0 12444 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_259
timestamp 1581320205
transform 1 0 12240 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_260
timestamp 1581320205
transform 1 0 11628 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_261
timestamp 1581320205
transform 1 0 11424 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_262
timestamp 1581320205
transform 1 0 11220 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_263
timestamp 1581320205
transform 1 0 11016 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_264
timestamp 1581320205
transform 1 0 10608 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_265
timestamp 1581320205
transform 1 0 10404 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_266
timestamp 1581320205
transform 1 0 10200 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_267
timestamp 1581320205
transform 1 0 9792 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_268
timestamp 1581320205
transform 1 0 9588 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_269
timestamp 1581320205
transform 1 0 9384 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_270
timestamp 1581320205
transform 1 0 9180 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_271
timestamp 1581320205
transform 1 0 8976 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_272
timestamp 1581320205
transform 1 0 7956 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_273
timestamp 1581320205
transform 1 0 7752 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_274
timestamp 1581320205
transform 1 0 7344 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_275
timestamp 1581320205
transform 1 0 7140 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_276
timestamp 1581320205
transform 1 0 6936 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_277
timestamp 1581320205
transform 1 0 6528 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_278
timestamp 1581320205
transform 1 0 6120 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_279
timestamp 1581320205
transform 1 0 5916 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_280
timestamp 1581320205
transform 1 0 5508 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_281
timestamp 1581320205
transform 1 0 5100 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_282
timestamp 1581320205
transform 1 0 4080 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_283
timestamp 1581320205
transform 1 0 3876 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_284
timestamp 1581320205
transform 1 0 3468 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_285
timestamp 1581320205
transform 1 0 2856 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_286
timestamp 1581320205
transform 1 0 2448 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_287
timestamp 1581320205
transform 1 0 2244 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_288
timestamp 1581320205
transform 1 0 2040 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_289
timestamp 1581320205
transform 1 0 1836 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_290
timestamp 1581320205
transform 1 0 1428 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_291
timestamp 1581320205
transform 1 0 1020 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_292
timestamp 1581320205
transform 1 0 816 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_293
timestamp 1581320205
transform 1 0 408 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_294
timestamp 1581320205
transform 1 0 204 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_295
timestamp 1581320205
transform 1 0 12852 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_296
timestamp 1581320205
transform 1 0 12648 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_297
timestamp 1581320205
transform 1 0 12240 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_298
timestamp 1581320205
transform 1 0 11832 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_299
timestamp 1581320205
transform 1 0 11628 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_300
timestamp 1581320205
transform 1 0 11220 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_301
timestamp 1581320205
transform 1 0 10812 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_302
timestamp 1581320205
transform 1 0 10404 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_303
timestamp 1581320205
transform 1 0 10200 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_304
timestamp 1581320205
transform 1 0 9792 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_305
timestamp 1581320205
transform 1 0 9180 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_306
timestamp 1581320205
transform 1 0 8772 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_307
timestamp 1581320205
transform 1 0 8568 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_308
timestamp 1581320205
transform 1 0 8364 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_309
timestamp 1581320205
transform 1 0 8160 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_310
timestamp 1581320205
transform 1 0 7956 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_311
timestamp 1581320205
transform 1 0 7752 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_312
timestamp 1581320205
transform 1 0 7344 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_313
timestamp 1581320205
transform 1 0 6732 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_314
timestamp 1581320205
transform 1 0 6528 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_315
timestamp 1581320205
transform 1 0 6324 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_316
timestamp 1581320205
transform 1 0 6120 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_317
timestamp 1581320205
transform 1 0 5304 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_318
timestamp 1581320205
transform 1 0 4488 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_319
timestamp 1581320205
transform 1 0 4284 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_320
timestamp 1581320205
transform 1 0 4080 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_321
timestamp 1581320205
transform 1 0 3876 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_322
timestamp 1581320205
transform 1 0 3468 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_323
timestamp 1581320205
transform 1 0 3264 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_324
timestamp 1581320205
transform 1 0 3060 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_325
timestamp 1581320205
transform 1 0 2856 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_326
timestamp 1581320205
transform 1 0 2652 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_327
timestamp 1581320205
transform 1 0 2244 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_328
timestamp 1581320205
transform 1 0 1836 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_329
timestamp 1581320205
transform 1 0 1428 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_330
timestamp 1581320205
transform 1 0 1224 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_331
timestamp 1581320205
transform 1 0 612 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_332
timestamp 1581320205
transform 1 0 12444 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_333
timestamp 1581320205
transform 1 0 12036 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_334
timestamp 1581320205
transform 1 0 11424 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_335
timestamp 1581320205
transform 1 0 11016 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_336
timestamp 1581320205
transform 1 0 10812 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_337
timestamp 1581320205
transform 1 0 10404 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_338
timestamp 1581320205
transform 1 0 9588 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_339
timestamp 1581320205
transform 1 0 9384 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_340
timestamp 1581320205
transform 1 0 8772 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_341
timestamp 1581320205
transform 1 0 8568 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_342
timestamp 1581320205
transform 1 0 8364 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_343
timestamp 1581320205
transform 1 0 8160 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_344
timestamp 1581320205
transform 1 0 7956 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_345
timestamp 1581320205
transform 1 0 7752 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_346
timestamp 1581320205
transform 1 0 7344 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_347
timestamp 1581320205
transform 1 0 7140 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_348
timestamp 1581320205
transform 1 0 6528 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_349
timestamp 1581320205
transform 1 0 6324 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_350
timestamp 1581320205
transform 1 0 5916 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_351
timestamp 1581320205
transform 1 0 5712 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_352
timestamp 1581320205
transform 1 0 5304 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_353
timestamp 1581320205
transform 1 0 5100 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_354
timestamp 1581320205
transform 1 0 4896 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_355
timestamp 1581320205
transform 1 0 4488 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_356
timestamp 1581320205
transform 1 0 4080 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_357
timestamp 1581320205
transform 1 0 3672 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_358
timestamp 1581320205
transform 1 0 3468 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_359
timestamp 1581320205
transform 1 0 3264 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_360
timestamp 1581320205
transform 1 0 3060 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_361
timestamp 1581320205
transform 1 0 2040 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_362
timestamp 1581320205
transform 1 0 1224 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_363
timestamp 1581320205
transform 1 0 1020 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_364
timestamp 1581320205
transform 1 0 612 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_365
timestamp 1581320205
transform 1 0 204 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_366
timestamp 1581320205
transform 1 0 12648 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_367
timestamp 1581320205
transform 1 0 12444 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_368
timestamp 1581320205
transform 1 0 12240 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_369
timestamp 1581320205
transform 1 0 11832 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_370
timestamp 1581320205
transform 1 0 11424 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_371
timestamp 1581320205
transform 1 0 10608 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_372
timestamp 1581320205
transform 1 0 10404 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_373
timestamp 1581320205
transform 1 0 10200 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_374
timestamp 1581320205
transform 1 0 9588 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_375
timestamp 1581320205
transform 1 0 9180 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_376
timestamp 1581320205
transform 1 0 8976 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_377
timestamp 1581320205
transform 1 0 8772 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_378
timestamp 1581320205
transform 1 0 8568 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_379
timestamp 1581320205
transform 1 0 8160 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_380
timestamp 1581320205
transform 1 0 7752 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_381
timestamp 1581320205
transform 1 0 7140 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_382
timestamp 1581320205
transform 1 0 6528 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_383
timestamp 1581320205
transform 1 0 6324 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_384
timestamp 1581320205
transform 1 0 6120 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_385
timestamp 1581320205
transform 1 0 5712 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_386
timestamp 1581320205
transform 1 0 5508 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_387
timestamp 1581320205
transform 1 0 5304 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_388
timestamp 1581320205
transform 1 0 4896 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_389
timestamp 1581320205
transform 1 0 4692 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_390
timestamp 1581320205
transform 1 0 4284 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_391
timestamp 1581320205
transform 1 0 2652 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_392
timestamp 1581320205
transform 1 0 2448 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_393
timestamp 1581320205
transform 1 0 2244 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_394
timestamp 1581320205
transform 1 0 1836 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_395
timestamp 1581320205
transform 1 0 1632 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_396
timestamp 1581320205
transform 1 0 1428 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_397
timestamp 1581320205
transform 1 0 1224 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_398
timestamp 1581320205
transform 1 0 1020 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_399
timestamp 1581320205
transform 1 0 12648 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_400
timestamp 1581320205
transform 1 0 12444 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_401
timestamp 1581320205
transform 1 0 12240 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_402
timestamp 1581320205
transform 1 0 12036 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_403
timestamp 1581320205
transform 1 0 11628 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_404
timestamp 1581320205
transform 1 0 11220 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_405
timestamp 1581320205
transform 1 0 11016 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_406
timestamp 1581320205
transform 1 0 10200 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_407
timestamp 1581320205
transform 1 0 9792 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_408
timestamp 1581320205
transform 1 0 9180 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_409
timestamp 1581320205
transform 1 0 8976 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_410
timestamp 1581320205
transform 1 0 8568 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_411
timestamp 1581320205
transform 1 0 8364 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_412
timestamp 1581320205
transform 1 0 8160 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_413
timestamp 1581320205
transform 1 0 7956 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_414
timestamp 1581320205
transform 1 0 7548 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_415
timestamp 1581320205
transform 1 0 7344 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_416
timestamp 1581320205
transform 1 0 6732 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_417
timestamp 1581320205
transform 1 0 6528 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_418
timestamp 1581320205
transform 1 0 6324 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_419
timestamp 1581320205
transform 1 0 6120 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_420
timestamp 1581320205
transform 1 0 5508 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_421
timestamp 1581320205
transform 1 0 5304 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_422
timestamp 1581320205
transform 1 0 5100 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_423
timestamp 1581320205
transform 1 0 4896 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_424
timestamp 1581320205
transform 1 0 4692 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_425
timestamp 1581320205
transform 1 0 4080 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_426
timestamp 1581320205
transform 1 0 3672 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_427
timestamp 1581320205
transform 1 0 3468 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_428
timestamp 1581320205
transform 1 0 3264 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_429
timestamp 1581320205
transform 1 0 3060 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_430
timestamp 1581320205
transform 1 0 2856 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_431
timestamp 1581320205
transform 1 0 2448 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_432
timestamp 1581320205
transform 1 0 2244 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_433
timestamp 1581320205
transform 1 0 1632 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_434
timestamp 1581320205
transform 1 0 1224 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_435
timestamp 1581320205
transform 1 0 1020 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_436
timestamp 1581320205
transform 1 0 612 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_437
timestamp 1581320205
transform 1 0 12648 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_438
timestamp 1581320205
transform 1 0 12444 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_439
timestamp 1581320205
transform 1 0 12240 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_440
timestamp 1581320205
transform 1 0 12036 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_441
timestamp 1581320205
transform 1 0 11628 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_442
timestamp 1581320205
transform 1 0 10404 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_443
timestamp 1581320205
transform 1 0 9792 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_444
timestamp 1581320205
transform 1 0 9588 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_445
timestamp 1581320205
transform 1 0 9384 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_446
timestamp 1581320205
transform 1 0 9180 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_447
timestamp 1581320205
transform 1 0 8568 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_448
timestamp 1581320205
transform 1 0 8364 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_449
timestamp 1581320205
transform 1 0 7344 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_450
timestamp 1581320205
transform 1 0 7140 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_451
timestamp 1581320205
transform 1 0 6936 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_452
timestamp 1581320205
transform 1 0 6528 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_453
timestamp 1581320205
transform 1 0 6120 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_454
timestamp 1581320205
transform 1 0 5916 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_455
timestamp 1581320205
transform 1 0 5100 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_456
timestamp 1581320205
transform 1 0 4896 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_457
timestamp 1581320205
transform 1 0 4488 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_458
timestamp 1581320205
transform 1 0 3876 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_459
timestamp 1581320205
transform 1 0 3468 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_460
timestamp 1581320205
transform 1 0 3060 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_461
timestamp 1581320205
transform 1 0 2856 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_462
timestamp 1581320205
transform 1 0 1836 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_463
timestamp 1581320205
transform 1 0 1224 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_464
timestamp 1581320205
transform 1 0 1020 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_465
timestamp 1581320205
transform 1 0 816 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_466
timestamp 1581320205
transform 1 0 612 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_467
timestamp 1581320205
transform 1 0 408 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_468
timestamp 1581320205
transform 1 0 204 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_469
timestamp 1581320205
transform 1 0 0 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_470
timestamp 1581320205
transform 1 0 12444 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_471
timestamp 1581320205
transform 1 0 12036 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_472
timestamp 1581320205
transform 1 0 11628 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_473
timestamp 1581320205
transform 1 0 11016 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_474
timestamp 1581320205
transform 1 0 10812 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_475
timestamp 1581320205
transform 1 0 10404 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_476
timestamp 1581320205
transform 1 0 10200 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_477
timestamp 1581320205
transform 1 0 9996 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_478
timestamp 1581320205
transform 1 0 9792 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_479
timestamp 1581320205
transform 1 0 9588 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_480
timestamp 1581320205
transform 1 0 9180 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_481
timestamp 1581320205
transform 1 0 8976 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_482
timestamp 1581320205
transform 1 0 7956 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_483
timestamp 1581320205
transform 1 0 7344 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_484
timestamp 1581320205
transform 1 0 6120 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_485
timestamp 1581320205
transform 1 0 5304 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_486
timestamp 1581320205
transform 1 0 5100 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_487
timestamp 1581320205
transform 1 0 4896 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_488
timestamp 1581320205
transform 1 0 4692 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_489
timestamp 1581320205
transform 1 0 4488 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_490
timestamp 1581320205
transform 1 0 4080 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_491
timestamp 1581320205
transform 1 0 3264 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_492
timestamp 1581320205
transform 1 0 3060 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_493
timestamp 1581320205
transform 1 0 2856 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_494
timestamp 1581320205
transform 1 0 2652 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_495
timestamp 1581320205
transform 1 0 1836 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_496
timestamp 1581320205
transform 1 0 1428 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_497
timestamp 1581320205
transform 1 0 1224 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_498
timestamp 1581320205
transform 1 0 1020 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_499
timestamp 1581320205
transform 1 0 816 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_500
timestamp 1581320205
transform 1 0 408 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_501
timestamp 1581320205
transform 1 0 204 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_502
timestamp 1581320205
transform 1 0 0 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_503
timestamp 1581320205
transform 1 0 12852 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_504
timestamp 1581320205
transform 1 0 12240 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_505
timestamp 1581320205
transform 1 0 11832 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_506
timestamp 1581320205
transform 1 0 11220 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_507
timestamp 1581320205
transform 1 0 11016 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_508
timestamp 1581320205
transform 1 0 10404 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_509
timestamp 1581320205
transform 1 0 9588 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_510
timestamp 1581320205
transform 1 0 9384 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_511
timestamp 1581320205
transform 1 0 9180 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_512
timestamp 1581320205
transform 1 0 8568 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_513
timestamp 1581320205
transform 1 0 7752 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_514
timestamp 1581320205
transform 1 0 7140 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_515
timestamp 1581320205
transform 1 0 6732 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_516
timestamp 1581320205
transform 1 0 6528 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_517
timestamp 1581320205
transform 1 0 6120 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_518
timestamp 1581320205
transform 1 0 5712 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_519
timestamp 1581320205
transform 1 0 5508 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_520
timestamp 1581320205
transform 1 0 5304 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_521
timestamp 1581320205
transform 1 0 4896 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_522
timestamp 1581320205
transform 1 0 4284 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_523
timestamp 1581320205
transform 1 0 3876 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_524
timestamp 1581320205
transform 1 0 3672 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_525
timestamp 1581320205
transform 1 0 3060 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_526
timestamp 1581320205
transform 1 0 2856 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_527
timestamp 1581320205
transform 1 0 2652 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_528
timestamp 1581320205
transform 1 0 2448 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_529
timestamp 1581320205
transform 1 0 2244 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_530
timestamp 1581320205
transform 1 0 2040 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_531
timestamp 1581320205
transform 1 0 1836 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_532
timestamp 1581320205
transform 1 0 1632 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_533
timestamp 1581320205
transform 1 0 1428 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_534
timestamp 1581320205
transform 1 0 1224 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_535
timestamp 1581320205
transform 1 0 1020 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_536
timestamp 1581320205
transform 1 0 816 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_537
timestamp 1581320205
transform 1 0 408 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_538
timestamp 1581320205
transform 1 0 0 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_539
timestamp 1581320205
transform 1 0 12240 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_540
timestamp 1581320205
transform 1 0 11628 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_541
timestamp 1581320205
transform 1 0 11424 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_542
timestamp 1581320205
transform 1 0 11016 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_543
timestamp 1581320205
transform 1 0 10812 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_544
timestamp 1581320205
transform 1 0 10608 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_545
timestamp 1581320205
transform 1 0 10404 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_546
timestamp 1581320205
transform 1 0 9384 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_547
timestamp 1581320205
transform 1 0 9180 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_548
timestamp 1581320205
transform 1 0 8772 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_549
timestamp 1581320205
transform 1 0 8568 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_550
timestamp 1581320205
transform 1 0 8364 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_551
timestamp 1581320205
transform 1 0 7956 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_552
timestamp 1581320205
transform 1 0 7344 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_553
timestamp 1581320205
transform 1 0 7140 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_554
timestamp 1581320205
transform 1 0 6936 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_555
timestamp 1581320205
transform 1 0 6528 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_556
timestamp 1581320205
transform 1 0 6324 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_557
timestamp 1581320205
transform 1 0 6120 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_558
timestamp 1581320205
transform 1 0 5916 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_559
timestamp 1581320205
transform 1 0 5304 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_560
timestamp 1581320205
transform 1 0 5100 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_561
timestamp 1581320205
transform 1 0 4896 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_562
timestamp 1581320205
transform 1 0 4080 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_563
timestamp 1581320205
transform 1 0 3876 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_564
timestamp 1581320205
transform 1 0 3468 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_565
timestamp 1581320205
transform 1 0 3264 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_566
timestamp 1581320205
transform 1 0 2856 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_567
timestamp 1581320205
transform 1 0 2652 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_568
timestamp 1581320205
transform 1 0 2448 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_569
timestamp 1581320205
transform 1 0 1632 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_570
timestamp 1581320205
transform 1 0 1428 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_571
timestamp 1581320205
transform 1 0 1224 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_572
timestamp 1581320205
transform 1 0 1020 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_573
timestamp 1581320205
transform 1 0 816 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_574
timestamp 1581320205
transform 1 0 612 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_575
timestamp 1581320205
transform 1 0 408 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_576
timestamp 1581320205
transform 1 0 0 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_577
timestamp 1581320205
transform 1 0 11628 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_578
timestamp 1581320205
transform 1 0 11424 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_579
timestamp 1581320205
transform 1 0 11016 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_580
timestamp 1581320205
transform 1 0 10608 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_581
timestamp 1581320205
transform 1 0 9996 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_582
timestamp 1581320205
transform 1 0 9384 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_583
timestamp 1581320205
transform 1 0 8772 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_584
timestamp 1581320205
transform 1 0 8568 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_585
timestamp 1581320205
transform 1 0 8364 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_586
timestamp 1581320205
transform 1 0 7956 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_587
timestamp 1581320205
transform 1 0 7752 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_588
timestamp 1581320205
transform 1 0 7548 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_589
timestamp 1581320205
transform 1 0 7344 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_590
timestamp 1581320205
transform 1 0 7140 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_591
timestamp 1581320205
transform 1 0 6732 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_592
timestamp 1581320205
transform 1 0 6528 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_593
timestamp 1581320205
transform 1 0 6324 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_594
timestamp 1581320205
transform 1 0 5916 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_595
timestamp 1581320205
transform 1 0 5304 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_596
timestamp 1581320205
transform 1 0 5100 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_597
timestamp 1581320205
transform 1 0 4896 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_598
timestamp 1581320205
transform 1 0 4692 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_599
timestamp 1581320205
transform 1 0 4488 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_600
timestamp 1581320205
transform 1 0 4080 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_601
timestamp 1581320205
transform 1 0 3672 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_602
timestamp 1581320205
transform 1 0 3264 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_603
timestamp 1581320205
transform 1 0 2856 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_604
timestamp 1581320205
transform 1 0 2652 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_605
timestamp 1581320205
transform 1 0 2040 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_606
timestamp 1581320205
transform 1 0 1428 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_607
timestamp 1581320205
transform 1 0 408 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_608
timestamp 1581320205
transform 1 0 12036 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_609
timestamp 1581320205
transform 1 0 11424 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_610
timestamp 1581320205
transform 1 0 10812 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_611
timestamp 1581320205
transform 1 0 10404 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_612
timestamp 1581320205
transform 1 0 9792 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_613
timestamp 1581320205
transform 1 0 9180 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_614
timestamp 1581320205
transform 1 0 8772 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_615
timestamp 1581320205
transform 1 0 8364 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_616
timestamp 1581320205
transform 1 0 8160 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_617
timestamp 1581320205
transform 1 0 7956 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_618
timestamp 1581320205
transform 1 0 6936 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_619
timestamp 1581320205
transform 1 0 6732 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_620
timestamp 1581320205
transform 1 0 6528 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_621
timestamp 1581320205
transform 1 0 6324 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_622
timestamp 1581320205
transform 1 0 5508 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_623
timestamp 1581320205
transform 1 0 5304 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_624
timestamp 1581320205
transform 1 0 5100 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_625
timestamp 1581320205
transform 1 0 4692 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_626
timestamp 1581320205
transform 1 0 4284 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_627
timestamp 1581320205
transform 1 0 3876 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_628
timestamp 1581320205
transform 1 0 3468 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_629
timestamp 1581320205
transform 1 0 2448 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_630
timestamp 1581320205
transform 1 0 2040 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_631
timestamp 1581320205
transform 1 0 1836 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_632
timestamp 1581320205
transform 1 0 1632 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_633
timestamp 1581320205
transform 1 0 1224 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_634
timestamp 1581320205
transform 1 0 1020 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_635
timestamp 1581320205
transform 1 0 408 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_636
timestamp 1581320205
transform 1 0 204 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_637
timestamp 1581320205
transform 1 0 12648 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_638
timestamp 1581320205
transform 1 0 12240 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_639
timestamp 1581320205
transform 1 0 12036 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_640
timestamp 1581320205
transform 1 0 11628 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_641
timestamp 1581320205
transform 1 0 11424 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_642
timestamp 1581320205
transform 1 0 11220 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_643
timestamp 1581320205
transform 1 0 10812 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_644
timestamp 1581320205
transform 1 0 10608 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_645
timestamp 1581320205
transform 1 0 10200 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_646
timestamp 1581320205
transform 1 0 9792 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_647
timestamp 1581320205
transform 1 0 9180 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_648
timestamp 1581320205
transform 1 0 8976 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_649
timestamp 1581320205
transform 1 0 8772 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_650
timestamp 1581320205
transform 1 0 8568 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_651
timestamp 1581320205
transform 1 0 8160 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_652
timestamp 1581320205
transform 1 0 7752 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_653
timestamp 1581320205
transform 1 0 7548 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_654
timestamp 1581320205
transform 1 0 7140 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_655
timestamp 1581320205
transform 1 0 6936 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_656
timestamp 1581320205
transform 1 0 6324 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_657
timestamp 1581320205
transform 1 0 6120 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_658
timestamp 1581320205
transform 1 0 5712 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_659
timestamp 1581320205
transform 1 0 4488 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_660
timestamp 1581320205
transform 1 0 3876 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_661
timestamp 1581320205
transform 1 0 3672 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_662
timestamp 1581320205
transform 1 0 3264 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_663
timestamp 1581320205
transform 1 0 2652 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_664
timestamp 1581320205
transform 1 0 2448 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_665
timestamp 1581320205
transform 1 0 1836 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_666
timestamp 1581320205
transform 1 0 1632 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_667
timestamp 1581320205
transform 1 0 1428 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_668
timestamp 1581320205
transform 1 0 1020 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_669
timestamp 1581320205
transform 1 0 612 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_670
timestamp 1581320205
transform 1 0 408 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_671
timestamp 1581320205
transform 1 0 204 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_672
timestamp 1581320205
transform 1 0 12852 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_673
timestamp 1581320205
transform 1 0 12648 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_674
timestamp 1581320205
transform 1 0 12240 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_675
timestamp 1581320205
transform 1 0 12036 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_676
timestamp 1581320205
transform 1 0 11628 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_677
timestamp 1581320205
transform 1 0 11424 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_678
timestamp 1581320205
transform 1 0 11016 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_679
timestamp 1581320205
transform 1 0 10812 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_680
timestamp 1581320205
transform 1 0 10404 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_681
timestamp 1581320205
transform 1 0 10200 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_682
timestamp 1581320205
transform 1 0 9996 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_683
timestamp 1581320205
transform 1 0 9792 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_684
timestamp 1581320205
transform 1 0 9588 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_685
timestamp 1581320205
transform 1 0 9384 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_686
timestamp 1581320205
transform 1 0 9180 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_687
timestamp 1581320205
transform 1 0 8568 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_688
timestamp 1581320205
transform 1 0 8364 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_689
timestamp 1581320205
transform 1 0 7344 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_690
timestamp 1581320205
transform 1 0 6732 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_691
timestamp 1581320205
transform 1 0 6120 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_692
timestamp 1581320205
transform 1 0 5304 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_693
timestamp 1581320205
transform 1 0 4692 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_694
timestamp 1581320205
transform 1 0 4488 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_695
timestamp 1581320205
transform 1 0 3876 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_696
timestamp 1581320205
transform 1 0 3264 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_697
timestamp 1581320205
transform 1 0 2856 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_698
timestamp 1581320205
transform 1 0 2040 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_699
timestamp 1581320205
transform 1 0 1836 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_700
timestamp 1581320205
transform 1 0 816 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_701
timestamp 1581320205
transform 1 0 0 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_702
timestamp 1581320205
transform 1 0 12852 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_703
timestamp 1581320205
transform 1 0 12648 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_704
timestamp 1581320205
transform 1 0 12444 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_705
timestamp 1581320205
transform 1 0 12240 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_706
timestamp 1581320205
transform 1 0 11832 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_707
timestamp 1581320205
transform 1 0 11016 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_708
timestamp 1581320205
transform 1 0 10812 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_709
timestamp 1581320205
transform 1 0 10200 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_710
timestamp 1581320205
transform 1 0 9996 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_711
timestamp 1581320205
transform 1 0 9792 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_712
timestamp 1581320205
transform 1 0 9588 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_713
timestamp 1581320205
transform 1 0 8976 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_714
timestamp 1581320205
transform 1 0 8364 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_715
timestamp 1581320205
transform 1 0 7752 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_716
timestamp 1581320205
transform 1 0 7548 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_717
timestamp 1581320205
transform 1 0 6324 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_718
timestamp 1581320205
transform 1 0 6120 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_719
timestamp 1581320205
transform 1 0 5712 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_720
timestamp 1581320205
transform 1 0 5508 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_721
timestamp 1581320205
transform 1 0 5304 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_722
timestamp 1581320205
transform 1 0 5100 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_723
timestamp 1581320205
transform 1 0 4896 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_724
timestamp 1581320205
transform 1 0 4488 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_725
timestamp 1581320205
transform 1 0 4080 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_726
timestamp 1581320205
transform 1 0 3060 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_727
timestamp 1581320205
transform 1 0 2856 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_728
timestamp 1581320205
transform 1 0 2040 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_729
timestamp 1581320205
transform 1 0 1632 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_730
timestamp 1581320205
transform 1 0 1020 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_731
timestamp 1581320205
transform 1 0 816 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_732
timestamp 1581320205
transform 1 0 612 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_733
timestamp 1581320205
transform 1 0 408 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_734
timestamp 1581320205
transform 1 0 0 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_735
timestamp 1581320205
transform 1 0 12852 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_736
timestamp 1581320205
transform 1 0 12444 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_737
timestamp 1581320205
transform 1 0 12240 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_738
timestamp 1581320205
transform 1 0 12036 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_739
timestamp 1581320205
transform 1 0 11220 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_740
timestamp 1581320205
transform 1 0 11016 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_741
timestamp 1581320205
transform 1 0 10812 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_742
timestamp 1581320205
transform 1 0 10608 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_743
timestamp 1581320205
transform 1 0 10200 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_744
timestamp 1581320205
transform 1 0 9996 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_745
timestamp 1581320205
transform 1 0 9384 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_746
timestamp 1581320205
transform 1 0 8364 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_747
timestamp 1581320205
transform 1 0 7752 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_748
timestamp 1581320205
transform 1 0 7344 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_749
timestamp 1581320205
transform 1 0 7140 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_750
timestamp 1581320205
transform 1 0 6732 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_751
timestamp 1581320205
transform 1 0 6324 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_752
timestamp 1581320205
transform 1 0 6120 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_753
timestamp 1581320205
transform 1 0 5916 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_754
timestamp 1581320205
transform 1 0 5712 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_755
timestamp 1581320205
transform 1 0 5508 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_756
timestamp 1581320205
transform 1 0 5100 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_757
timestamp 1581320205
transform 1 0 4896 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_758
timestamp 1581320205
transform 1 0 4692 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_759
timestamp 1581320205
transform 1 0 4284 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_760
timestamp 1581320205
transform 1 0 3876 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_761
timestamp 1581320205
transform 1 0 3672 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_762
timestamp 1581320205
transform 1 0 3468 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_763
timestamp 1581320205
transform 1 0 3264 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_764
timestamp 1581320205
transform 1 0 2856 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_765
timestamp 1581320205
transform 1 0 2652 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_766
timestamp 1581320205
transform 1 0 2448 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_767
timestamp 1581320205
transform 1 0 2040 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_768
timestamp 1581320205
transform 1 0 1632 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_769
timestamp 1581320205
transform 1 0 1020 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_770
timestamp 1581320205
transform 1 0 816 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_771
timestamp 1581320205
transform 1 0 0 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_772
timestamp 1581320205
transform 1 0 12852 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_773
timestamp 1581320205
transform 1 0 12444 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_774
timestamp 1581320205
transform 1 0 11424 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_775
timestamp 1581320205
transform 1 0 10404 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_776
timestamp 1581320205
transform 1 0 10200 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_777
timestamp 1581320205
transform 1 0 9792 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_778
timestamp 1581320205
transform 1 0 8772 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_779
timestamp 1581320205
transform 1 0 8568 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_780
timestamp 1581320205
transform 1 0 8364 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_781
timestamp 1581320205
transform 1 0 7956 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_782
timestamp 1581320205
transform 1 0 7752 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_783
timestamp 1581320205
transform 1 0 7140 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_784
timestamp 1581320205
transform 1 0 6528 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_785
timestamp 1581320205
transform 1 0 6324 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_786
timestamp 1581320205
transform 1 0 6120 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_787
timestamp 1581320205
transform 1 0 5712 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_788
timestamp 1581320205
transform 1 0 5508 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_789
timestamp 1581320205
transform 1 0 5304 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_790
timestamp 1581320205
transform 1 0 4896 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_791
timestamp 1581320205
transform 1 0 4692 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_792
timestamp 1581320205
transform 1 0 4488 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_793
timestamp 1581320205
transform 1 0 3876 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_794
timestamp 1581320205
transform 1 0 3468 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_795
timestamp 1581320205
transform 1 0 3060 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_796
timestamp 1581320205
transform 1 0 2652 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_797
timestamp 1581320205
transform 1 0 1836 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_798
timestamp 1581320205
transform 1 0 1224 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_799
timestamp 1581320205
transform 1 0 408 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_800
timestamp 1581320205
transform 1 0 12852 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_801
timestamp 1581320205
transform 1 0 11832 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_802
timestamp 1581320205
transform 1 0 11628 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_803
timestamp 1581320205
transform 1 0 11220 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_804
timestamp 1581320205
transform 1 0 11016 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_805
timestamp 1581320205
transform 1 0 10608 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_806
timestamp 1581320205
transform 1 0 9996 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_807
timestamp 1581320205
transform 1 0 9384 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_808
timestamp 1581320205
transform 1 0 9180 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_809
timestamp 1581320205
transform 1 0 8976 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_810
timestamp 1581320205
transform 1 0 8160 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_811
timestamp 1581320205
transform 1 0 7956 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_812
timestamp 1581320205
transform 1 0 7752 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_813
timestamp 1581320205
transform 1 0 7344 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_814
timestamp 1581320205
transform 1 0 7140 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_815
timestamp 1581320205
transform 1 0 6936 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_816
timestamp 1581320205
transform 1 0 5712 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_817
timestamp 1581320205
transform 1 0 5508 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_818
timestamp 1581320205
transform 1 0 5304 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_819
timestamp 1581320205
transform 1 0 4284 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_820
timestamp 1581320205
transform 1 0 4080 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_821
timestamp 1581320205
transform 1 0 3672 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_822
timestamp 1581320205
transform 1 0 3468 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_823
timestamp 1581320205
transform 1 0 3264 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_824
timestamp 1581320205
transform 1 0 2652 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_825
timestamp 1581320205
transform 1 0 2244 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_826
timestamp 1581320205
transform 1 0 2040 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_827
timestamp 1581320205
transform 1 0 1632 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_828
timestamp 1581320205
transform 1 0 1428 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_829
timestamp 1581320205
transform 1 0 408 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_830
timestamp 1581320205
transform 1 0 12852 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_831
timestamp 1581320205
transform 1 0 12444 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_832
timestamp 1581320205
transform 1 0 12240 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_833
timestamp 1581320205
transform 1 0 12036 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_834
timestamp 1581320205
transform 1 0 11628 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_835
timestamp 1581320205
transform 1 0 11424 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_836
timestamp 1581320205
transform 1 0 11016 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_837
timestamp 1581320205
transform 1 0 10608 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_838
timestamp 1581320205
transform 1 0 10404 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_839
timestamp 1581320205
transform 1 0 10200 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_840
timestamp 1581320205
transform 1 0 9384 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_841
timestamp 1581320205
transform 1 0 8976 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_842
timestamp 1581320205
transform 1 0 8160 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_843
timestamp 1581320205
transform 1 0 7752 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_844
timestamp 1581320205
transform 1 0 7344 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_845
timestamp 1581320205
transform 1 0 7140 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_846
timestamp 1581320205
transform 1 0 6528 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_847
timestamp 1581320205
transform 1 0 5712 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_848
timestamp 1581320205
transform 1 0 4284 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_849
timestamp 1581320205
transform 1 0 4080 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_850
timestamp 1581320205
transform 1 0 3672 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_851
timestamp 1581320205
transform 1 0 2856 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_852
timestamp 1581320205
transform 1 0 2448 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_853
timestamp 1581320205
transform 1 0 1836 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_854
timestamp 1581320205
transform 1 0 612 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_855
timestamp 1581320205
transform 1 0 408 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_856
timestamp 1581320205
transform 1 0 0 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_857
timestamp 1581320205
transform 1 0 12444 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_858
timestamp 1581320205
transform 1 0 12036 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_859
timestamp 1581320205
transform 1 0 11424 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_860
timestamp 1581320205
transform 1 0 11016 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_861
timestamp 1581320205
transform 1 0 10812 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_862
timestamp 1581320205
transform 1 0 10608 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_863
timestamp 1581320205
transform 1 0 10200 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_864
timestamp 1581320205
transform 1 0 9996 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_865
timestamp 1581320205
transform 1 0 9792 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_866
timestamp 1581320205
transform 1 0 9588 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_867
timestamp 1581320205
transform 1 0 8364 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_868
timestamp 1581320205
transform 1 0 7956 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_869
timestamp 1581320205
transform 1 0 7344 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_870
timestamp 1581320205
transform 1 0 6936 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_871
timestamp 1581320205
transform 1 0 6732 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_872
timestamp 1581320205
transform 1 0 6528 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_873
timestamp 1581320205
transform 1 0 6324 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_874
timestamp 1581320205
transform 1 0 5916 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_875
timestamp 1581320205
transform 1 0 5304 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_876
timestamp 1581320205
transform 1 0 4896 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_877
timestamp 1581320205
transform 1 0 4692 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_878
timestamp 1581320205
transform 1 0 4284 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_879
timestamp 1581320205
transform 1 0 4080 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_880
timestamp 1581320205
transform 1 0 3672 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_881
timestamp 1581320205
transform 1 0 2652 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_882
timestamp 1581320205
transform 1 0 2244 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_883
timestamp 1581320205
transform 1 0 2040 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_884
timestamp 1581320205
transform 1 0 1836 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_885
timestamp 1581320205
transform 1 0 1632 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_886
timestamp 1581320205
transform 1 0 1224 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_887
timestamp 1581320205
transform 1 0 1020 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_888
timestamp 1581320205
transform 1 0 816 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_889
timestamp 1581320205
transform 1 0 204 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_890
timestamp 1581320205
transform 1 0 0 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_891
timestamp 1581320205
transform 1 0 12240 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_892
timestamp 1581320205
transform 1 0 12036 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_893
timestamp 1581320205
transform 1 0 11832 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_894
timestamp 1581320205
transform 1 0 11424 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_895
timestamp 1581320205
transform 1 0 11220 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_896
timestamp 1581320205
transform 1 0 10404 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_897
timestamp 1581320205
transform 1 0 9792 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_898
timestamp 1581320205
transform 1 0 9588 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_899
timestamp 1581320205
transform 1 0 9384 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_900
timestamp 1581320205
transform 1 0 9180 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_901
timestamp 1581320205
transform 1 0 8976 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_902
timestamp 1581320205
transform 1 0 8772 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_903
timestamp 1581320205
transform 1 0 8568 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_904
timestamp 1581320205
transform 1 0 8160 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_905
timestamp 1581320205
transform 1 0 7956 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_906
timestamp 1581320205
transform 1 0 7548 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_907
timestamp 1581320205
transform 1 0 7344 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_908
timestamp 1581320205
transform 1 0 6732 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_909
timestamp 1581320205
transform 1 0 6324 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_910
timestamp 1581320205
transform 1 0 5916 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_911
timestamp 1581320205
transform 1 0 5304 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_912
timestamp 1581320205
transform 1 0 5100 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_913
timestamp 1581320205
transform 1 0 4692 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_914
timestamp 1581320205
transform 1 0 4488 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_915
timestamp 1581320205
transform 1 0 4284 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_916
timestamp 1581320205
transform 1 0 4080 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_917
timestamp 1581320205
transform 1 0 3876 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_918
timestamp 1581320205
transform 1 0 3468 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_919
timestamp 1581320205
transform 1 0 3264 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_920
timestamp 1581320205
transform 1 0 3060 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_921
timestamp 1581320205
transform 1 0 2652 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_922
timestamp 1581320205
transform 1 0 2448 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_923
timestamp 1581320205
transform 1 0 2244 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_924
timestamp 1581320205
transform 1 0 2040 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_925
timestamp 1581320205
transform 1 0 1836 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_926
timestamp 1581320205
transform 1 0 1428 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_927
timestamp 1581320205
transform 1 0 1224 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_928
timestamp 1581320205
transform 1 0 816 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_929
timestamp 1581320205
transform 1 0 204 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_930
timestamp 1581320205
transform 1 0 12648 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_931
timestamp 1581320205
transform 1 0 12444 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_932
timestamp 1581320205
transform 1 0 12036 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_933
timestamp 1581320205
transform 1 0 11832 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_934
timestamp 1581320205
transform 1 0 11424 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_935
timestamp 1581320205
transform 1 0 11220 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_936
timestamp 1581320205
transform 1 0 10812 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_937
timestamp 1581320205
transform 1 0 10404 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_938
timestamp 1581320205
transform 1 0 8976 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_939
timestamp 1581320205
transform 1 0 8568 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_940
timestamp 1581320205
transform 1 0 8160 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_941
timestamp 1581320205
transform 1 0 7956 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_942
timestamp 1581320205
transform 1 0 7140 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_943
timestamp 1581320205
transform 1 0 6936 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_944
timestamp 1581320205
transform 1 0 6528 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_945
timestamp 1581320205
transform 1 0 5712 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_946
timestamp 1581320205
transform 1 0 5508 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_947
timestamp 1581320205
transform 1 0 5304 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_948
timestamp 1581320205
transform 1 0 4692 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_949
timestamp 1581320205
transform 1 0 4488 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_950
timestamp 1581320205
transform 1 0 4284 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_951
timestamp 1581320205
transform 1 0 3672 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_952
timestamp 1581320205
transform 1 0 3264 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_953
timestamp 1581320205
transform 1 0 2652 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_954
timestamp 1581320205
transform 1 0 2448 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_955
timestamp 1581320205
transform 1 0 2244 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_956
timestamp 1581320205
transform 1 0 2040 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_957
timestamp 1581320205
transform 1 0 1836 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_958
timestamp 1581320205
transform 1 0 1632 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_959
timestamp 1581320205
transform 1 0 1224 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_960
timestamp 1581320205
transform 1 0 1020 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_961
timestamp 1581320205
transform 1 0 204 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_962
timestamp 1581320205
transform 1 0 11832 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_963
timestamp 1581320205
transform 1 0 11628 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_964
timestamp 1581320205
transform 1 0 11220 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_965
timestamp 1581320205
transform 1 0 11016 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_966
timestamp 1581320205
transform 1 0 10812 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_967
timestamp 1581320205
transform 1 0 10608 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_968
timestamp 1581320205
transform 1 0 9792 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_969
timestamp 1581320205
transform 1 0 9588 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_970
timestamp 1581320205
transform 1 0 9384 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_971
timestamp 1581320205
transform 1 0 9180 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_972
timestamp 1581320205
transform 1 0 8976 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_973
timestamp 1581320205
transform 1 0 8772 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_974
timestamp 1581320205
transform 1 0 8568 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_975
timestamp 1581320205
transform 1 0 8160 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_976
timestamp 1581320205
transform 1 0 7956 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_977
timestamp 1581320205
transform 1 0 7752 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_978
timestamp 1581320205
transform 1 0 7548 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_979
timestamp 1581320205
transform 1 0 6936 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_980
timestamp 1581320205
transform 1 0 6732 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_981
timestamp 1581320205
transform 1 0 5304 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_982
timestamp 1581320205
transform 1 0 4488 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_983
timestamp 1581320205
transform 1 0 4080 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_984
timestamp 1581320205
transform 1 0 3876 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_985
timestamp 1581320205
transform 1 0 3672 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_986
timestamp 1581320205
transform 1 0 3468 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_987
timestamp 1581320205
transform 1 0 2856 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_988
timestamp 1581320205
transform 1 0 1632 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_989
timestamp 1581320205
transform 1 0 1224 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_990
timestamp 1581320205
transform 1 0 816 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_991
timestamp 1581320205
transform 1 0 612 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_992
timestamp 1581320205
transform 1 0 204 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_993
timestamp 1581320205
transform 1 0 0 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_994
timestamp 1581320205
transform 1 0 11628 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_995
timestamp 1581320205
transform 1 0 11220 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_996
timestamp 1581320205
transform 1 0 10812 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_997
timestamp 1581320205
transform 1 0 10608 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_998
timestamp 1581320205
transform 1 0 9996 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_999
timestamp 1581320205
transform 1 0 9792 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1000
timestamp 1581320205
transform 1 0 9384 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1001
timestamp 1581320205
transform 1 0 8976 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1002
timestamp 1581320205
transform 1 0 8568 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1003
timestamp 1581320205
transform 1 0 8364 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1004
timestamp 1581320205
transform 1 0 7956 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1005
timestamp 1581320205
transform 1 0 7548 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1006
timestamp 1581320205
transform 1 0 6732 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1007
timestamp 1581320205
transform 1 0 6528 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1008
timestamp 1581320205
transform 1 0 6324 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1009
timestamp 1581320205
transform 1 0 5712 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1010
timestamp 1581320205
transform 1 0 5508 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1011
timestamp 1581320205
transform 1 0 5100 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1012
timestamp 1581320205
transform 1 0 4488 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1013
timestamp 1581320205
transform 1 0 3876 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1014
timestamp 1581320205
transform 1 0 3468 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1015
timestamp 1581320205
transform 1 0 3060 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1016
timestamp 1581320205
transform 1 0 2652 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1017
timestamp 1581320205
transform 1 0 1632 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1018
timestamp 1581320205
transform 1 0 12648 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1019
timestamp 1581320205
transform 1 0 12036 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1020
timestamp 1581320205
transform 1 0 11628 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1021
timestamp 1581320205
transform 1 0 11424 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1022
timestamp 1581320205
transform 1 0 11220 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1023
timestamp 1581320205
transform 1 0 11016 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1024
timestamp 1581320205
transform 1 0 10608 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1025
timestamp 1581320205
transform 1 0 10404 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1026
timestamp 1581320205
transform 1 0 9588 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1027
timestamp 1581320205
transform 1 0 8976 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1028
timestamp 1581320205
transform 1 0 8772 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1029
timestamp 1581320205
transform 1 0 8364 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1030
timestamp 1581320205
transform 1 0 8160 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1031
timestamp 1581320205
transform 1 0 7956 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1032
timestamp 1581320205
transform 1 0 7752 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1033
timestamp 1581320205
transform 1 0 7548 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1034
timestamp 1581320205
transform 1 0 7344 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1035
timestamp 1581320205
transform 1 0 6528 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1036
timestamp 1581320205
transform 1 0 6120 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1037
timestamp 1581320205
transform 1 0 5304 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1038
timestamp 1581320205
transform 1 0 5100 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1039
timestamp 1581320205
transform 1 0 4896 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1040
timestamp 1581320205
transform 1 0 4692 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1041
timestamp 1581320205
transform 1 0 4488 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1042
timestamp 1581320205
transform 1 0 3876 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1043
timestamp 1581320205
transform 1 0 3468 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1044
timestamp 1581320205
transform 1 0 3264 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1045
timestamp 1581320205
transform 1 0 3060 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1046
timestamp 1581320205
transform 1 0 2652 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1047
timestamp 1581320205
transform 1 0 2244 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1048
timestamp 1581320205
transform 1 0 2040 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1049
timestamp 1581320205
transform 1 0 1836 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1050
timestamp 1581320205
transform 1 0 1224 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1051
timestamp 1581320205
transform 1 0 1020 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1052
timestamp 1581320205
transform 1 0 816 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1053
timestamp 1581320205
transform 1 0 408 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1054
timestamp 1581320205
transform 1 0 0 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_0
timestamp 1581320205
transform 1 0 13056 0 1 7817
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_1
timestamp 1581320205
transform 1 0 11424 0 1 7817
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_2
timestamp 1581320205
transform 1 0 9792 0 1 7817
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_3
timestamp 1581320205
transform 1 0 8160 0 1 7817
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_4
timestamp 1581320205
transform 1 0 6528 0 1 7817
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_5
timestamp 1581320205
transform 1 0 4896 0 1 7817
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_6
timestamp 1581320205
transform 1 0 3264 0 1 7817
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_7
timestamp 1581320205
transform 1 0 1632 0 1 7817
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_8
timestamp 1581320205
transform 1 0 0 0 1 7817
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_9
timestamp 1581320205
transform 1 0 13056 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_10
timestamp 1581320205
transform 1 0 11424 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_11
timestamp 1581320205
transform 1 0 9792 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_12
timestamp 1581320205
transform 1 0 8160 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_13
timestamp 1581320205
transform 1 0 6528 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_14
timestamp 1581320205
transform 1 0 4896 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_15
timestamp 1581320205
transform 1 0 3264 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_16
timestamp 1581320205
transform 1 0 1632 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_17
timestamp 1581320205
transform 1 0 0 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_18
timestamp 1581320205
transform 1 0 13056 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_19
timestamp 1581320205
transform 1 0 11424 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_20
timestamp 1581320205
transform 1 0 9792 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_21
timestamp 1581320205
transform 1 0 8160 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_22
timestamp 1581320205
transform 1 0 6528 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_23
timestamp 1581320205
transform 1 0 4896 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_24
timestamp 1581320205
transform 1 0 3264 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_25
timestamp 1581320205
transform 1 0 1632 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_26
timestamp 1581320205
transform 1 0 0 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_27
timestamp 1581320205
transform 1 0 13056 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_28
timestamp 1581320205
transform 1 0 11424 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_29
timestamp 1581320205
transform 1 0 9792 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_30
timestamp 1581320205
transform 1 0 8160 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_31
timestamp 1581320205
transform 1 0 6528 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_32
timestamp 1581320205
transform 1 0 4896 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_33
timestamp 1581320205
transform 1 0 3264 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_34
timestamp 1581320205
transform 1 0 1632 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_35
timestamp 1581320205
transform 1 0 0 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_36
timestamp 1581320205
transform 1 0 13056 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_37
timestamp 1581320205
transform 1 0 11424 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_38
timestamp 1581320205
transform 1 0 9792 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_39
timestamp 1581320205
transform 1 0 8160 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_40
timestamp 1581320205
transform 1 0 6528 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_41
timestamp 1581320205
transform 1 0 4896 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_42
timestamp 1581320205
transform 1 0 3264 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_43
timestamp 1581320205
transform 1 0 1632 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_44
timestamp 1581320205
transform 1 0 0 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_45
timestamp 1581320205
transform 1 0 13056 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_46
timestamp 1581320205
transform 1 0 11424 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_47
timestamp 1581320205
transform 1 0 9792 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_48
timestamp 1581320205
transform 1 0 8160 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_49
timestamp 1581320205
transform 1 0 6528 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_50
timestamp 1581320205
transform 1 0 4896 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_51
timestamp 1581320205
transform 1 0 3264 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_52
timestamp 1581320205
transform 1 0 1632 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_53
timestamp 1581320205
transform 1 0 0 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_54
timestamp 1581320205
transform 1 0 13056 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_55
timestamp 1581320205
transform 1 0 11424 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_56
timestamp 1581320205
transform 1 0 9792 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_57
timestamp 1581320205
transform 1 0 8160 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_58
timestamp 1581320205
transform 1 0 6528 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_59
timestamp 1581320205
transform 1 0 4896 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_60
timestamp 1581320205
transform 1 0 3264 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_61
timestamp 1581320205
transform 1 0 1632 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_62
timestamp 1581320205
transform 1 0 0 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_63
timestamp 1581320205
transform 1 0 13056 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_64
timestamp 1581320205
transform 1 0 11424 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_65
timestamp 1581320205
transform 1 0 9792 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_66
timestamp 1581320205
transform 1 0 8160 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_67
timestamp 1581320205
transform 1 0 6528 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_68
timestamp 1581320205
transform 1 0 4896 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_69
timestamp 1581320205
transform 1 0 3264 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_70
timestamp 1581320205
transform 1 0 1632 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_71
timestamp 1581320205
transform 1 0 0 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_72
timestamp 1581320205
transform 1 0 13056 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_73
timestamp 1581320205
transform 1 0 11424 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_74
timestamp 1581320205
transform 1 0 9792 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_75
timestamp 1581320205
transform 1 0 8160 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_76
timestamp 1581320205
transform 1 0 6528 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_77
timestamp 1581320205
transform 1 0 4896 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_78
timestamp 1581320205
transform 1 0 3264 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_79
timestamp 1581320205
transform 1 0 1632 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_80
timestamp 1581320205
transform 1 0 0 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_81
timestamp 1581320205
transform 1 0 13056 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_82
timestamp 1581320205
transform 1 0 11424 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_83
timestamp 1581320205
transform 1 0 9792 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_84
timestamp 1581320205
transform 1 0 8160 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_85
timestamp 1581320205
transform 1 0 6528 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_86
timestamp 1581320205
transform 1 0 4896 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_87
timestamp 1581320205
transform 1 0 3264 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_88
timestamp 1581320205
transform 1 0 1632 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_89
timestamp 1581320205
transform 1 0 0 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_90
timestamp 1581320205
transform 1 0 13056 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_91
timestamp 1581320205
transform 1 0 11424 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_92
timestamp 1581320205
transform 1 0 9792 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_93
timestamp 1581320205
transform 1 0 8160 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_94
timestamp 1581320205
transform 1 0 6528 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_95
timestamp 1581320205
transform 1 0 4896 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_96
timestamp 1581320205
transform 1 0 3264 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_97
timestamp 1581320205
transform 1 0 1632 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_98
timestamp 1581320205
transform 1 0 0 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_99
timestamp 1581320205
transform 1 0 13056 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_100
timestamp 1581320205
transform 1 0 11424 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_101
timestamp 1581320205
transform 1 0 9792 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_102
timestamp 1581320205
transform 1 0 8160 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_103
timestamp 1581320205
transform 1 0 6528 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_104
timestamp 1581320205
transform 1 0 4896 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_105
timestamp 1581320205
transform 1 0 3264 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_106
timestamp 1581320205
transform 1 0 1632 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_107
timestamp 1581320205
transform 1 0 0 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_108
timestamp 1581320205
transform 1 0 13056 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_109
timestamp 1581320205
transform 1 0 11424 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_110
timestamp 1581320205
transform 1 0 9792 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_111
timestamp 1581320205
transform 1 0 8160 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_112
timestamp 1581320205
transform 1 0 6528 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_113
timestamp 1581320205
transform 1 0 4896 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_114
timestamp 1581320205
transform 1 0 3264 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_115
timestamp 1581320205
transform 1 0 1632 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_116
timestamp 1581320205
transform 1 0 0 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_117
timestamp 1581320205
transform 1 0 13056 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_118
timestamp 1581320205
transform 1 0 11424 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_119
timestamp 1581320205
transform 1 0 9792 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_120
timestamp 1581320205
transform 1 0 8160 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_121
timestamp 1581320205
transform 1 0 6528 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_122
timestamp 1581320205
transform 1 0 4896 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_123
timestamp 1581320205
transform 1 0 3264 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_124
timestamp 1581320205
transform 1 0 1632 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_125
timestamp 1581320205
transform 1 0 0 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_126
timestamp 1581320205
transform 1 0 13056 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_127
timestamp 1581320205
transform 1 0 11424 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_128
timestamp 1581320205
transform 1 0 9792 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_129
timestamp 1581320205
transform 1 0 8160 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_130
timestamp 1581320205
transform 1 0 6528 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_131
timestamp 1581320205
transform 1 0 4896 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_132
timestamp 1581320205
transform 1 0 3264 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_133
timestamp 1581320205
transform 1 0 1632 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_134
timestamp 1581320205
transform 1 0 0 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_135
timestamp 1581320205
transform 1 0 13056 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_136
timestamp 1581320205
transform 1 0 11424 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_137
timestamp 1581320205
transform 1 0 9792 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_138
timestamp 1581320205
transform 1 0 8160 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_139
timestamp 1581320205
transform 1 0 6528 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_140
timestamp 1581320205
transform 1 0 4896 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_141
timestamp 1581320205
transform 1 0 3264 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_142
timestamp 1581320205
transform 1 0 1632 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_143
timestamp 1581320205
transform 1 0 0 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_144
timestamp 1581320205
transform 1 0 13056 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_145
timestamp 1581320205
transform 1 0 11424 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_146
timestamp 1581320205
transform 1 0 9792 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_147
timestamp 1581320205
transform 1 0 8160 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_148
timestamp 1581320205
transform 1 0 6528 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_149
timestamp 1581320205
transform 1 0 4896 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_150
timestamp 1581320205
transform 1 0 3264 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_151
timestamp 1581320205
transform 1 0 1632 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_152
timestamp 1581320205
transform 1 0 0 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_153
timestamp 1581320205
transform 1 0 13056 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_154
timestamp 1581320205
transform 1 0 11424 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_155
timestamp 1581320205
transform 1 0 9792 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_156
timestamp 1581320205
transform 1 0 8160 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_157
timestamp 1581320205
transform 1 0 6528 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_158
timestamp 1581320205
transform 1 0 4896 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_159
timestamp 1581320205
transform 1 0 3264 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_160
timestamp 1581320205
transform 1 0 1632 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_161
timestamp 1581320205
transform 1 0 0 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_162
timestamp 1581320205
transform 1 0 13056 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_163
timestamp 1581320205
transform 1 0 11424 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_164
timestamp 1581320205
transform 1 0 9792 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_165
timestamp 1581320205
transform 1 0 8160 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_166
timestamp 1581320205
transform 1 0 6528 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_167
timestamp 1581320205
transform 1 0 4896 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_168
timestamp 1581320205
transform 1 0 3264 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_169
timestamp 1581320205
transform 1 0 1632 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_170
timestamp 1581320205
transform 1 0 0 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_171
timestamp 1581320205
transform 1 0 13056 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_172
timestamp 1581320205
transform 1 0 11424 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_173
timestamp 1581320205
transform 1 0 9792 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_174
timestamp 1581320205
transform 1 0 8160 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_175
timestamp 1581320205
transform 1 0 6528 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_176
timestamp 1581320205
transform 1 0 4896 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_177
timestamp 1581320205
transform 1 0 3264 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_178
timestamp 1581320205
transform 1 0 1632 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_179
timestamp 1581320205
transform 1 0 0 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_180
timestamp 1581320205
transform 1 0 13056 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_181
timestamp 1581320205
transform 1 0 11424 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_182
timestamp 1581320205
transform 1 0 9792 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_183
timestamp 1581320205
transform 1 0 8160 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_184
timestamp 1581320205
transform 1 0 6528 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_185
timestamp 1581320205
transform 1 0 4896 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_186
timestamp 1581320205
transform 1 0 3264 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_187
timestamp 1581320205
transform 1 0 1632 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_188
timestamp 1581320205
transform 1 0 0 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_189
timestamp 1581320205
transform 1 0 13056 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_190
timestamp 1581320205
transform 1 0 11424 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_191
timestamp 1581320205
transform 1 0 9792 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_192
timestamp 1581320205
transform 1 0 8160 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_193
timestamp 1581320205
transform 1 0 6528 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_194
timestamp 1581320205
transform 1 0 4896 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_195
timestamp 1581320205
transform 1 0 3264 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_196
timestamp 1581320205
transform 1 0 1632 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_197
timestamp 1581320205
transform 1 0 0 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_198
timestamp 1581320205
transform 1 0 13056 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_199
timestamp 1581320205
transform 1 0 11424 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_200
timestamp 1581320205
transform 1 0 9792 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_201
timestamp 1581320205
transform 1 0 8160 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_202
timestamp 1581320205
transform 1 0 6528 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_203
timestamp 1581320205
transform 1 0 4896 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_204
timestamp 1581320205
transform 1 0 3264 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_205
timestamp 1581320205
transform 1 0 1632 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_206
timestamp 1581320205
transform 1 0 0 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_207
timestamp 1581320205
transform 1 0 13056 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_208
timestamp 1581320205
transform 1 0 11424 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_209
timestamp 1581320205
transform 1 0 9792 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_210
timestamp 1581320205
transform 1 0 8160 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_211
timestamp 1581320205
transform 1 0 6528 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_212
timestamp 1581320205
transform 1 0 4896 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_213
timestamp 1581320205
transform 1 0 3264 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_214
timestamp 1581320205
transform 1 0 1632 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_215
timestamp 1581320205
transform 1 0 0 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_216
timestamp 1581320205
transform 1 0 13056 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_217
timestamp 1581320205
transform 1 0 11424 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_218
timestamp 1581320205
transform 1 0 9792 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_219
timestamp 1581320205
transform 1 0 8160 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_220
timestamp 1581320205
transform 1 0 6528 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_221
timestamp 1581320205
transform 1 0 4896 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_222
timestamp 1581320205
transform 1 0 3264 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_223
timestamp 1581320205
transform 1 0 1632 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_224
timestamp 1581320205
transform 1 0 0 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_225
timestamp 1581320205
transform 1 0 13056 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_226
timestamp 1581320205
transform 1 0 11424 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_227
timestamp 1581320205
transform 1 0 9792 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_228
timestamp 1581320205
transform 1 0 8160 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_229
timestamp 1581320205
transform 1 0 6528 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_230
timestamp 1581320205
transform 1 0 4896 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_231
timestamp 1581320205
transform 1 0 3264 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_232
timestamp 1581320205
transform 1 0 1632 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_233
timestamp 1581320205
transform 1 0 0 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_234
timestamp 1581320205
transform 1 0 13056 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_235
timestamp 1581320205
transform 1 0 11424 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_236
timestamp 1581320205
transform 1 0 9792 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_237
timestamp 1581320205
transform 1 0 8160 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_238
timestamp 1581320205
transform 1 0 6528 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_239
timestamp 1581320205
transform 1 0 4896 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_240
timestamp 1581320205
transform 1 0 3264 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_241
timestamp 1581320205
transform 1 0 1632 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_242
timestamp 1581320205
transform 1 0 0 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_243
timestamp 1581320205
transform 1 0 13056 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_244
timestamp 1581320205
transform 1 0 11424 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_245
timestamp 1581320205
transform 1 0 9792 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_246
timestamp 1581320205
transform 1 0 8160 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_247
timestamp 1581320205
transform 1 0 6528 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_248
timestamp 1581320205
transform 1 0 4896 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_249
timestamp 1581320205
transform 1 0 3264 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_250
timestamp 1581320205
transform 1 0 1632 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_251
timestamp 1581320205
transform 1 0 0 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_252
timestamp 1581320205
transform 1 0 13056 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_253
timestamp 1581320205
transform 1 0 11424 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_254
timestamp 1581320205
transform 1 0 9792 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_255
timestamp 1581320205
transform 1 0 8160 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_256
timestamp 1581320205
transform 1 0 6528 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_257
timestamp 1581320205
transform 1 0 4896 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_258
timestamp 1581320205
transform 1 0 3264 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_259
timestamp 1581320205
transform 1 0 1632 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_260
timestamp 1581320205
transform 1 0 0 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_261
timestamp 1581320205
transform 1 0 13056 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_262
timestamp 1581320205
transform 1 0 11424 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_263
timestamp 1581320205
transform 1 0 9792 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_264
timestamp 1581320205
transform 1 0 8160 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_265
timestamp 1581320205
transform 1 0 6528 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_266
timestamp 1581320205
transform 1 0 4896 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_267
timestamp 1581320205
transform 1 0 3264 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_268
timestamp 1581320205
transform 1 0 1632 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_269
timestamp 1581320205
transform 1 0 0 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_270
timestamp 1581320205
transform 1 0 13056 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_271
timestamp 1581320205
transform 1 0 11424 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_272
timestamp 1581320205
transform 1 0 9792 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_273
timestamp 1581320205
transform 1 0 8160 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_274
timestamp 1581320205
transform 1 0 6528 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_275
timestamp 1581320205
transform 1 0 4896 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_276
timestamp 1581320205
transform 1 0 3264 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_277
timestamp 1581320205
transform 1 0 1632 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_278
timestamp 1581320205
transform 1 0 0 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_279
timestamp 1581320205
transform 1 0 13056 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_280
timestamp 1581320205
transform 1 0 11424 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_281
timestamp 1581320205
transform 1 0 9792 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_282
timestamp 1581320205
transform 1 0 8160 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_283
timestamp 1581320205
transform 1 0 6528 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_284
timestamp 1581320205
transform 1 0 4896 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_285
timestamp 1581320205
transform 1 0 3264 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_286
timestamp 1581320205
transform 1 0 1632 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_287
timestamp 1581320205
transform 1 0 0 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_288
timestamp 1581320205
transform 1 0 13056 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_289
timestamp 1581320205
transform 1 0 11424 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_290
timestamp 1581320205
transform 1 0 9792 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_291
timestamp 1581320205
transform 1 0 8160 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_292
timestamp 1581320205
transform 1 0 6528 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_293
timestamp 1581320205
transform 1 0 4896 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_294
timestamp 1581320205
transform 1 0 3264 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_295
timestamp 1581320205
transform 1 0 1632 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_296
timestamp 1581320205
transform 1 0 0 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_precharge_array  sky130_rom_krom_rom_precharge_array_0
timestamp 1581320205
transform 1 0 0 0 1 128
box 0 -212 13164 408
<< labels >>
rlabel metal2 s 61 368 89 396 4 precharge
port 3 nsew
rlabel metal2 s 19 1013 47 1041 4 wl_0_0
port 5 nsew
rlabel metal2 s 19 1217 47 1245 4 wl_0_1
port 7 nsew
rlabel metal2 s 19 1421 47 1449 4 wl_0_2
port 9 nsew
rlabel metal2 s 19 1625 47 1653 4 wl_0_3
port 11 nsew
rlabel metal2 s 19 1829 47 1857 4 wl_0_4
port 13 nsew
rlabel metal2 s 19 2033 47 2061 4 wl_0_5
port 15 nsew
rlabel metal2 s 19 2237 47 2265 4 wl_0_6
port 17 nsew
rlabel metal2 s 19 2441 47 2469 4 wl_0_7
port 19 nsew
rlabel metal2 s 19 2749 47 2777 4 wl_0_8
port 21 nsew
rlabel metal2 s 19 2953 47 2981 4 wl_0_9
port 23 nsew
rlabel metal2 s 19 3157 47 3185 4 wl_0_10
port 25 nsew
rlabel metal2 s 19 3361 47 3389 4 wl_0_11
port 27 nsew
rlabel metal2 s 19 3565 47 3593 4 wl_0_12
port 29 nsew
rlabel metal2 s 19 3769 47 3797 4 wl_0_13
port 31 nsew
rlabel metal2 s 19 3973 47 4001 4 wl_0_14
port 33 nsew
rlabel metal2 s 19 4177 47 4205 4 wl_0_15
port 35 nsew
rlabel metal2 s 19 4485 47 4513 4 wl_0_16
port 37 nsew
rlabel metal2 s 19 4689 47 4717 4 wl_0_17
port 39 nsew
rlabel metal2 s 19 4893 47 4921 4 wl_0_18
port 41 nsew
rlabel metal2 s 19 5097 47 5125 4 wl_0_19
port 43 nsew
rlabel metal2 s 19 5301 47 5329 4 wl_0_20
port 45 nsew
rlabel metal2 s 19 5505 47 5533 4 wl_0_21
port 47 nsew
rlabel metal2 s 19 5709 47 5737 4 wl_0_22
port 49 nsew
rlabel metal2 s 19 5913 47 5941 4 wl_0_23
port 51 nsew
rlabel metal2 s 19 6221 47 6249 4 wl_0_24
port 53 nsew
rlabel metal2 s 19 6425 47 6453 4 wl_0_25
port 55 nsew
rlabel metal2 s 19 6629 47 6657 4 wl_0_26
port 57 nsew
rlabel metal2 s 19 6833 47 6861 4 wl_0_27
port 59 nsew
rlabel metal2 s 19 7037 47 7065 4 wl_0_28
port 61 nsew
rlabel metal2 s 19 7241 47 7269 4 wl_0_29
port 63 nsew
rlabel metal2 s 19 7445 47 7473 4 wl_0_30
port 65 nsew
rlabel metal2 s 19 7649 47 7677 4 wl_0_31
port 67 nsew
rlabel metal1 s 128 -14 156 14 4 bl_0_0
port 69 nsew
rlabel metal1 s 332 -14 360 14 4 bl_0_1
port 71 nsew
rlabel metal1 s 536 -14 564 14 4 bl_0_2
port 73 nsew
rlabel metal1 s 740 -14 768 14 4 bl_0_3
port 75 nsew
rlabel metal1 s 944 -14 972 14 4 bl_0_4
port 77 nsew
rlabel metal1 s 1148 -14 1176 14 4 bl_0_5
port 79 nsew
rlabel metal1 s 1352 -14 1380 14 4 bl_0_6
port 81 nsew
rlabel metal1 s 1556 -14 1584 14 4 bl_0_7
port 83 nsew
rlabel metal1 s 1760 -14 1788 14 4 bl_0_8
port 85 nsew
rlabel metal1 s 1964 -14 1992 14 4 bl_0_9
port 87 nsew
rlabel metal1 s 2168 -14 2196 14 4 bl_0_10
port 89 nsew
rlabel metal1 s 2372 -14 2400 14 4 bl_0_11
port 91 nsew
rlabel metal1 s 2576 -14 2604 14 4 bl_0_12
port 93 nsew
rlabel metal1 s 2780 -14 2808 14 4 bl_0_13
port 95 nsew
rlabel metal1 s 2984 -14 3012 14 4 bl_0_14
port 97 nsew
rlabel metal1 s 3188 -14 3216 14 4 bl_0_15
port 99 nsew
rlabel metal1 s 3392 -14 3420 14 4 bl_0_16
port 101 nsew
rlabel metal1 s 3596 -14 3624 14 4 bl_0_17
port 103 nsew
rlabel metal1 s 3800 -14 3828 14 4 bl_0_18
port 105 nsew
rlabel metal1 s 4004 -14 4032 14 4 bl_0_19
port 107 nsew
rlabel metal1 s 4208 -14 4236 14 4 bl_0_20
port 109 nsew
rlabel metal1 s 4412 -14 4440 14 4 bl_0_21
port 111 nsew
rlabel metal1 s 4616 -14 4644 14 4 bl_0_22
port 113 nsew
rlabel metal1 s 4820 -14 4848 14 4 bl_0_23
port 115 nsew
rlabel metal1 s 5024 -14 5052 14 4 bl_0_24
port 117 nsew
rlabel metal1 s 5228 -14 5256 14 4 bl_0_25
port 119 nsew
rlabel metal1 s 5432 -14 5460 14 4 bl_0_26
port 121 nsew
rlabel metal1 s 5636 -14 5664 14 4 bl_0_27
port 123 nsew
rlabel metal1 s 5840 -14 5868 14 4 bl_0_28
port 125 nsew
rlabel metal1 s 6044 -14 6072 14 4 bl_0_29
port 127 nsew
rlabel metal1 s 6248 -14 6276 14 4 bl_0_30
port 129 nsew
rlabel metal1 s 6452 -14 6480 14 4 bl_0_31
port 131 nsew
rlabel metal1 s 6656 -14 6684 14 4 bl_0_32
port 133 nsew
rlabel metal1 s 6860 -14 6888 14 4 bl_0_33
port 135 nsew
rlabel metal1 s 7064 -14 7092 14 4 bl_0_34
port 137 nsew
rlabel metal1 s 7268 -14 7296 14 4 bl_0_35
port 139 nsew
rlabel metal1 s 7472 -14 7500 14 4 bl_0_36
port 141 nsew
rlabel metal1 s 7676 -14 7704 14 4 bl_0_37
port 143 nsew
rlabel metal1 s 7880 -14 7908 14 4 bl_0_38
port 145 nsew
rlabel metal1 s 8084 -14 8112 14 4 bl_0_39
port 147 nsew
rlabel metal1 s 8288 -14 8316 14 4 bl_0_40
port 149 nsew
rlabel metal1 s 8492 -14 8520 14 4 bl_0_41
port 151 nsew
rlabel metal1 s 8696 -14 8724 14 4 bl_0_42
port 153 nsew
rlabel metal1 s 8900 -14 8928 14 4 bl_0_43
port 155 nsew
rlabel metal1 s 9104 -14 9132 14 4 bl_0_44
port 157 nsew
rlabel metal1 s 9308 -14 9336 14 4 bl_0_45
port 159 nsew
rlabel metal1 s 9512 -14 9540 14 4 bl_0_46
port 161 nsew
rlabel metal1 s 9716 -14 9744 14 4 bl_0_47
port 163 nsew
rlabel metal1 s 9920 -14 9948 14 4 bl_0_48
port 165 nsew
rlabel metal1 s 10124 -14 10152 14 4 bl_0_49
port 167 nsew
rlabel metal1 s 10328 -14 10356 14 4 bl_0_50
port 169 nsew
rlabel metal1 s 10532 -14 10560 14 4 bl_0_51
port 171 nsew
rlabel metal1 s 10736 -14 10764 14 4 bl_0_52
port 173 nsew
rlabel metal1 s 10940 -14 10968 14 4 bl_0_53
port 175 nsew
rlabel metal1 s 11144 -14 11172 14 4 bl_0_54
port 177 nsew
rlabel metal1 s 11348 -14 11376 14 4 bl_0_55
port 179 nsew
rlabel metal1 s 11552 -14 11580 14 4 bl_0_56
port 181 nsew
rlabel metal1 s 11756 -14 11784 14 4 bl_0_57
port 183 nsew
rlabel metal1 s 11960 -14 11988 14 4 bl_0_58
port 185 nsew
rlabel metal1 s 12164 -14 12192 14 4 bl_0_59
port 187 nsew
rlabel metal1 s 12368 -14 12396 14 4 bl_0_60
port 189 nsew
rlabel metal1 s 12572 -14 12600 14 4 bl_0_61
port 191 nsew
rlabel metal1 s 12776 -14 12804 14 4 bl_0_62
port 193 nsew
rlabel metal1 s 12980 -14 13008 14 4 bl_0_63
port 195 nsew
rlabel metal1 s 13277 368 13305 396 4 precharge_r
port 197 nsew
rlabel metal2 s 230 2595 13124 2623 4 gnd
port 199 nsew
rlabel metal2 s 230 4331 13124 4359 4 gnd
port 199 nsew
rlabel metal2 s 230 6067 13124 6095 4 gnd
port 199 nsew
rlabel metal1 s 12994 7980 13022 8008 4 gnd
port 199 nsew
rlabel metal1 s 114 7980 142 8008 4 gnd
port 199 nsew
rlabel metal2 s 230 859 13124 887 4 gnd
port 199 nsew
rlabel metal2 s 12 -32 40 32 4 vdd
port 201 nsew
<< properties >>
string FIXED_BBOX 0 0 13305 974
<< end >>
