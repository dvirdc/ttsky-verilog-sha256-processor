magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1260 -878 11103 3301
<< poly >>
rect 87 641 117 1252
rect 291 845 321 1252
rect 495 1049 525 1252
rect 586 1051 652 1067
rect 586 1049 602 1051
rect 495 1019 602 1049
rect 586 1017 602 1019
rect 636 1017 652 1051
rect 586 1001 652 1017
rect 382 847 448 863
rect 382 845 398 847
rect 291 815 398 845
rect 382 813 398 815
rect 432 813 448 847
rect 382 797 448 813
rect 178 643 244 659
rect 178 641 194 643
rect 87 611 194 641
rect 178 609 194 611
rect 228 609 244 643
rect 699 641 729 1252
rect 903 845 933 1252
rect 1107 1049 1137 1252
rect 1198 1051 1264 1067
rect 1198 1049 1214 1051
rect 1107 1019 1214 1049
rect 1198 1017 1214 1019
rect 1248 1017 1264 1051
rect 1198 1001 1264 1017
rect 994 847 1060 863
rect 994 845 1010 847
rect 903 815 1010 845
rect 994 813 1010 815
rect 1044 813 1060 847
rect 994 797 1060 813
rect 790 643 856 659
rect 790 641 806 643
rect 699 611 806 641
rect 178 593 244 609
rect 790 609 806 611
rect 840 609 856 643
rect 1311 641 1341 1252
rect 1515 845 1545 1252
rect 1719 1049 1749 1252
rect 1810 1051 1876 1067
rect 1810 1049 1826 1051
rect 1719 1019 1826 1049
rect 1810 1017 1826 1019
rect 1860 1017 1876 1051
rect 1810 1001 1876 1017
rect 1606 847 1672 863
rect 1606 845 1622 847
rect 1515 815 1622 845
rect 1606 813 1622 815
rect 1656 813 1672 847
rect 1606 797 1672 813
rect 1402 643 1468 659
rect 1402 641 1418 643
rect 1311 611 1418 641
rect 790 593 856 609
rect 1402 609 1418 611
rect 1452 609 1468 643
rect 1923 641 1953 1252
rect 2127 845 2157 1252
rect 2331 1049 2361 1252
rect 2422 1051 2488 1067
rect 2422 1049 2438 1051
rect 2331 1019 2438 1049
rect 2422 1017 2438 1019
rect 2472 1017 2488 1051
rect 2422 1001 2488 1017
rect 2218 847 2284 863
rect 2218 845 2234 847
rect 2127 815 2234 845
rect 2218 813 2234 815
rect 2268 813 2284 847
rect 2218 797 2284 813
rect 2014 643 2080 659
rect 2014 641 2030 643
rect 1923 611 2030 641
rect 1402 593 1468 609
rect 2014 609 2030 611
rect 2064 609 2080 643
rect 2535 641 2565 1252
rect 2739 845 2769 1252
rect 2943 1049 2973 1252
rect 3034 1051 3100 1067
rect 3034 1049 3050 1051
rect 2943 1019 3050 1049
rect 3034 1017 3050 1019
rect 3084 1017 3100 1051
rect 3034 1001 3100 1017
rect 2830 847 2896 863
rect 2830 845 2846 847
rect 2739 815 2846 845
rect 2830 813 2846 815
rect 2880 813 2896 847
rect 2830 797 2896 813
rect 2626 643 2692 659
rect 2626 641 2642 643
rect 2535 611 2642 641
rect 2014 593 2080 609
rect 2626 609 2642 611
rect 2676 609 2692 643
rect 3147 641 3177 1252
rect 3351 845 3381 1252
rect 3555 1049 3585 1252
rect 3646 1051 3712 1067
rect 3646 1049 3662 1051
rect 3555 1019 3662 1049
rect 3646 1017 3662 1019
rect 3696 1017 3712 1051
rect 3646 1001 3712 1017
rect 3442 847 3508 863
rect 3442 845 3458 847
rect 3351 815 3458 845
rect 3442 813 3458 815
rect 3492 813 3508 847
rect 3442 797 3508 813
rect 3238 643 3304 659
rect 3238 641 3254 643
rect 3147 611 3254 641
rect 2626 593 2692 609
rect 3238 609 3254 611
rect 3288 609 3304 643
rect 3759 641 3789 1252
rect 3963 845 3993 1252
rect 4167 1049 4197 1252
rect 4258 1051 4324 1067
rect 4258 1049 4274 1051
rect 4167 1019 4274 1049
rect 4258 1017 4274 1019
rect 4308 1017 4324 1051
rect 4258 1001 4324 1017
rect 4054 847 4120 863
rect 4054 845 4070 847
rect 3963 815 4070 845
rect 4054 813 4070 815
rect 4104 813 4120 847
rect 4054 797 4120 813
rect 3850 643 3916 659
rect 3850 641 3866 643
rect 3759 611 3866 641
rect 3238 593 3304 609
rect 3850 609 3866 611
rect 3900 609 3916 643
rect 4371 641 4401 1252
rect 4575 845 4605 1252
rect 4779 1049 4809 1252
rect 4870 1051 4936 1067
rect 4870 1049 4886 1051
rect 4779 1019 4886 1049
rect 4870 1017 4886 1019
rect 4920 1017 4936 1051
rect 4870 1001 4936 1017
rect 4666 847 4732 863
rect 4666 845 4682 847
rect 4575 815 4682 845
rect 4666 813 4682 815
rect 4716 813 4732 847
rect 4666 797 4732 813
rect 4462 643 4528 659
rect 4462 641 4478 643
rect 4371 611 4478 641
rect 3850 593 3916 609
rect 4462 609 4478 611
rect 4512 609 4528 643
rect 4983 641 5013 1252
rect 5187 845 5217 1252
rect 5391 1049 5421 1252
rect 5482 1051 5548 1067
rect 5482 1049 5498 1051
rect 5391 1019 5498 1049
rect 5482 1017 5498 1019
rect 5532 1017 5548 1051
rect 5482 1001 5548 1017
rect 5278 847 5344 863
rect 5278 845 5294 847
rect 5187 815 5294 845
rect 5278 813 5294 815
rect 5328 813 5344 847
rect 5278 797 5344 813
rect 5074 643 5140 659
rect 5074 641 5090 643
rect 4983 611 5090 641
rect 4462 593 4528 609
rect 5074 609 5090 611
rect 5124 609 5140 643
rect 5595 641 5625 1252
rect 5799 845 5829 1252
rect 6003 1049 6033 1252
rect 6094 1051 6160 1067
rect 6094 1049 6110 1051
rect 6003 1019 6110 1049
rect 6094 1017 6110 1019
rect 6144 1017 6160 1051
rect 6094 1001 6160 1017
rect 5890 847 5956 863
rect 5890 845 5906 847
rect 5799 815 5906 845
rect 5890 813 5906 815
rect 5940 813 5956 847
rect 5890 797 5956 813
rect 5686 643 5752 659
rect 5686 641 5702 643
rect 5595 611 5702 641
rect 5074 593 5140 609
rect 5686 609 5702 611
rect 5736 609 5752 643
rect 6207 641 6237 1252
rect 6411 845 6441 1252
rect 6615 1049 6645 1252
rect 6706 1051 6772 1067
rect 6706 1049 6722 1051
rect 6615 1019 6722 1049
rect 6706 1017 6722 1019
rect 6756 1017 6772 1051
rect 6706 1001 6772 1017
rect 6502 847 6568 863
rect 6502 845 6518 847
rect 6411 815 6518 845
rect 6502 813 6518 815
rect 6552 813 6568 847
rect 6502 797 6568 813
rect 6298 643 6364 659
rect 6298 641 6314 643
rect 6207 611 6314 641
rect 5686 593 5752 609
rect 6298 609 6314 611
rect 6348 609 6364 643
rect 6819 641 6849 1252
rect 7023 845 7053 1252
rect 7227 1049 7257 1252
rect 7318 1051 7384 1067
rect 7318 1049 7334 1051
rect 7227 1019 7334 1049
rect 7318 1017 7334 1019
rect 7368 1017 7384 1051
rect 7318 1001 7384 1017
rect 7114 847 7180 863
rect 7114 845 7130 847
rect 7023 815 7130 845
rect 7114 813 7130 815
rect 7164 813 7180 847
rect 7114 797 7180 813
rect 6910 643 6976 659
rect 6910 641 6926 643
rect 6819 611 6926 641
rect 6298 593 6364 609
rect 6910 609 6926 611
rect 6960 609 6976 643
rect 7431 641 7461 1252
rect 7635 845 7665 1252
rect 7839 1049 7869 1252
rect 7930 1051 7996 1067
rect 7930 1049 7946 1051
rect 7839 1019 7946 1049
rect 7930 1017 7946 1019
rect 7980 1017 7996 1051
rect 7930 1001 7996 1017
rect 7726 847 7792 863
rect 7726 845 7742 847
rect 7635 815 7742 845
rect 7726 813 7742 815
rect 7776 813 7792 847
rect 7726 797 7792 813
rect 7522 643 7588 659
rect 7522 641 7538 643
rect 7431 611 7538 641
rect 6910 593 6976 609
rect 7522 609 7538 611
rect 7572 609 7588 643
rect 8043 641 8073 1252
rect 8247 845 8277 1252
rect 8451 1049 8481 1252
rect 8542 1051 8608 1067
rect 8542 1049 8558 1051
rect 8451 1019 8558 1049
rect 8542 1017 8558 1019
rect 8592 1017 8608 1051
rect 8542 1001 8608 1017
rect 8338 847 8404 863
rect 8338 845 8354 847
rect 8247 815 8354 845
rect 8338 813 8354 815
rect 8388 813 8404 847
rect 8338 797 8404 813
rect 8134 643 8200 659
rect 8134 641 8150 643
rect 8043 611 8150 641
rect 7522 593 7588 609
rect 8134 609 8150 611
rect 8184 609 8200 643
rect 8655 641 8685 1252
rect 8859 845 8889 1252
rect 9063 1049 9093 1252
rect 9154 1051 9220 1067
rect 9154 1049 9170 1051
rect 9063 1019 9170 1049
rect 9154 1017 9170 1019
rect 9204 1017 9220 1051
rect 9154 1001 9220 1017
rect 8950 847 9016 863
rect 8950 845 8966 847
rect 8859 815 8966 845
rect 8950 813 8966 815
rect 9000 813 9016 847
rect 8950 797 9016 813
rect 8746 643 8812 659
rect 8746 641 8762 643
rect 8655 611 8762 641
rect 8134 593 8200 609
rect 8746 609 8762 611
rect 8796 609 8812 643
rect 9267 641 9297 1252
rect 9471 845 9501 1252
rect 9675 1049 9705 1252
rect 9766 1051 9832 1067
rect 9766 1049 9782 1051
rect 9675 1019 9782 1049
rect 9766 1017 9782 1019
rect 9816 1017 9832 1051
rect 9766 1001 9832 1017
rect 9562 847 9628 863
rect 9562 845 9578 847
rect 9471 815 9578 845
rect 9562 813 9578 815
rect 9612 813 9628 847
rect 9562 797 9628 813
rect 9358 643 9424 659
rect 9358 641 9374 643
rect 9267 611 9374 641
rect 8746 593 8812 609
rect 9358 609 9374 611
rect 9408 609 9424 643
rect 9358 593 9424 609
<< polycont >>
rect 602 1017 636 1051
rect 398 813 432 847
rect 194 609 228 643
rect 1214 1017 1248 1051
rect 1010 813 1044 847
rect 806 609 840 643
rect 1826 1017 1860 1051
rect 1622 813 1656 847
rect 1418 609 1452 643
rect 2438 1017 2472 1051
rect 2234 813 2268 847
rect 2030 609 2064 643
rect 3050 1017 3084 1051
rect 2846 813 2880 847
rect 2642 609 2676 643
rect 3662 1017 3696 1051
rect 3458 813 3492 847
rect 3254 609 3288 643
rect 4274 1017 4308 1051
rect 4070 813 4104 847
rect 3866 609 3900 643
rect 4886 1017 4920 1051
rect 4682 813 4716 847
rect 4478 609 4512 643
rect 5498 1017 5532 1051
rect 5294 813 5328 847
rect 5090 609 5124 643
rect 6110 1017 6144 1051
rect 5906 813 5940 847
rect 5702 609 5736 643
rect 6722 1017 6756 1051
rect 6518 813 6552 847
rect 6314 609 6348 643
rect 7334 1017 7368 1051
rect 7130 813 7164 847
rect 6926 609 6960 643
rect 7946 1017 7980 1051
rect 7742 813 7776 847
rect 7538 609 7572 643
rect 8558 1017 8592 1051
rect 8354 813 8388 847
rect 8150 609 8184 643
rect 9170 1017 9204 1051
rect 8966 813 9000 847
rect 8762 609 8796 643
rect 9782 1017 9816 1051
rect 9578 813 9612 847
rect 9374 609 9408 643
<< locali >>
rect 586 1017 602 1051
rect 636 1017 652 1051
rect 1198 1017 1214 1051
rect 1248 1017 1264 1051
rect 1810 1017 1826 1051
rect 1860 1017 1876 1051
rect 2422 1017 2438 1051
rect 2472 1017 2488 1051
rect 3034 1017 3050 1051
rect 3084 1017 3100 1051
rect 3646 1017 3662 1051
rect 3696 1017 3712 1051
rect 4258 1017 4274 1051
rect 4308 1017 4324 1051
rect 4870 1017 4886 1051
rect 4920 1017 4936 1051
rect 5482 1017 5498 1051
rect 5532 1017 5548 1051
rect 6094 1017 6110 1051
rect 6144 1017 6160 1051
rect 6706 1017 6722 1051
rect 6756 1017 6772 1051
rect 7318 1017 7334 1051
rect 7368 1017 7384 1051
rect 7930 1017 7946 1051
rect 7980 1017 7996 1051
rect 8542 1017 8558 1051
rect 8592 1017 8608 1051
rect 9154 1017 9170 1051
rect 9204 1017 9220 1051
rect 9766 1017 9782 1051
rect 9816 1017 9832 1051
rect 382 813 398 847
rect 432 813 448 847
rect 994 813 1010 847
rect 1044 813 1060 847
rect 1606 813 1622 847
rect 1656 813 1672 847
rect 2218 813 2234 847
rect 2268 813 2284 847
rect 2830 813 2846 847
rect 2880 813 2896 847
rect 3442 813 3458 847
rect 3492 813 3508 847
rect 4054 813 4070 847
rect 4104 813 4120 847
rect 4666 813 4682 847
rect 4716 813 4732 847
rect 5278 813 5294 847
rect 5328 813 5344 847
rect 5890 813 5906 847
rect 5940 813 5956 847
rect 6502 813 6518 847
rect 6552 813 6568 847
rect 7114 813 7130 847
rect 7164 813 7180 847
rect 7726 813 7742 847
rect 7776 813 7792 847
rect 8338 813 8354 847
rect 8388 813 8404 847
rect 8950 813 8966 847
rect 9000 813 9016 847
rect 9562 813 9578 847
rect 9612 813 9628 847
rect 178 609 194 643
rect 228 609 244 643
rect 790 609 806 643
rect 840 609 856 643
rect 1402 609 1418 643
rect 1452 609 1468 643
rect 2014 609 2030 643
rect 2064 609 2080 643
rect 2626 609 2642 643
rect 2676 609 2692 643
rect 3238 609 3254 643
rect 3288 609 3304 643
rect 3850 609 3866 643
rect 3900 609 3916 643
rect 4462 609 4478 643
rect 4512 609 4528 643
rect 5074 609 5090 643
rect 5124 609 5140 643
rect 5686 609 5702 643
rect 5736 609 5752 643
rect 6298 609 6314 643
rect 6348 609 6364 643
rect 6910 609 6926 643
rect 6960 609 6976 643
rect 7522 609 7538 643
rect 7572 609 7588 643
rect 8134 609 8150 643
rect 8184 609 8200 643
rect 8746 609 8762 643
rect 8796 609 8812 643
rect 9358 609 9374 643
rect 9408 609 9424 643
<< viali >>
rect 602 1017 636 1051
rect 1214 1017 1248 1051
rect 1826 1017 1860 1051
rect 2438 1017 2472 1051
rect 3050 1017 3084 1051
rect 3662 1017 3696 1051
rect 4274 1017 4308 1051
rect 4886 1017 4920 1051
rect 5498 1017 5532 1051
rect 6110 1017 6144 1051
rect 6722 1017 6756 1051
rect 7334 1017 7368 1051
rect 7946 1017 7980 1051
rect 8558 1017 8592 1051
rect 9170 1017 9204 1051
rect 9782 1017 9816 1051
rect 398 813 432 847
rect 1010 813 1044 847
rect 1622 813 1656 847
rect 2234 813 2268 847
rect 2846 813 2880 847
rect 3458 813 3492 847
rect 4070 813 4104 847
rect 4682 813 4716 847
rect 5294 813 5328 847
rect 5906 813 5940 847
rect 6518 813 6552 847
rect 7130 813 7164 847
rect 7742 813 7776 847
rect 8354 813 8388 847
rect 8966 813 9000 847
rect 9578 813 9612 847
rect 194 609 228 643
rect 806 609 840 643
rect 1418 609 1452 643
rect 2030 609 2064 643
rect 2642 609 2676 643
rect 3254 609 3288 643
rect 3866 609 3900 643
rect 4478 609 4512 643
rect 5090 609 5124 643
rect 5702 609 5736 643
rect 6314 609 6348 643
rect 6926 609 6960 643
rect 7538 609 7572 643
rect 8150 609 8184 643
rect 8762 609 8796 643
rect 9374 609 9408 643
<< metal1 >>
rect 80 1854 108 2006
rect 172 1948 178 2000
rect 230 1948 236 2000
rect 284 1854 312 2006
rect 376 1948 382 2000
rect 434 1948 440 2000
rect 488 1854 516 2006
rect 580 1948 586 2000
rect 638 1948 644 2000
rect 692 1854 720 2006
rect 784 1948 790 2000
rect 842 1948 848 2000
rect 896 1854 924 2006
rect 988 1948 994 2000
rect 1046 1948 1052 2000
rect 1100 1854 1128 2006
rect 1192 1948 1198 2000
rect 1250 1948 1256 2000
rect 1304 1854 1332 2006
rect 1396 1948 1402 2000
rect 1454 1948 1460 2000
rect 1508 1854 1536 2006
rect 1600 1948 1606 2000
rect 1658 1948 1664 2000
rect 1712 1854 1740 2006
rect 1804 1948 1810 2000
rect 1862 1948 1868 2000
rect 1916 1854 1944 2006
rect 2008 1948 2014 2000
rect 2066 1948 2072 2000
rect 2120 1854 2148 2006
rect 2212 1948 2218 2000
rect 2270 1948 2276 2000
rect 2324 1854 2352 2006
rect 2416 1948 2422 2000
rect 2474 1948 2480 2000
rect 2528 1854 2556 2006
rect 2620 1948 2626 2000
rect 2678 1948 2684 2000
rect 2732 1854 2760 2006
rect 2824 1948 2830 2000
rect 2882 1948 2888 2000
rect 2936 1854 2964 2006
rect 3028 1948 3034 2000
rect 3086 1948 3092 2000
rect 3140 1854 3168 2006
rect 3232 1948 3238 2000
rect 3290 1948 3296 2000
rect 3344 1854 3372 2006
rect 3436 1948 3442 2000
rect 3494 1948 3500 2000
rect 3548 1854 3576 2006
rect 3640 1948 3646 2000
rect 3698 1948 3704 2000
rect 3752 1854 3780 2006
rect 3844 1948 3850 2000
rect 3902 1948 3908 2000
rect 3956 1854 3984 2006
rect 4048 1948 4054 2000
rect 4106 1948 4112 2000
rect 4160 1854 4188 2006
rect 4252 1948 4258 2000
rect 4310 1948 4316 2000
rect 4364 1854 4392 2006
rect 4456 1948 4462 2000
rect 4514 1948 4520 2000
rect 4568 1854 4596 2006
rect 4660 1948 4666 2000
rect 4718 1948 4724 2000
rect 4772 1854 4800 2006
rect 4864 1948 4870 2000
rect 4922 1948 4928 2000
rect 4976 1854 5004 2006
rect 5068 1948 5074 2000
rect 5126 1948 5132 2000
rect 5180 1854 5208 2006
rect 5272 1948 5278 2000
rect 5330 1948 5336 2000
rect 5384 1854 5412 2006
rect 5476 1948 5482 2000
rect 5534 1948 5540 2000
rect 5588 1854 5616 2006
rect 5680 1948 5686 2000
rect 5738 1948 5744 2000
rect 5792 1854 5820 2006
rect 5884 1948 5890 2000
rect 5942 1948 5948 2000
rect 5996 1854 6024 2006
rect 6088 1948 6094 2000
rect 6146 1948 6152 2000
rect 6200 1854 6228 2006
rect 6292 1948 6298 2000
rect 6350 1948 6356 2000
rect 6404 1854 6432 2006
rect 6496 1948 6502 2000
rect 6554 1948 6560 2000
rect 6608 1854 6636 2006
rect 6700 1948 6706 2000
rect 6758 1948 6764 2000
rect 6812 1854 6840 2006
rect 6904 1948 6910 2000
rect 6962 1948 6968 2000
rect 7016 1854 7044 2006
rect 7108 1948 7114 2000
rect 7166 1948 7172 2000
rect 7220 1854 7248 2006
rect 7312 1948 7318 2000
rect 7370 1948 7376 2000
rect 7424 1854 7452 2006
rect 7516 1948 7522 2000
rect 7574 1948 7580 2000
rect 7628 1854 7656 2006
rect 7720 1948 7726 2000
rect 7778 1948 7784 2000
rect 7832 1854 7860 2006
rect 7924 1948 7930 2000
rect 7982 1948 7988 2000
rect 8036 1854 8064 2006
rect 8128 1948 8134 2000
rect 8186 1948 8192 2000
rect 8240 1854 8268 2006
rect 8332 1948 8338 2000
rect 8390 1948 8396 2000
rect 8444 1854 8472 2006
rect 8536 1948 8542 2000
rect 8594 1948 8600 2000
rect 8648 1854 8676 2006
rect 8740 1948 8746 2000
rect 8798 1948 8804 2000
rect 8852 1854 8880 2006
rect 8944 1948 8950 2000
rect 9002 1948 9008 2000
rect 9056 1854 9084 2006
rect 9148 1948 9154 2000
rect 9206 1948 9212 2000
rect 9260 1854 9288 2006
rect 9352 1948 9358 2000
rect 9410 1948 9416 2000
rect 9464 1854 9492 2006
rect 9556 1948 9562 2000
rect 9614 1948 9620 2000
rect 9668 1854 9696 2006
rect 9760 1948 9766 2000
rect 9818 1948 9824 2000
rect 80 434 108 1224
rect 179 600 185 652
rect 237 600 243 652
rect 284 434 312 1224
rect 383 804 389 856
rect 441 804 447 856
rect 488 434 516 1224
rect 587 1008 593 1060
rect 645 1008 651 1060
rect 692 434 720 1224
rect 791 600 797 652
rect 849 600 855 652
rect 896 434 924 1224
rect 995 804 1001 856
rect 1053 804 1059 856
rect 1100 434 1128 1224
rect 1199 1008 1205 1060
rect 1257 1008 1263 1060
rect 1304 434 1332 1224
rect 1403 600 1409 652
rect 1461 600 1467 652
rect 1508 434 1536 1224
rect 1607 804 1613 856
rect 1665 804 1671 856
rect 1712 434 1740 1224
rect 1811 1008 1817 1060
rect 1869 1008 1875 1060
rect 1916 434 1944 1224
rect 2015 600 2021 652
rect 2073 600 2079 652
rect 2120 434 2148 1224
rect 2219 804 2225 856
rect 2277 804 2283 856
rect 2324 434 2352 1224
rect 2423 1008 2429 1060
rect 2481 1008 2487 1060
rect 2528 434 2556 1224
rect 2627 600 2633 652
rect 2685 600 2691 652
rect 2732 434 2760 1224
rect 2831 804 2837 856
rect 2889 804 2895 856
rect 2936 434 2964 1224
rect 3035 1008 3041 1060
rect 3093 1008 3099 1060
rect 3140 434 3168 1224
rect 3239 600 3245 652
rect 3297 600 3303 652
rect 3344 434 3372 1224
rect 3443 804 3449 856
rect 3501 804 3507 856
rect 3548 434 3576 1224
rect 3647 1008 3653 1060
rect 3705 1008 3711 1060
rect 3752 434 3780 1224
rect 3851 600 3857 652
rect 3909 600 3915 652
rect 3956 434 3984 1224
rect 4055 804 4061 856
rect 4113 804 4119 856
rect 4160 434 4188 1224
rect 4259 1008 4265 1060
rect 4317 1008 4323 1060
rect 4364 434 4392 1224
rect 4463 600 4469 652
rect 4521 600 4527 652
rect 4568 434 4596 1224
rect 4667 804 4673 856
rect 4725 804 4731 856
rect 4772 434 4800 1224
rect 4871 1008 4877 1060
rect 4929 1008 4935 1060
rect 4976 434 5004 1224
rect 5075 600 5081 652
rect 5133 600 5139 652
rect 5180 434 5208 1224
rect 5279 804 5285 856
rect 5337 804 5343 856
rect 5384 434 5412 1224
rect 5483 1008 5489 1060
rect 5541 1008 5547 1060
rect 5588 434 5616 1224
rect 5687 600 5693 652
rect 5745 600 5751 652
rect 5792 434 5820 1224
rect 5891 804 5897 856
rect 5949 804 5955 856
rect 5996 434 6024 1224
rect 6095 1008 6101 1060
rect 6153 1008 6159 1060
rect 6200 434 6228 1224
rect 6299 600 6305 652
rect 6357 600 6363 652
rect 6404 434 6432 1224
rect 6503 804 6509 856
rect 6561 804 6567 856
rect 6608 434 6636 1224
rect 6707 1008 6713 1060
rect 6765 1008 6771 1060
rect 6812 434 6840 1224
rect 6911 600 6917 652
rect 6969 600 6975 652
rect 7016 434 7044 1224
rect 7115 804 7121 856
rect 7173 804 7179 856
rect 7220 434 7248 1224
rect 7319 1008 7325 1060
rect 7377 1008 7383 1060
rect 7424 434 7452 1224
rect 7523 600 7529 652
rect 7581 600 7587 652
rect 7628 434 7656 1224
rect 7727 804 7733 856
rect 7785 804 7791 856
rect 7832 434 7860 1224
rect 7931 1008 7937 1060
rect 7989 1008 7995 1060
rect 8036 434 8064 1224
rect 8135 600 8141 652
rect 8193 600 8199 652
rect 8240 434 8268 1224
rect 8339 804 8345 856
rect 8397 804 8403 856
rect 8444 434 8472 1224
rect 8543 1008 8549 1060
rect 8601 1008 8607 1060
rect 8648 434 8676 1224
rect 8747 600 8753 652
rect 8805 600 8811 652
rect 8852 434 8880 1224
rect 8951 804 8957 856
rect 9009 804 9015 856
rect 9056 434 9084 1224
rect 9155 1008 9161 1060
rect 9213 1008 9219 1060
rect 9260 434 9288 1224
rect 9359 600 9365 652
rect 9417 600 9423 652
rect 9464 434 9492 1224
rect 9563 804 9569 856
rect 9621 804 9627 856
rect 9668 434 9696 1224
rect 9767 1008 9773 1060
rect 9825 1008 9831 1060
rect 62 382 68 434
rect 120 382 126 434
rect 266 382 272 434
rect 324 382 330 434
rect 470 382 476 434
rect 528 382 534 434
rect 674 382 680 434
rect 732 382 738 434
rect 878 382 884 434
rect 936 382 942 434
rect 1082 382 1088 434
rect 1140 382 1146 434
rect 1286 382 1292 434
rect 1344 382 1350 434
rect 1490 382 1496 434
rect 1548 382 1554 434
rect 1694 382 1700 434
rect 1752 382 1758 434
rect 1898 382 1904 434
rect 1956 382 1962 434
rect 2102 382 2108 434
rect 2160 382 2166 434
rect 2306 382 2312 434
rect 2364 382 2370 434
rect 2510 382 2516 434
rect 2568 382 2574 434
rect 2714 382 2720 434
rect 2772 382 2778 434
rect 2918 382 2924 434
rect 2976 382 2982 434
rect 3122 382 3128 434
rect 3180 382 3186 434
rect 3326 382 3332 434
rect 3384 382 3390 434
rect 3530 382 3536 434
rect 3588 382 3594 434
rect 3734 382 3740 434
rect 3792 382 3798 434
rect 3938 382 3944 434
rect 3996 382 4002 434
rect 4142 382 4148 434
rect 4200 382 4206 434
rect 4346 382 4352 434
rect 4404 382 4410 434
rect 4550 382 4556 434
rect 4608 382 4614 434
rect 4754 382 4760 434
rect 4812 382 4818 434
rect 4958 382 4964 434
rect 5016 382 5022 434
rect 5162 382 5168 434
rect 5220 382 5226 434
rect 5366 382 5372 434
rect 5424 382 5430 434
rect 5570 382 5576 434
rect 5628 382 5634 434
rect 5774 382 5780 434
rect 5832 382 5838 434
rect 5978 382 5984 434
rect 6036 382 6042 434
rect 6182 382 6188 434
rect 6240 382 6246 434
rect 6386 382 6392 434
rect 6444 382 6450 434
rect 6590 382 6596 434
rect 6648 382 6654 434
rect 6794 382 6800 434
rect 6852 382 6858 434
rect 6998 382 7004 434
rect 7056 382 7062 434
rect 7202 382 7208 434
rect 7260 382 7266 434
rect 7406 382 7412 434
rect 7464 382 7470 434
rect 7610 382 7616 434
rect 7668 382 7674 434
rect 7814 382 7820 434
rect 7872 382 7878 434
rect 8018 382 8024 434
rect 8076 382 8082 434
rect 8222 382 8228 434
rect 8280 382 8286 434
rect 8426 382 8432 434
rect 8484 382 8490 434
rect 8630 382 8636 434
rect 8688 382 8694 434
rect 8834 382 8840 434
rect 8892 382 8898 434
rect 9038 382 9044 434
rect 9096 382 9102 434
rect 9242 382 9248 434
rect 9300 382 9306 434
rect 9446 382 9452 434
rect 9504 382 9510 434
rect 9650 382 9656 434
rect 9708 382 9714 434
<< via1 >>
rect 178 1948 230 2000
rect 382 1948 434 2000
rect 586 1948 638 2000
rect 790 1948 842 2000
rect 994 1948 1046 2000
rect 1198 1948 1250 2000
rect 1402 1948 1454 2000
rect 1606 1948 1658 2000
rect 1810 1948 1862 2000
rect 2014 1948 2066 2000
rect 2218 1948 2270 2000
rect 2422 1948 2474 2000
rect 2626 1948 2678 2000
rect 2830 1948 2882 2000
rect 3034 1948 3086 2000
rect 3238 1948 3290 2000
rect 3442 1948 3494 2000
rect 3646 1948 3698 2000
rect 3850 1948 3902 2000
rect 4054 1948 4106 2000
rect 4258 1948 4310 2000
rect 4462 1948 4514 2000
rect 4666 1948 4718 2000
rect 4870 1948 4922 2000
rect 5074 1948 5126 2000
rect 5278 1948 5330 2000
rect 5482 1948 5534 2000
rect 5686 1948 5738 2000
rect 5890 1948 5942 2000
rect 6094 1948 6146 2000
rect 6298 1948 6350 2000
rect 6502 1948 6554 2000
rect 6706 1948 6758 2000
rect 6910 1948 6962 2000
rect 7114 1948 7166 2000
rect 7318 1948 7370 2000
rect 7522 1948 7574 2000
rect 7726 1948 7778 2000
rect 7930 1948 7982 2000
rect 8134 1948 8186 2000
rect 8338 1948 8390 2000
rect 8542 1948 8594 2000
rect 8746 1948 8798 2000
rect 8950 1948 9002 2000
rect 9154 1948 9206 2000
rect 9358 1948 9410 2000
rect 9562 1948 9614 2000
rect 9766 1948 9818 2000
rect 185 643 237 652
rect 185 609 194 643
rect 194 609 228 643
rect 228 609 237 643
rect 185 600 237 609
rect 389 847 441 856
rect 389 813 398 847
rect 398 813 432 847
rect 432 813 441 847
rect 389 804 441 813
rect 593 1051 645 1060
rect 593 1017 602 1051
rect 602 1017 636 1051
rect 636 1017 645 1051
rect 593 1008 645 1017
rect 797 643 849 652
rect 797 609 806 643
rect 806 609 840 643
rect 840 609 849 643
rect 797 600 849 609
rect 1001 847 1053 856
rect 1001 813 1010 847
rect 1010 813 1044 847
rect 1044 813 1053 847
rect 1001 804 1053 813
rect 1205 1051 1257 1060
rect 1205 1017 1214 1051
rect 1214 1017 1248 1051
rect 1248 1017 1257 1051
rect 1205 1008 1257 1017
rect 1409 643 1461 652
rect 1409 609 1418 643
rect 1418 609 1452 643
rect 1452 609 1461 643
rect 1409 600 1461 609
rect 1613 847 1665 856
rect 1613 813 1622 847
rect 1622 813 1656 847
rect 1656 813 1665 847
rect 1613 804 1665 813
rect 1817 1051 1869 1060
rect 1817 1017 1826 1051
rect 1826 1017 1860 1051
rect 1860 1017 1869 1051
rect 1817 1008 1869 1017
rect 2021 643 2073 652
rect 2021 609 2030 643
rect 2030 609 2064 643
rect 2064 609 2073 643
rect 2021 600 2073 609
rect 2225 847 2277 856
rect 2225 813 2234 847
rect 2234 813 2268 847
rect 2268 813 2277 847
rect 2225 804 2277 813
rect 2429 1051 2481 1060
rect 2429 1017 2438 1051
rect 2438 1017 2472 1051
rect 2472 1017 2481 1051
rect 2429 1008 2481 1017
rect 2633 643 2685 652
rect 2633 609 2642 643
rect 2642 609 2676 643
rect 2676 609 2685 643
rect 2633 600 2685 609
rect 2837 847 2889 856
rect 2837 813 2846 847
rect 2846 813 2880 847
rect 2880 813 2889 847
rect 2837 804 2889 813
rect 3041 1051 3093 1060
rect 3041 1017 3050 1051
rect 3050 1017 3084 1051
rect 3084 1017 3093 1051
rect 3041 1008 3093 1017
rect 3245 643 3297 652
rect 3245 609 3254 643
rect 3254 609 3288 643
rect 3288 609 3297 643
rect 3245 600 3297 609
rect 3449 847 3501 856
rect 3449 813 3458 847
rect 3458 813 3492 847
rect 3492 813 3501 847
rect 3449 804 3501 813
rect 3653 1051 3705 1060
rect 3653 1017 3662 1051
rect 3662 1017 3696 1051
rect 3696 1017 3705 1051
rect 3653 1008 3705 1017
rect 3857 643 3909 652
rect 3857 609 3866 643
rect 3866 609 3900 643
rect 3900 609 3909 643
rect 3857 600 3909 609
rect 4061 847 4113 856
rect 4061 813 4070 847
rect 4070 813 4104 847
rect 4104 813 4113 847
rect 4061 804 4113 813
rect 4265 1051 4317 1060
rect 4265 1017 4274 1051
rect 4274 1017 4308 1051
rect 4308 1017 4317 1051
rect 4265 1008 4317 1017
rect 4469 643 4521 652
rect 4469 609 4478 643
rect 4478 609 4512 643
rect 4512 609 4521 643
rect 4469 600 4521 609
rect 4673 847 4725 856
rect 4673 813 4682 847
rect 4682 813 4716 847
rect 4716 813 4725 847
rect 4673 804 4725 813
rect 4877 1051 4929 1060
rect 4877 1017 4886 1051
rect 4886 1017 4920 1051
rect 4920 1017 4929 1051
rect 4877 1008 4929 1017
rect 5081 643 5133 652
rect 5081 609 5090 643
rect 5090 609 5124 643
rect 5124 609 5133 643
rect 5081 600 5133 609
rect 5285 847 5337 856
rect 5285 813 5294 847
rect 5294 813 5328 847
rect 5328 813 5337 847
rect 5285 804 5337 813
rect 5489 1051 5541 1060
rect 5489 1017 5498 1051
rect 5498 1017 5532 1051
rect 5532 1017 5541 1051
rect 5489 1008 5541 1017
rect 5693 643 5745 652
rect 5693 609 5702 643
rect 5702 609 5736 643
rect 5736 609 5745 643
rect 5693 600 5745 609
rect 5897 847 5949 856
rect 5897 813 5906 847
rect 5906 813 5940 847
rect 5940 813 5949 847
rect 5897 804 5949 813
rect 6101 1051 6153 1060
rect 6101 1017 6110 1051
rect 6110 1017 6144 1051
rect 6144 1017 6153 1051
rect 6101 1008 6153 1017
rect 6305 643 6357 652
rect 6305 609 6314 643
rect 6314 609 6348 643
rect 6348 609 6357 643
rect 6305 600 6357 609
rect 6509 847 6561 856
rect 6509 813 6518 847
rect 6518 813 6552 847
rect 6552 813 6561 847
rect 6509 804 6561 813
rect 6713 1051 6765 1060
rect 6713 1017 6722 1051
rect 6722 1017 6756 1051
rect 6756 1017 6765 1051
rect 6713 1008 6765 1017
rect 6917 643 6969 652
rect 6917 609 6926 643
rect 6926 609 6960 643
rect 6960 609 6969 643
rect 6917 600 6969 609
rect 7121 847 7173 856
rect 7121 813 7130 847
rect 7130 813 7164 847
rect 7164 813 7173 847
rect 7121 804 7173 813
rect 7325 1051 7377 1060
rect 7325 1017 7334 1051
rect 7334 1017 7368 1051
rect 7368 1017 7377 1051
rect 7325 1008 7377 1017
rect 7529 643 7581 652
rect 7529 609 7538 643
rect 7538 609 7572 643
rect 7572 609 7581 643
rect 7529 600 7581 609
rect 7733 847 7785 856
rect 7733 813 7742 847
rect 7742 813 7776 847
rect 7776 813 7785 847
rect 7733 804 7785 813
rect 7937 1051 7989 1060
rect 7937 1017 7946 1051
rect 7946 1017 7980 1051
rect 7980 1017 7989 1051
rect 7937 1008 7989 1017
rect 8141 643 8193 652
rect 8141 609 8150 643
rect 8150 609 8184 643
rect 8184 609 8193 643
rect 8141 600 8193 609
rect 8345 847 8397 856
rect 8345 813 8354 847
rect 8354 813 8388 847
rect 8388 813 8397 847
rect 8345 804 8397 813
rect 8549 1051 8601 1060
rect 8549 1017 8558 1051
rect 8558 1017 8592 1051
rect 8592 1017 8601 1051
rect 8549 1008 8601 1017
rect 8753 643 8805 652
rect 8753 609 8762 643
rect 8762 609 8796 643
rect 8796 609 8805 643
rect 8753 600 8805 609
rect 8957 847 9009 856
rect 8957 813 8966 847
rect 8966 813 9000 847
rect 9000 813 9009 847
rect 8957 804 9009 813
rect 9161 1051 9213 1060
rect 9161 1017 9170 1051
rect 9170 1017 9204 1051
rect 9204 1017 9213 1051
rect 9161 1008 9213 1017
rect 9365 643 9417 652
rect 9365 609 9374 643
rect 9374 609 9408 643
rect 9408 609 9417 643
rect 9365 600 9417 609
rect 9569 847 9621 856
rect 9569 813 9578 847
rect 9578 813 9612 847
rect 9612 813 9621 847
rect 9569 804 9621 813
rect 9773 1051 9825 1060
rect 9773 1017 9782 1051
rect 9782 1017 9816 1051
rect 9816 1017 9825 1051
rect 9773 1008 9825 1017
rect 68 382 120 434
rect 272 382 324 434
rect 476 382 528 434
rect 680 382 732 434
rect 884 382 936 434
rect 1088 382 1140 434
rect 1292 382 1344 434
rect 1496 382 1548 434
rect 1700 382 1752 434
rect 1904 382 1956 434
rect 2108 382 2160 434
rect 2312 382 2364 434
rect 2516 382 2568 434
rect 2720 382 2772 434
rect 2924 382 2976 434
rect 3128 382 3180 434
rect 3332 382 3384 434
rect 3536 382 3588 434
rect 3740 382 3792 434
rect 3944 382 3996 434
rect 4148 382 4200 434
rect 4352 382 4404 434
rect 4556 382 4608 434
rect 4760 382 4812 434
rect 4964 382 5016 434
rect 5168 382 5220 434
rect 5372 382 5424 434
rect 5576 382 5628 434
rect 5780 382 5832 434
rect 5984 382 6036 434
rect 6188 382 6240 434
rect 6392 382 6444 434
rect 6596 382 6648 434
rect 6800 382 6852 434
rect 7004 382 7056 434
rect 7208 382 7260 434
rect 7412 382 7464 434
rect 7616 382 7668 434
rect 7820 382 7872 434
rect 8024 382 8076 434
rect 8228 382 8280 434
rect 8432 382 8484 434
rect 8636 382 8688 434
rect 8840 382 8892 434
rect 9044 382 9096 434
rect 9248 382 9300 434
rect 9452 382 9504 434
rect 9656 382 9708 434
<< metal2 >>
rect 26 2000 9832 2006
rect 26 1948 178 2000
rect 230 1948 382 2000
rect 434 1948 586 2000
rect 638 1948 790 2000
rect 842 1948 994 2000
rect 1046 1948 1198 2000
rect 1250 1948 1402 2000
rect 1454 1948 1606 2000
rect 1658 1948 1810 2000
rect 1862 1948 2014 2000
rect 2066 1948 2218 2000
rect 2270 1948 2422 2000
rect 2474 1948 2626 2000
rect 2678 1948 2830 2000
rect 2882 1948 3034 2000
rect 3086 1948 3238 2000
rect 3290 1948 3442 2000
rect 3494 1948 3646 2000
rect 3698 1948 3850 2000
rect 3902 1948 4054 2000
rect 4106 1948 4258 2000
rect 4310 1948 4462 2000
rect 4514 1948 4666 2000
rect 4718 1948 4870 2000
rect 4922 1948 5074 2000
rect 5126 1948 5278 2000
rect 5330 1948 5482 2000
rect 5534 1948 5686 2000
rect 5738 1948 5890 2000
rect 5942 1948 6094 2000
rect 6146 1948 6298 2000
rect 6350 1948 6502 2000
rect 6554 1948 6706 2000
rect 6758 1948 6910 2000
rect 6962 1948 7114 2000
rect 7166 1948 7318 2000
rect 7370 1948 7522 2000
rect 7574 1948 7726 2000
rect 7778 1948 7930 2000
rect 7982 1948 8134 2000
rect 8186 1948 8338 2000
rect 8390 1948 8542 2000
rect 8594 1948 8746 2000
rect 8798 1948 8950 2000
rect 9002 1948 9154 2000
rect 9206 1948 9358 2000
rect 9410 1948 9562 2000
rect 9614 1948 9766 2000
rect 9818 1948 9832 2000
rect 26 1942 9832 1948
rect 587 1048 593 1060
rect 0 1020 593 1048
rect 587 1008 593 1020
rect 645 1048 651 1060
rect 1199 1048 1205 1060
rect 645 1020 1205 1048
rect 645 1008 651 1020
rect 1199 1008 1205 1020
rect 1257 1048 1263 1060
rect 1811 1048 1817 1060
rect 1257 1020 1817 1048
rect 1257 1008 1263 1020
rect 1811 1008 1817 1020
rect 1869 1048 1875 1060
rect 2423 1048 2429 1060
rect 1869 1020 2429 1048
rect 1869 1008 1875 1020
rect 2423 1008 2429 1020
rect 2481 1048 2487 1060
rect 3035 1048 3041 1060
rect 2481 1020 3041 1048
rect 2481 1008 2487 1020
rect 3035 1008 3041 1020
rect 3093 1048 3099 1060
rect 3647 1048 3653 1060
rect 3093 1020 3653 1048
rect 3093 1008 3099 1020
rect 3647 1008 3653 1020
rect 3705 1048 3711 1060
rect 4259 1048 4265 1060
rect 3705 1020 4265 1048
rect 3705 1008 3711 1020
rect 4259 1008 4265 1020
rect 4317 1048 4323 1060
rect 4871 1048 4877 1060
rect 4317 1020 4877 1048
rect 4317 1008 4323 1020
rect 4871 1008 4877 1020
rect 4929 1048 4935 1060
rect 5483 1048 5489 1060
rect 4929 1020 5489 1048
rect 4929 1008 4935 1020
rect 5483 1008 5489 1020
rect 5541 1048 5547 1060
rect 6095 1048 6101 1060
rect 5541 1020 6101 1048
rect 5541 1008 5547 1020
rect 6095 1008 6101 1020
rect 6153 1048 6159 1060
rect 6707 1048 6713 1060
rect 6153 1020 6713 1048
rect 6153 1008 6159 1020
rect 6707 1008 6713 1020
rect 6765 1048 6771 1060
rect 7319 1048 7325 1060
rect 6765 1020 7325 1048
rect 6765 1008 6771 1020
rect 7319 1008 7325 1020
rect 7377 1048 7383 1060
rect 7931 1048 7937 1060
rect 7377 1020 7937 1048
rect 7377 1008 7383 1020
rect 7931 1008 7937 1020
rect 7989 1048 7995 1060
rect 8543 1048 8549 1060
rect 7989 1020 8549 1048
rect 7989 1008 7995 1020
rect 8543 1008 8549 1020
rect 8601 1048 8607 1060
rect 9155 1048 9161 1060
rect 8601 1020 9161 1048
rect 8601 1008 8607 1020
rect 9155 1008 9161 1020
rect 9213 1048 9219 1060
rect 9767 1048 9773 1060
rect 9213 1020 9773 1048
rect 9213 1008 9219 1020
rect 9767 1008 9773 1020
rect 9825 1008 9831 1060
rect 383 844 389 856
rect 0 816 389 844
rect 383 804 389 816
rect 441 844 447 856
rect 995 844 1001 856
rect 441 816 1001 844
rect 441 804 447 816
rect 995 804 1001 816
rect 1053 844 1059 856
rect 1607 844 1613 856
rect 1053 816 1613 844
rect 1053 804 1059 816
rect 1607 804 1613 816
rect 1665 844 1671 856
rect 2219 844 2225 856
rect 1665 816 2225 844
rect 1665 804 1671 816
rect 2219 804 2225 816
rect 2277 844 2283 856
rect 2831 844 2837 856
rect 2277 816 2837 844
rect 2277 804 2283 816
rect 2831 804 2837 816
rect 2889 844 2895 856
rect 3443 844 3449 856
rect 2889 816 3449 844
rect 2889 804 2895 816
rect 3443 804 3449 816
rect 3501 844 3507 856
rect 4055 844 4061 856
rect 3501 816 4061 844
rect 3501 804 3507 816
rect 4055 804 4061 816
rect 4113 844 4119 856
rect 4667 844 4673 856
rect 4113 816 4673 844
rect 4113 804 4119 816
rect 4667 804 4673 816
rect 4725 844 4731 856
rect 5279 844 5285 856
rect 4725 816 5285 844
rect 4725 804 4731 816
rect 5279 804 5285 816
rect 5337 844 5343 856
rect 5891 844 5897 856
rect 5337 816 5897 844
rect 5337 804 5343 816
rect 5891 804 5897 816
rect 5949 844 5955 856
rect 6503 844 6509 856
rect 5949 816 6509 844
rect 5949 804 5955 816
rect 6503 804 6509 816
rect 6561 844 6567 856
rect 7115 844 7121 856
rect 6561 816 7121 844
rect 6561 804 6567 816
rect 7115 804 7121 816
rect 7173 844 7179 856
rect 7727 844 7733 856
rect 7173 816 7733 844
rect 7173 804 7179 816
rect 7727 804 7733 816
rect 7785 844 7791 856
rect 8339 844 8345 856
rect 7785 816 8345 844
rect 7785 804 7791 816
rect 8339 804 8345 816
rect 8397 844 8403 856
rect 8951 844 8957 856
rect 8397 816 8957 844
rect 8397 804 8403 816
rect 8951 804 8957 816
rect 9009 844 9015 856
rect 9563 844 9569 856
rect 9009 816 9569 844
rect 9009 804 9015 816
rect 9563 804 9569 816
rect 9621 844 9627 856
rect 9621 816 9792 844
rect 9621 804 9627 816
rect 179 640 185 652
rect 0 612 185 640
rect 179 600 185 612
rect 237 640 243 652
rect 791 640 797 652
rect 237 612 797 640
rect 237 600 243 612
rect 791 600 797 612
rect 849 640 855 652
rect 1403 640 1409 652
rect 849 612 1409 640
rect 849 600 855 612
rect 1403 600 1409 612
rect 1461 640 1467 652
rect 2015 640 2021 652
rect 1461 612 2021 640
rect 1461 600 1467 612
rect 2015 600 2021 612
rect 2073 640 2079 652
rect 2627 640 2633 652
rect 2073 612 2633 640
rect 2073 600 2079 612
rect 2627 600 2633 612
rect 2685 640 2691 652
rect 3239 640 3245 652
rect 2685 612 3245 640
rect 2685 600 2691 612
rect 3239 600 3245 612
rect 3297 640 3303 652
rect 3851 640 3857 652
rect 3297 612 3857 640
rect 3297 600 3303 612
rect 3851 600 3857 612
rect 3909 640 3915 652
rect 4463 640 4469 652
rect 3909 612 4469 640
rect 3909 600 3915 612
rect 4463 600 4469 612
rect 4521 640 4527 652
rect 5075 640 5081 652
rect 4521 612 5081 640
rect 4521 600 4527 612
rect 5075 600 5081 612
rect 5133 640 5139 652
rect 5687 640 5693 652
rect 5133 612 5693 640
rect 5133 600 5139 612
rect 5687 600 5693 612
rect 5745 640 5751 652
rect 6299 640 6305 652
rect 5745 612 6305 640
rect 5745 600 5751 612
rect 6299 600 6305 612
rect 6357 640 6363 652
rect 6911 640 6917 652
rect 6357 612 6917 640
rect 6357 600 6363 612
rect 6911 600 6917 612
rect 6969 640 6975 652
rect 7523 640 7529 652
rect 6969 612 7529 640
rect 6969 600 6975 612
rect 7523 600 7529 612
rect 7581 640 7587 652
rect 8135 640 8141 652
rect 7581 612 8141 640
rect 7581 600 7587 612
rect 8135 600 8141 612
rect 8193 640 8199 652
rect 8747 640 8753 652
rect 8193 612 8753 640
rect 8193 600 8199 612
rect 8747 600 8753 612
rect 8805 640 8811 652
rect 9359 640 9365 652
rect 8805 612 9365 640
rect 8805 600 8811 612
rect 9359 600 9365 612
rect 9417 640 9423 652
rect 9417 612 9792 640
rect 9417 600 9423 612
rect 62 382 68 434
rect 120 422 126 434
rect 266 422 272 434
rect 120 394 272 422
rect 120 382 126 394
rect 266 382 272 394
rect 324 422 330 434
rect 470 422 476 434
rect 324 394 476 422
rect 324 382 330 394
rect 470 382 476 394
rect 528 382 534 434
rect 674 382 680 434
rect 732 422 738 434
rect 878 422 884 434
rect 732 394 884 422
rect 732 382 738 394
rect 878 382 884 394
rect 936 422 942 434
rect 1082 422 1088 434
rect 936 394 1088 422
rect 936 382 942 394
rect 1082 382 1088 394
rect 1140 382 1146 434
rect 1286 382 1292 434
rect 1344 422 1350 434
rect 1490 422 1496 434
rect 1344 394 1496 422
rect 1344 382 1350 394
rect 1490 382 1496 394
rect 1548 422 1554 434
rect 1694 422 1700 434
rect 1548 394 1700 422
rect 1548 382 1554 394
rect 1694 382 1700 394
rect 1752 382 1758 434
rect 1898 382 1904 434
rect 1956 422 1962 434
rect 2102 422 2108 434
rect 1956 394 2108 422
rect 1956 382 1962 394
rect 2102 382 2108 394
rect 2160 422 2166 434
rect 2306 422 2312 434
rect 2160 394 2312 422
rect 2160 382 2166 394
rect 2306 382 2312 394
rect 2364 382 2370 434
rect 2510 382 2516 434
rect 2568 422 2574 434
rect 2714 422 2720 434
rect 2568 394 2720 422
rect 2568 382 2574 394
rect 2714 382 2720 394
rect 2772 422 2778 434
rect 2918 422 2924 434
rect 2772 394 2924 422
rect 2772 382 2778 394
rect 2918 382 2924 394
rect 2976 382 2982 434
rect 3122 382 3128 434
rect 3180 422 3186 434
rect 3326 422 3332 434
rect 3180 394 3332 422
rect 3180 382 3186 394
rect 3326 382 3332 394
rect 3384 422 3390 434
rect 3530 422 3536 434
rect 3384 394 3536 422
rect 3384 382 3390 394
rect 3530 382 3536 394
rect 3588 382 3594 434
rect 3734 382 3740 434
rect 3792 422 3798 434
rect 3938 422 3944 434
rect 3792 394 3944 422
rect 3792 382 3798 394
rect 3938 382 3944 394
rect 3996 422 4002 434
rect 4142 422 4148 434
rect 3996 394 4148 422
rect 3996 382 4002 394
rect 4142 382 4148 394
rect 4200 382 4206 434
rect 4346 382 4352 434
rect 4404 422 4410 434
rect 4550 422 4556 434
rect 4404 394 4556 422
rect 4404 382 4410 394
rect 4550 382 4556 394
rect 4608 422 4614 434
rect 4754 422 4760 434
rect 4608 394 4760 422
rect 4608 382 4614 394
rect 4754 382 4760 394
rect 4812 382 4818 434
rect 4958 382 4964 434
rect 5016 422 5022 434
rect 5162 422 5168 434
rect 5016 394 5168 422
rect 5016 382 5022 394
rect 5162 382 5168 394
rect 5220 422 5226 434
rect 5366 422 5372 434
rect 5220 394 5372 422
rect 5220 382 5226 394
rect 5366 382 5372 394
rect 5424 382 5430 434
rect 5570 382 5576 434
rect 5628 422 5634 434
rect 5774 422 5780 434
rect 5628 394 5780 422
rect 5628 382 5634 394
rect 5774 382 5780 394
rect 5832 422 5838 434
rect 5978 422 5984 434
rect 5832 394 5984 422
rect 5832 382 5838 394
rect 5978 382 5984 394
rect 6036 382 6042 434
rect 6182 382 6188 434
rect 6240 422 6246 434
rect 6386 422 6392 434
rect 6240 394 6392 422
rect 6240 382 6246 394
rect 6386 382 6392 394
rect 6444 422 6450 434
rect 6590 422 6596 434
rect 6444 394 6596 422
rect 6444 382 6450 394
rect 6590 382 6596 394
rect 6648 382 6654 434
rect 6794 382 6800 434
rect 6852 422 6858 434
rect 6998 422 7004 434
rect 6852 394 7004 422
rect 6852 382 6858 394
rect 6998 382 7004 394
rect 7056 422 7062 434
rect 7202 422 7208 434
rect 7056 394 7208 422
rect 7056 382 7062 394
rect 7202 382 7208 394
rect 7260 382 7266 434
rect 7406 382 7412 434
rect 7464 422 7470 434
rect 7610 422 7616 434
rect 7464 394 7616 422
rect 7464 382 7470 394
rect 7610 382 7616 394
rect 7668 422 7674 434
rect 7814 422 7820 434
rect 7668 394 7820 422
rect 7668 382 7674 394
rect 7814 382 7820 394
rect 7872 382 7878 434
rect 8018 382 8024 434
rect 8076 422 8082 434
rect 8222 422 8228 434
rect 8076 394 8228 422
rect 8076 382 8082 394
rect 8222 382 8228 394
rect 8280 422 8286 434
rect 8426 422 8432 434
rect 8280 394 8432 422
rect 8280 382 8286 394
rect 8426 382 8432 394
rect 8484 382 8490 434
rect 8630 382 8636 434
rect 8688 422 8694 434
rect 8834 422 8840 434
rect 8688 394 8840 422
rect 8688 382 8694 394
rect 8834 382 8840 394
rect 8892 422 8898 434
rect 9038 422 9044 434
rect 8892 394 9044 422
rect 8892 382 8898 394
rect 9038 382 9044 394
rect 9096 382 9102 434
rect 9242 382 9248 434
rect 9300 422 9306 434
rect 9446 422 9452 434
rect 9300 394 9452 422
rect 9300 382 9306 394
rect 9446 382 9452 394
rect 9504 422 9510 434
rect 9650 422 9656 434
rect 9504 394 9656 422
rect 9504 382 9510 394
rect 9650 382 9656 394
rect 9708 382 9714 434
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_0
timestamp 1581321264
transform 1 0 9588 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_1
timestamp 1581321264
transform 1 0 9384 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_2
timestamp 1581321264
transform 1 0 9180 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_3
timestamp 1581321264
transform 1 0 8976 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_4
timestamp 1581321264
transform 1 0 8772 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_5
timestamp 1581321264
transform 1 0 8568 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_6
timestamp 1581321264
transform 1 0 8364 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_7
timestamp 1581321264
transform 1 0 8160 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_8
timestamp 1581321264
transform 1 0 7956 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_9
timestamp 1581321264
transform 1 0 7752 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_10
timestamp 1581321264
transform 1 0 7548 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_11
timestamp 1581321264
transform 1 0 7344 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_12
timestamp 1581321264
transform 1 0 7140 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_13
timestamp 1581321264
transform 1 0 6936 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_14
timestamp 1581321264
transform 1 0 6732 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_15
timestamp 1581321264
transform 1 0 6528 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_16
timestamp 1581321264
transform 1 0 6324 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_17
timestamp 1581321264
transform 1 0 6120 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_18
timestamp 1581321264
transform 1 0 5916 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_19
timestamp 1581321264
transform 1 0 5712 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_20
timestamp 1581321264
transform 1 0 5508 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_21
timestamp 1581321264
transform 1 0 5304 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_22
timestamp 1581321264
transform 1 0 5100 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_23
timestamp 1581321264
transform 1 0 4896 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_24
timestamp 1581321264
transform 1 0 4692 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_25
timestamp 1581321264
transform 1 0 4488 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_26
timestamp 1581321264
transform 1 0 4284 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_27
timestamp 1581321264
transform 1 0 4080 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_28
timestamp 1581321264
transform 1 0 3876 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_29
timestamp 1581321264
transform 1 0 3672 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_30
timestamp 1581321264
transform 1 0 3468 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_31
timestamp 1581321264
transform 1 0 3264 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_32
timestamp 1581321264
transform 1 0 3060 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_33
timestamp 1581321264
transform 1 0 2856 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_34
timestamp 1581321264
transform 1 0 2652 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_35
timestamp 1581321264
transform 1 0 2448 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_36
timestamp 1581321264
transform 1 0 2244 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_37
timestamp 1581321264
transform 1 0 2040 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_38
timestamp 1581321264
transform 1 0 1836 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_39
timestamp 1581321264
transform 1 0 1632 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_40
timestamp 1581321264
transform 1 0 1428 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_41
timestamp 1581321264
transform 1 0 1224 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_42
timestamp 1581321264
transform 1 0 1020 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_43
timestamp 1581321264
transform 1 0 816 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_44
timestamp 1581321264
transform 1 0 612 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_45
timestamp 1581321264
transform 1 0 408 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_46
timestamp 1581321264
transform 1 0 204 0 1 1224
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_47
timestamp 1581321264
transform 1 0 0 0 1 1224
box 1 0 255 817
<< labels >>
rlabel metal2 s 0 612 9792 640 4 sel_0
port 3 nsew
rlabel metal2 s 0 816 9792 844 4 sel_1
port 5 nsew
rlabel metal2 s 0 1020 9792 1048 4 sel_2
port 7 nsew
rlabel metal1 s 80 408 108 1224 4 bl_out_0
port 9 nsew
rlabel metal1 s 692 408 720 1224 4 bl_out_1
port 11 nsew
rlabel metal1 s 1304 408 1332 1224 4 bl_out_2
port 13 nsew
rlabel metal1 s 1916 408 1944 1224 4 bl_out_3
port 15 nsew
rlabel metal1 s 2528 408 2556 1224 4 bl_out_4
port 17 nsew
rlabel metal1 s 3140 408 3168 1224 4 bl_out_5
port 19 nsew
rlabel metal1 s 3752 408 3780 1224 4 bl_out_6
port 21 nsew
rlabel metal1 s 4364 408 4392 1224 4 bl_out_7
port 23 nsew
rlabel metal1 s 4976 408 5004 1224 4 bl_out_8
port 25 nsew
rlabel metal1 s 5588 408 5616 1224 4 bl_out_9
port 27 nsew
rlabel metal1 s 6200 408 6228 1224 4 bl_out_10
port 29 nsew
rlabel metal1 s 6812 408 6840 1224 4 bl_out_11
port 31 nsew
rlabel metal1 s 7424 408 7452 1224 4 bl_out_12
port 33 nsew
rlabel metal1 s 8036 408 8064 1224 4 bl_out_13
port 35 nsew
rlabel metal1 s 8648 408 8676 1224 4 bl_out_14
port 37 nsew
rlabel metal1 s 9260 408 9288 1224 4 bl_out_15
port 39 nsew
rlabel metal2 s 26 1942 9832 2006 4 gnd
port 41 nsew
rlabel metal1 s 80 1854 108 2006 4 bl_0
port 43 nsew
rlabel metal1 s 284 1854 312 2006 4 bl_1
port 45 nsew
rlabel metal1 s 488 1854 516 2006 4 bl_2
port 47 nsew
rlabel metal1 s 692 1854 720 2006 4 bl_3
port 49 nsew
rlabel metal1 s 896 1854 924 2006 4 bl_4
port 51 nsew
rlabel metal1 s 1100 1854 1128 2006 4 bl_5
port 53 nsew
rlabel metal1 s 1304 1854 1332 2006 4 bl_6
port 55 nsew
rlabel metal1 s 1508 1854 1536 2006 4 bl_7
port 57 nsew
rlabel metal1 s 1712 1854 1740 2006 4 bl_8
port 59 nsew
rlabel metal1 s 1916 1854 1944 2006 4 bl_9
port 61 nsew
rlabel metal1 s 2120 1854 2148 2006 4 bl_10
port 63 nsew
rlabel metal1 s 2324 1854 2352 2006 4 bl_11
port 65 nsew
rlabel metal1 s 2528 1854 2556 2006 4 bl_12
port 67 nsew
rlabel metal1 s 2732 1854 2760 2006 4 bl_13
port 69 nsew
rlabel metal1 s 2936 1854 2964 2006 4 bl_14
port 71 nsew
rlabel metal1 s 3140 1854 3168 2006 4 bl_15
port 73 nsew
rlabel metal1 s 3344 1854 3372 2006 4 bl_16
port 75 nsew
rlabel metal1 s 3548 1854 3576 2006 4 bl_17
port 77 nsew
rlabel metal1 s 3752 1854 3780 2006 4 bl_18
port 79 nsew
rlabel metal1 s 3956 1854 3984 2006 4 bl_19
port 81 nsew
rlabel metal1 s 4160 1854 4188 2006 4 bl_20
port 83 nsew
rlabel metal1 s 4364 1854 4392 2006 4 bl_21
port 85 nsew
rlabel metal1 s 4568 1854 4596 2006 4 bl_22
port 87 nsew
rlabel metal1 s 4772 1854 4800 2006 4 bl_23
port 89 nsew
rlabel metal1 s 4976 1854 5004 2006 4 bl_24
port 91 nsew
rlabel metal1 s 5180 1854 5208 2006 4 bl_25
port 93 nsew
rlabel metal1 s 5384 1854 5412 2006 4 bl_26
port 95 nsew
rlabel metal1 s 5588 1854 5616 2006 4 bl_27
port 97 nsew
rlabel metal1 s 5792 1854 5820 2006 4 bl_28
port 99 nsew
rlabel metal1 s 5996 1854 6024 2006 4 bl_29
port 101 nsew
rlabel metal1 s 6200 1854 6228 2006 4 bl_30
port 103 nsew
rlabel metal1 s 6404 1854 6432 2006 4 bl_31
port 105 nsew
rlabel metal1 s 6608 1854 6636 2006 4 bl_32
port 107 nsew
rlabel metal1 s 6812 1854 6840 2006 4 bl_33
port 109 nsew
rlabel metal1 s 7016 1854 7044 2006 4 bl_34
port 111 nsew
rlabel metal1 s 7220 1854 7248 2006 4 bl_35
port 113 nsew
rlabel metal1 s 7424 1854 7452 2006 4 bl_36
port 115 nsew
rlabel metal1 s 7628 1854 7656 2006 4 bl_37
port 117 nsew
rlabel metal1 s 7832 1854 7860 2006 4 bl_38
port 119 nsew
rlabel metal1 s 8036 1854 8064 2006 4 bl_39
port 121 nsew
rlabel metal1 s 8240 1854 8268 2006 4 bl_40
port 123 nsew
rlabel metal1 s 8444 1854 8472 2006 4 bl_41
port 125 nsew
rlabel metal1 s 8648 1854 8676 2006 4 bl_42
port 127 nsew
rlabel metal1 s 8852 1854 8880 2006 4 bl_43
port 129 nsew
rlabel metal1 s 9056 1854 9084 2006 4 bl_44
port 131 nsew
rlabel metal1 s 9260 1854 9288 2006 4 bl_45
port 133 nsew
rlabel metal1 s 9464 1854 9492 2006 4 bl_46
port 135 nsew
rlabel metal1 s 9668 1854 9696 2006 4 bl_47
port 137 nsew
<< properties >>
string FIXED_BBOX 0 0 9792 981
<< end >>
