magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1308 -1216 2171 4388
<< locali >>
rect 194 60 260 94
rect 602 60 668 94
<< metal1 >>
rect 0 2833 817 2861
rect 0 2408 844 2436
rect 0 2160 816 2188
rect 0 1881 817 1909
rect 0 1456 844 1484
rect 0 844 816 872
rect 0 222 844 250
<< metal2 >>
rect 189 3098 217 3126
rect 329 3098 357 3126
rect 597 3098 625 3126
rect 737 3098 765 3126
use sky130_rom_krom_rom_address_control_buf  sky130_rom_krom_rom_address_control_buf_0
timestamp 1581321264
transform -1 0 816 0 1 0
box -95 44 456 3128
use sky130_rom_krom_rom_address_control_buf  sky130_rom_krom_rom_address_control_buf_1
timestamp 1581321264
transform -1 0 408 0 1 0
box -95 44 456 3128
<< labels >>
rlabel metal1 s 0 2160 816 2188 4 clk
port 3 nsew
rlabel metal1 s 0 2833 28 2861 4 vdd
port 5 nsew
rlabel metal1 s 0 1881 28 1909 4 vdd
port 5 nsew
rlabel metal1 s 0 844 28 872 4 vdd
port 5 nsew
rlabel metal1 s 816 2408 844 2436 4 gnd
port 7 nsew
rlabel metal1 s 816 1456 844 1484 4 gnd
port 7 nsew
rlabel metal1 s 816 222 844 250 4 gnd
port 7 nsew
rlabel metal2 s 189 3098 217 3126 4 A0_out
port 9 nsew
rlabel metal2 s 329 3098 357 3126 4 Abar0_out
port 11 nsew
rlabel locali s 227 77 227 77 4 A0_in
port 12 nsew
rlabel metal2 s 597 3098 625 3126 4 A1_out
port 14 nsew
rlabel metal2 s 737 3098 765 3126 4 Abar1_out
port 16 nsew
rlabel locali s 635 77 635 77 4 A1_in
port 17 nsew
<< properties >>
string FIXED_BBOX 0 0 816 3098
<< end >>
