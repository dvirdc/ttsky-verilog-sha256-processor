magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1216 -1310 2472 2071
<< nwell >>
rect 774 -50 942 118
<< pwell >>
rect 169 -17 303 85
<< psubdiff >>
rect 195 51 277 59
rect 195 17 219 51
rect 253 17 277 51
rect 195 9 277 17
<< nsubdiff >>
rect 817 51 899 59
rect 817 17 841 51
rect 875 17 899 51
rect 817 9 899 17
<< psubdiffcont >>
rect 219 17 253 51
<< nsubdiffcont >>
rect 841 17 875 51
<< locali >>
rect 60 563 94 629
rect 1160 546 1194 613
rect 60 359 94 425
rect 1160 342 1194 409
rect 60 155 94 221
rect 1160 138 1194 205
rect 203 17 219 51
rect 253 17 269 51
rect 825 17 841 51
rect 875 17 891 51
<< viali >>
rect 219 17 253 51
rect 841 17 875 51
<< metal1 >>
rect 222 63 250 730
rect 844 63 872 730
rect 213 51 259 63
rect 213 17 219 51
rect 253 17 259 51
rect 213 5 259 17
rect 835 51 881 63
rect 835 17 841 51
rect 875 17 881 51
rect 835 5 881 17
use sky130_rom_krom_pinv_dec_2  sky130_rom_krom_pinv_dec_2_0
timestamp 1581321264
transform 1 0 0 0 1 512
box 44 -50 1212 299
use sky130_rom_krom_pinv_dec_2  sky130_rom_krom_pinv_dec_2_1
timestamp 1581321264
transform 1 0 0 0 1 308
box 44 -50 1212 299
use sky130_rom_krom_pinv_dec_2  sky130_rom_krom_pinv_dec_2_2
timestamp 1581321264
transform 1 0 0 0 1 104
box 44 -50 1212 299
<< labels >>
rlabel locali s 77 188 77 188 4 in_0
port 2 nsew
rlabel locali s 1177 188 1177 188 4 out_0
port 3 nsew
rlabel locali s 77 392 77 392 4 in_1
port 4 nsew
rlabel locali s 1177 392 1177 392 4 out_1
port 5 nsew
rlabel locali s 77 596 77 596 4 in_2
port 6 nsew
rlabel locali s 1177 596 1177 596 4 out_2
port 7 nsew
rlabel metal1 s 222 6 250 34 4 gnd
port 9 nsew
rlabel metal1 s 222 702 250 730 4 gnd
port 9 nsew
rlabel metal1 s 844 702 872 730 4 vdd
port 11 nsew
rlabel metal1 s 844 6 872 34 4 vdd
port 11 nsew
<< properties >>
string FIXED_BBOX 774 -50 942 0
<< end >>
