magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1296 -1277 1664 3436
<< nwell >>
rect -36 1017 404 2176
<< pwell >>
rect 232 149 334 159
rect 28 25 334 149
<< scnmos >>
rect 114 51 144 123
<< scpmos >>
rect 114 1844 144 2068
<< ndiff >>
rect 54 104 114 123
rect 54 70 62 104
rect 96 70 114 104
rect 54 51 114 70
rect 144 104 204 123
rect 144 70 162 104
rect 196 70 204 104
rect 144 51 204 70
<< pdiff >>
rect 54 1973 114 2068
rect 54 1939 62 1973
rect 96 1939 114 1973
rect 54 1844 114 1939
rect 144 1973 204 2068
rect 144 1939 162 1973
rect 196 1939 204 1973
rect 144 1844 204 1939
<< ndiffc >>
rect 62 70 96 104
rect 162 70 196 104
<< pdiffc >>
rect 62 1939 96 1973
rect 162 1939 196 1973
<< psubdiff >>
rect 258 109 308 133
rect 258 75 266 109
rect 300 75 308 109
rect 258 51 308 75
<< nsubdiff >>
rect 258 2031 308 2055
rect 258 1997 266 2031
rect 300 1997 308 2031
rect 258 1973 308 1997
<< psubdiffcont >>
rect 266 75 300 109
<< nsubdiffcont >>
rect 266 1997 300 2031
<< poly >>
rect 114 2068 144 2094
rect 114 1054 144 1844
rect 48 1038 144 1054
rect 48 1004 64 1038
rect 98 1004 144 1038
rect 48 988 144 1004
rect 114 123 144 988
rect 114 25 144 51
<< polycont >>
rect 64 1004 98 1038
<< locali >>
rect 0 2102 368 2136
rect 62 1973 96 2102
rect 266 2031 300 2102
rect 62 1923 96 1939
rect 162 1973 196 1989
rect 266 1981 300 1997
rect 64 1038 98 1054
rect 64 988 98 1004
rect 162 1038 196 1939
rect 162 1004 213 1038
rect 62 104 96 120
rect 62 17 96 70
rect 162 104 196 1004
rect 162 54 196 70
rect 266 109 300 125
rect 266 17 300 75
rect 0 -17 368 17
<< labels >>
rlabel locali s 81 1021 81 1021 4 A
port 1 nsew
rlabel locali s 196 1021 196 1021 4 Z
port 2 nsew
rlabel locali s 184 0 184 0 4 gnd
port 3 nsew
rlabel locali s 184 2119 184 2119 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 368 1872
<< end >>
