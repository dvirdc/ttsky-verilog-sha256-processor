VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO sky130_rom_krom
   CLASS BLOCK ;
   SIZE 302.89 BY 61.28 ;
   SYMMETRY X Y R90 ;
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met1 ;
         RECT  -6.975 14.57 -6.715 14.83 ;
      END
   END clk0
   PIN cs0
      DIRECTION INPUT ;
      PORT
         LAYER met1 ;
         RECT  2.245 9.535 2.505 9.795 ;
      END
   END cs0
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met1 ;
         RECT  24.13 7.905 24.39 8.165 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met1 ;
         RECT  26.17 7.905 26.43 8.165 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met1 ;
         RECT  28.21 7.905 28.47 8.165 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met1 ;
         RECT  1.64 35.25 1.9 35.51 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met1 ;
         RECT  3.68 35.25 3.94 35.51 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met1 ;
         RECT  5.72 35.25 5.98 35.51 ;
      END
   END addr0[5]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  73.415 -0.045 73.675 0.215 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  74.955 -0.045 75.215 0.215 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  76.495 -0.045 76.755 0.215 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  78.035 -0.045 78.295 0.215 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  79.575 -0.045 79.835 0.215 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  81.115 -0.045 81.375 0.215 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  82.655 -0.045 82.915 0.215 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  84.195 -0.045 84.455 0.215 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  85.735 -0.045 85.995 0.215 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  87.275 -0.045 87.535 0.215 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  88.815 -0.045 89.075 0.215 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  90.355 -0.045 90.615 0.215 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  91.895 -0.045 92.155 0.215 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  93.435 -0.045 93.695 0.215 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  94.975 -0.045 95.235 0.215 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  96.515 -0.045 96.775 0.215 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  98.055 -0.045 98.315 0.215 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  99.595 -0.045 99.855 0.215 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  101.135 -0.045 101.395 0.215 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  102.675 -0.045 102.935 0.215 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  104.215 -0.045 104.475 0.215 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  105.755 -0.045 106.015 0.215 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  107.295 -0.045 107.555 0.215 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  108.835 -0.045 109.095 0.215 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  110.375 -0.045 110.635 0.215 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  111.915 -0.045 112.175 0.215 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  113.455 -0.045 113.715 0.215 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  114.995 -0.045 115.255 0.215 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  116.535 -0.045 116.795 0.215 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  118.075 -0.045 118.335 0.215 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  119.615 -0.045 119.875 0.215 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met1 ;
         RECT  121.155 -0.045 121.415 0.215 ;
      END
   END dout0[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  -7.48 67.02 310.37 68.76 ;
         LAYER met4 ;
         RECT  -7.48 -7.48 -5.74 68.76 ;
         LAYER met4 ;
         RECT  308.63 -7.48 310.37 68.76 ;
         LAYER met3 ;
         RECT  -7.48 -7.48 310.37 -5.74 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  -4.0 63.54 306.89 65.28 ;
         LAYER met3 ;
         RECT  -4.0 -4.0 306.89 -2.26 ;
         LAYER met4 ;
         RECT  305.15 -4.0 306.89 65.28 ;
         LAYER met4 ;
         RECT  -4.0 -4.0 -2.26 65.28 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 1.965 9.255 ;
      RECT  0.62 9.255 1.965 10.075 ;
      RECT  1.965 0.62 2.785 9.255 ;
      RECT  2.785 9.255 302.27 10.075 ;
      RECT  2.785 0.62 23.85 7.625 ;
      RECT  2.785 7.625 23.85 8.445 ;
      RECT  2.785 8.445 23.85 9.255 ;
      RECT  23.85 0.62 24.67 7.625 ;
      RECT  23.85 8.445 24.67 9.255 ;
      RECT  24.67 0.62 302.27 7.625 ;
      RECT  24.67 8.445 302.27 9.255 ;
      RECT  24.67 7.625 25.89 8.445 ;
      RECT  26.71 7.625 27.93 8.445 ;
      RECT  28.75 7.625 302.27 8.445 ;
      RECT  0.62 10.075 1.36 34.97 ;
      RECT  0.62 34.97 1.36 35.79 ;
      RECT  0.62 35.79 1.36 60.66 ;
      RECT  1.36 10.075 1.965 34.97 ;
      RECT  1.36 35.79 1.965 60.66 ;
      RECT  1.965 10.075 2.18 34.97 ;
      RECT  1.965 35.79 2.18 60.66 ;
      RECT  2.18 10.075 2.785 34.97 ;
      RECT  2.18 34.97 2.785 35.79 ;
      RECT  2.18 35.79 2.785 60.66 ;
      RECT  2.785 10.075 3.4 34.97 ;
      RECT  2.785 34.97 3.4 35.79 ;
      RECT  2.785 35.79 3.4 60.66 ;
      RECT  3.4 10.075 4.22 34.97 ;
      RECT  3.4 35.79 4.22 60.66 ;
      RECT  4.22 10.075 302.27 34.97 ;
      RECT  4.22 35.79 302.27 60.66 ;
      RECT  4.22 34.97 5.44 35.79 ;
      RECT  6.26 34.97 302.27 35.79 ;
   LAYER  met2 ;
      RECT  0.62 0.62 302.27 60.66 ;
   LAYER  met3 ;
      RECT  0.62 0.62 302.27 60.66 ;
   LAYER  met4 ;
      RECT  0.62 0.62 302.27 60.66 ;
   END
END    sky130_rom_krom
END    LIBRARY
