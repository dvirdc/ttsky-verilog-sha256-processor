magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1266 -1344 10781 4796
<< poly >>
rect 0 3388 66 3404
rect 0 3354 16 3388
rect 50 3386 66 3388
rect 1736 3388 1802 3404
rect 1736 3386 1752 3388
rect 50 3356 1752 3386
rect 50 3354 66 3356
rect 0 3338 66 3354
rect 1736 3354 1752 3356
rect 1786 3386 1802 3388
rect 3472 3388 3538 3404
rect 3472 3386 3488 3388
rect 1786 3356 3488 3386
rect 1786 3354 1802 3356
rect 1736 3338 1802 3354
rect 3472 3354 3488 3356
rect 3522 3386 3538 3388
rect 5208 3388 5274 3404
rect 5208 3386 5224 3388
rect 3522 3356 5224 3386
rect 3522 3354 3538 3356
rect 3472 3338 3538 3354
rect 5208 3354 5224 3356
rect 5258 3386 5274 3388
rect 6944 3388 7010 3404
rect 6944 3386 6960 3388
rect 5258 3356 6960 3386
rect 5258 3354 5274 3356
rect 5208 3338 5274 3354
rect 6944 3354 6960 3356
rect 6994 3386 7010 3388
rect 8680 3388 8746 3404
rect 8680 3386 8696 3388
rect 6994 3356 8696 3386
rect 6994 3354 7010 3356
rect 6944 3338 7010 3354
rect 8680 3354 8696 3356
rect 8730 3386 8746 3388
rect 9192 3388 9258 3404
rect 9192 3386 9208 3388
rect 8730 3356 9208 3386
rect 8730 3354 8746 3356
rect 8680 3338 8746 3354
rect 9192 3354 9208 3356
rect 9242 3354 9258 3388
rect 9192 3338 9258 3354
rect 0 3184 66 3200
rect 0 3150 16 3184
rect 50 3182 66 3184
rect 1736 3184 1802 3200
rect 1736 3182 1752 3184
rect 50 3152 1752 3182
rect 50 3150 66 3152
rect 0 3134 66 3150
rect 1736 3150 1752 3152
rect 1786 3182 1802 3184
rect 3472 3184 3538 3200
rect 3472 3182 3488 3184
rect 1786 3152 3488 3182
rect 1786 3150 1802 3152
rect 1736 3134 1802 3150
rect 3472 3150 3488 3152
rect 3522 3182 3538 3184
rect 5208 3184 5274 3200
rect 5208 3182 5224 3184
rect 3522 3152 5224 3182
rect 3522 3150 3538 3152
rect 3472 3134 3538 3150
rect 5208 3150 5224 3152
rect 5258 3182 5274 3184
rect 6944 3184 7010 3200
rect 6944 3182 6960 3184
rect 5258 3152 6960 3182
rect 5258 3150 5274 3152
rect 5208 3134 5274 3150
rect 6944 3150 6960 3152
rect 6994 3182 7010 3184
rect 8680 3184 8746 3200
rect 8680 3182 8696 3184
rect 6994 3152 8696 3182
rect 6994 3150 7010 3152
rect 6944 3134 7010 3150
rect 8680 3150 8696 3152
rect 8730 3182 8746 3184
rect 9192 3184 9258 3200
rect 9192 3182 9208 3184
rect 8730 3152 9208 3182
rect 8730 3150 8746 3152
rect 8680 3134 8746 3150
rect 9192 3150 9208 3152
rect 9242 3150 9258 3184
rect 9192 3134 9258 3150
rect 0 2980 66 2996
rect 0 2946 16 2980
rect 50 2978 66 2980
rect 1736 2980 1802 2996
rect 1736 2978 1752 2980
rect 50 2948 1752 2978
rect 50 2946 66 2948
rect 0 2930 66 2946
rect 1736 2946 1752 2948
rect 1786 2978 1802 2980
rect 3472 2980 3538 2996
rect 3472 2978 3488 2980
rect 1786 2948 3488 2978
rect 1786 2946 1802 2948
rect 1736 2930 1802 2946
rect 3472 2946 3488 2948
rect 3522 2978 3538 2980
rect 5208 2980 5274 2996
rect 5208 2978 5224 2980
rect 3522 2948 5224 2978
rect 3522 2946 3538 2948
rect 3472 2930 3538 2946
rect 5208 2946 5224 2948
rect 5258 2978 5274 2980
rect 6944 2980 7010 2996
rect 6944 2978 6960 2980
rect 5258 2948 6960 2978
rect 5258 2946 5274 2948
rect 5208 2930 5274 2946
rect 6944 2946 6960 2948
rect 6994 2978 7010 2980
rect 8680 2980 8746 2996
rect 8680 2978 8696 2980
rect 6994 2948 8696 2978
rect 6994 2946 7010 2948
rect 6944 2930 7010 2946
rect 8680 2946 8696 2948
rect 8730 2978 8746 2980
rect 9192 2980 9258 2996
rect 9192 2978 9208 2980
rect 8730 2948 9208 2978
rect 8730 2946 8746 2948
rect 8680 2930 8746 2946
rect 9192 2946 9208 2948
rect 9242 2946 9258 2980
rect 9192 2930 9258 2946
rect 0 2776 66 2792
rect 0 2742 16 2776
rect 50 2774 66 2776
rect 1736 2776 1802 2792
rect 1736 2774 1752 2776
rect 50 2744 1752 2774
rect 50 2742 66 2744
rect 0 2726 66 2742
rect 1736 2742 1752 2744
rect 1786 2774 1802 2776
rect 3472 2776 3538 2792
rect 3472 2774 3488 2776
rect 1786 2744 3488 2774
rect 1786 2742 1802 2744
rect 1736 2726 1802 2742
rect 3472 2742 3488 2744
rect 3522 2774 3538 2776
rect 5208 2776 5274 2792
rect 5208 2774 5224 2776
rect 3522 2744 5224 2774
rect 3522 2742 3538 2744
rect 3472 2726 3538 2742
rect 5208 2742 5224 2744
rect 5258 2774 5274 2776
rect 6944 2776 7010 2792
rect 6944 2774 6960 2776
rect 5258 2744 6960 2774
rect 5258 2742 5274 2744
rect 5208 2726 5274 2742
rect 6944 2742 6960 2744
rect 6994 2774 7010 2776
rect 8680 2776 8746 2792
rect 8680 2774 8696 2776
rect 6994 2744 8696 2774
rect 6994 2742 7010 2744
rect 6944 2726 7010 2742
rect 8680 2742 8696 2744
rect 8730 2774 8746 2776
rect 9192 2776 9258 2792
rect 9192 2774 9208 2776
rect 8730 2744 9208 2774
rect 8730 2742 8746 2744
rect 8680 2726 8746 2742
rect 9192 2742 9208 2744
rect 9242 2742 9258 2776
rect 9192 2726 9258 2742
rect 0 2572 66 2588
rect 0 2538 16 2572
rect 50 2570 66 2572
rect 1736 2572 1802 2588
rect 1736 2570 1752 2572
rect 50 2540 1752 2570
rect 50 2538 66 2540
rect 0 2522 66 2538
rect 1736 2538 1752 2540
rect 1786 2570 1802 2572
rect 3472 2572 3538 2588
rect 3472 2570 3488 2572
rect 1786 2540 3488 2570
rect 1786 2538 1802 2540
rect 1736 2522 1802 2538
rect 3472 2538 3488 2540
rect 3522 2570 3538 2572
rect 5208 2572 5274 2588
rect 5208 2570 5224 2572
rect 3522 2540 5224 2570
rect 3522 2538 3538 2540
rect 3472 2522 3538 2538
rect 5208 2538 5224 2540
rect 5258 2570 5274 2572
rect 6944 2572 7010 2588
rect 6944 2570 6960 2572
rect 5258 2540 6960 2570
rect 5258 2538 5274 2540
rect 5208 2522 5274 2538
rect 6944 2538 6960 2540
rect 6994 2570 7010 2572
rect 8680 2572 8746 2588
rect 8680 2570 8696 2572
rect 6994 2540 8696 2570
rect 6994 2538 7010 2540
rect 6944 2522 7010 2538
rect 8680 2538 8696 2540
rect 8730 2570 8746 2572
rect 9192 2572 9258 2588
rect 9192 2570 9208 2572
rect 8730 2540 9208 2570
rect 8730 2538 8746 2540
rect 8680 2522 8746 2538
rect 9192 2538 9208 2540
rect 9242 2538 9258 2572
rect 9192 2522 9258 2538
rect 0 2368 66 2384
rect 0 2334 16 2368
rect 50 2366 66 2368
rect 1736 2368 1802 2384
rect 1736 2366 1752 2368
rect 50 2336 1752 2366
rect 50 2334 66 2336
rect 0 2318 66 2334
rect 1736 2334 1752 2336
rect 1786 2366 1802 2368
rect 3472 2368 3538 2384
rect 3472 2366 3488 2368
rect 1786 2336 3488 2366
rect 1786 2334 1802 2336
rect 1736 2318 1802 2334
rect 3472 2334 3488 2336
rect 3522 2366 3538 2368
rect 5208 2368 5274 2384
rect 5208 2366 5224 2368
rect 3522 2336 5224 2366
rect 3522 2334 3538 2336
rect 3472 2318 3538 2334
rect 5208 2334 5224 2336
rect 5258 2366 5274 2368
rect 6944 2368 7010 2384
rect 6944 2366 6960 2368
rect 5258 2336 6960 2366
rect 5258 2334 5274 2336
rect 5208 2318 5274 2334
rect 6944 2334 6960 2336
rect 6994 2366 7010 2368
rect 8680 2368 8746 2384
rect 8680 2366 8696 2368
rect 6994 2336 8696 2366
rect 6994 2334 7010 2336
rect 6944 2318 7010 2334
rect 8680 2334 8696 2336
rect 8730 2366 8746 2368
rect 9192 2368 9258 2384
rect 9192 2366 9208 2368
rect 8730 2336 9208 2366
rect 8730 2334 8746 2336
rect 8680 2318 8746 2334
rect 9192 2334 9208 2336
rect 9242 2334 9258 2368
rect 9192 2318 9258 2334
rect 0 2164 66 2180
rect 0 2130 16 2164
rect 50 2162 66 2164
rect 1736 2164 1802 2180
rect 1736 2162 1752 2164
rect 50 2132 1752 2162
rect 50 2130 66 2132
rect 0 2114 66 2130
rect 1736 2130 1752 2132
rect 1786 2162 1802 2164
rect 3472 2164 3538 2180
rect 3472 2162 3488 2164
rect 1786 2132 3488 2162
rect 1786 2130 1802 2132
rect 1736 2114 1802 2130
rect 3472 2130 3488 2132
rect 3522 2162 3538 2164
rect 5208 2164 5274 2180
rect 5208 2162 5224 2164
rect 3522 2132 5224 2162
rect 3522 2130 3538 2132
rect 3472 2114 3538 2130
rect 5208 2130 5224 2132
rect 5258 2162 5274 2164
rect 6944 2164 7010 2180
rect 6944 2162 6960 2164
rect 5258 2132 6960 2162
rect 5258 2130 5274 2132
rect 5208 2114 5274 2130
rect 6944 2130 6960 2132
rect 6994 2162 7010 2164
rect 8680 2164 8746 2180
rect 8680 2162 8696 2164
rect 6994 2132 8696 2162
rect 6994 2130 7010 2132
rect 6944 2114 7010 2130
rect 8680 2130 8696 2132
rect 8730 2162 8746 2164
rect 9192 2164 9258 2180
rect 9192 2162 9208 2164
rect 8730 2132 9208 2162
rect 8730 2130 8746 2132
rect 8680 2114 8746 2130
rect 9192 2130 9208 2132
rect 9242 2130 9258 2164
rect 9192 2114 9258 2130
rect 0 1960 66 1976
rect 0 1926 16 1960
rect 50 1958 66 1960
rect 1736 1960 1802 1976
rect 1736 1958 1752 1960
rect 50 1928 1752 1958
rect 50 1926 66 1928
rect 0 1910 66 1926
rect 1736 1926 1752 1928
rect 1786 1958 1802 1960
rect 3472 1960 3538 1976
rect 3472 1958 3488 1960
rect 1786 1928 3488 1958
rect 1786 1926 1802 1928
rect 1736 1910 1802 1926
rect 3472 1926 3488 1928
rect 3522 1958 3538 1960
rect 5208 1960 5274 1976
rect 5208 1958 5224 1960
rect 3522 1928 5224 1958
rect 3522 1926 3538 1928
rect 3472 1910 3538 1926
rect 5208 1926 5224 1928
rect 5258 1958 5274 1960
rect 6944 1960 7010 1976
rect 6944 1958 6960 1960
rect 5258 1928 6960 1958
rect 5258 1926 5274 1928
rect 5208 1910 5274 1926
rect 6944 1926 6960 1928
rect 6994 1958 7010 1960
rect 8680 1960 8746 1976
rect 8680 1958 8696 1960
rect 6994 1928 8696 1958
rect 6994 1926 7010 1928
rect 6944 1910 7010 1926
rect 8680 1926 8696 1928
rect 8730 1958 8746 1960
rect 9192 1960 9258 1976
rect 9192 1958 9208 1960
rect 8730 1928 9208 1958
rect 8730 1926 8746 1928
rect 8680 1910 8746 1926
rect 9192 1926 9208 1928
rect 9242 1926 9258 1960
rect 9192 1910 9258 1926
rect 0 1756 66 1772
rect 0 1722 16 1756
rect 50 1754 66 1756
rect 1736 1756 1802 1772
rect 1736 1754 1752 1756
rect 50 1724 1752 1754
rect 50 1722 66 1724
rect 0 1706 66 1722
rect 1736 1722 1752 1724
rect 1786 1754 1802 1756
rect 3472 1756 3538 1772
rect 3472 1754 3488 1756
rect 1786 1724 3488 1754
rect 1786 1722 1802 1724
rect 1736 1706 1802 1722
rect 3472 1722 3488 1724
rect 3522 1754 3538 1756
rect 5208 1756 5274 1772
rect 5208 1754 5224 1756
rect 3522 1724 5224 1754
rect 3522 1722 3538 1724
rect 3472 1706 3538 1722
rect 5208 1722 5224 1724
rect 5258 1754 5274 1756
rect 6944 1756 7010 1772
rect 6944 1754 6960 1756
rect 5258 1724 6960 1754
rect 5258 1722 5274 1724
rect 5208 1706 5274 1722
rect 6944 1722 6960 1724
rect 6994 1754 7010 1756
rect 8680 1756 8746 1772
rect 8680 1754 8696 1756
rect 6994 1724 8696 1754
rect 6994 1722 7010 1724
rect 6944 1706 7010 1722
rect 8680 1722 8696 1724
rect 8730 1754 8746 1756
rect 9192 1756 9258 1772
rect 9192 1754 9208 1756
rect 8730 1724 9208 1754
rect 8730 1722 8746 1724
rect 8680 1706 8746 1722
rect 9192 1722 9208 1724
rect 9242 1722 9258 1756
rect 9192 1706 9258 1722
rect 0 1552 66 1568
rect 0 1518 16 1552
rect 50 1550 66 1552
rect 1736 1552 1802 1568
rect 1736 1550 1752 1552
rect 50 1520 1752 1550
rect 50 1518 66 1520
rect 0 1502 66 1518
rect 1736 1518 1752 1520
rect 1786 1550 1802 1552
rect 3472 1552 3538 1568
rect 3472 1550 3488 1552
rect 1786 1520 3488 1550
rect 1786 1518 1802 1520
rect 1736 1502 1802 1518
rect 3472 1518 3488 1520
rect 3522 1550 3538 1552
rect 5208 1552 5274 1568
rect 5208 1550 5224 1552
rect 3522 1520 5224 1550
rect 3522 1518 3538 1520
rect 3472 1502 3538 1518
rect 5208 1518 5224 1520
rect 5258 1550 5274 1552
rect 6944 1552 7010 1568
rect 6944 1550 6960 1552
rect 5258 1520 6960 1550
rect 5258 1518 5274 1520
rect 5208 1502 5274 1518
rect 6944 1518 6960 1520
rect 6994 1550 7010 1552
rect 8680 1552 8746 1568
rect 8680 1550 8696 1552
rect 6994 1520 8696 1550
rect 6994 1518 7010 1520
rect 6944 1502 7010 1518
rect 8680 1518 8696 1520
rect 8730 1550 8746 1552
rect 9192 1552 9258 1568
rect 9192 1550 9208 1552
rect 8730 1520 9208 1550
rect 8730 1518 8746 1520
rect 8680 1502 8746 1518
rect 9192 1518 9208 1520
rect 9242 1518 9258 1552
rect 9192 1502 9258 1518
rect 0 1348 66 1364
rect 0 1314 16 1348
rect 50 1346 66 1348
rect 1736 1348 1802 1364
rect 1736 1346 1752 1348
rect 50 1316 1752 1346
rect 50 1314 66 1316
rect 0 1298 66 1314
rect 1736 1314 1752 1316
rect 1786 1346 1802 1348
rect 3472 1348 3538 1364
rect 3472 1346 3488 1348
rect 1786 1316 3488 1346
rect 1786 1314 1802 1316
rect 1736 1298 1802 1314
rect 3472 1314 3488 1316
rect 3522 1346 3538 1348
rect 5208 1348 5274 1364
rect 5208 1346 5224 1348
rect 3522 1316 5224 1346
rect 3522 1314 3538 1316
rect 3472 1298 3538 1314
rect 5208 1314 5224 1316
rect 5258 1346 5274 1348
rect 6944 1348 7010 1364
rect 6944 1346 6960 1348
rect 5258 1316 6960 1346
rect 5258 1314 5274 1316
rect 5208 1298 5274 1314
rect 6944 1314 6960 1316
rect 6994 1346 7010 1348
rect 8680 1348 8746 1364
rect 8680 1346 8696 1348
rect 6994 1316 8696 1346
rect 6994 1314 7010 1316
rect 6944 1298 7010 1314
rect 8680 1314 8696 1316
rect 8730 1346 8746 1348
rect 9192 1348 9258 1364
rect 9192 1346 9208 1348
rect 8730 1316 9208 1346
rect 8730 1314 8746 1316
rect 8680 1298 8746 1314
rect 9192 1314 9208 1316
rect 9242 1314 9258 1348
rect 9192 1298 9258 1314
rect 0 1144 66 1160
rect 0 1110 16 1144
rect 50 1142 66 1144
rect 1736 1144 1802 1160
rect 1736 1142 1752 1144
rect 50 1112 1752 1142
rect 50 1110 66 1112
rect 0 1094 66 1110
rect 1736 1110 1752 1112
rect 1786 1142 1802 1144
rect 3472 1144 3538 1160
rect 3472 1142 3488 1144
rect 1786 1112 3488 1142
rect 1786 1110 1802 1112
rect 1736 1094 1802 1110
rect 3472 1110 3488 1112
rect 3522 1142 3538 1144
rect 5208 1144 5274 1160
rect 5208 1142 5224 1144
rect 3522 1112 5224 1142
rect 3522 1110 3538 1112
rect 3472 1094 3538 1110
rect 5208 1110 5224 1112
rect 5258 1142 5274 1144
rect 6944 1144 7010 1160
rect 6944 1142 6960 1144
rect 5258 1112 6960 1142
rect 5258 1110 5274 1112
rect 5208 1094 5274 1110
rect 6944 1110 6960 1112
rect 6994 1142 7010 1144
rect 8680 1144 8746 1160
rect 8680 1142 8696 1144
rect 6994 1112 8696 1142
rect 6994 1110 7010 1112
rect 6944 1094 7010 1110
rect 8680 1110 8696 1112
rect 8730 1142 8746 1144
rect 9192 1144 9258 1160
rect 9192 1142 9208 1144
rect 8730 1112 9208 1142
rect 8730 1110 8746 1112
rect 8680 1094 8746 1110
rect 9192 1110 9208 1112
rect 9242 1110 9258 1144
rect 9192 1094 9258 1110
rect 0 940 66 956
rect 0 906 16 940
rect 50 938 66 940
rect 1736 940 1802 956
rect 1736 938 1752 940
rect 50 908 1752 938
rect 50 906 66 908
rect 0 890 66 906
rect 1736 906 1752 908
rect 1786 938 1802 940
rect 3472 940 3538 956
rect 3472 938 3488 940
rect 1786 908 3488 938
rect 1786 906 1802 908
rect 1736 890 1802 906
rect 3472 906 3488 908
rect 3522 938 3538 940
rect 5208 940 5274 956
rect 5208 938 5224 940
rect 3522 908 5224 938
rect 3522 906 3538 908
rect 3472 890 3538 906
rect 5208 906 5224 908
rect 5258 938 5274 940
rect 6944 940 7010 956
rect 6944 938 6960 940
rect 5258 908 6960 938
rect 5258 906 5274 908
rect 5208 890 5274 906
rect 6944 906 6960 908
rect 6994 938 7010 940
rect 8680 940 8746 956
rect 8680 938 8696 940
rect 6994 908 8696 938
rect 6994 906 7010 908
rect 6944 890 7010 906
rect 8680 906 8696 908
rect 8730 938 8746 940
rect 9192 940 9258 956
rect 9192 938 9208 940
rect 8730 908 9208 938
rect 8730 906 8746 908
rect 8680 890 8746 906
rect 9192 906 9208 908
rect 9242 906 9258 940
rect 9192 890 9258 906
<< polycont >>
rect 16 3354 50 3388
rect 1752 3354 1786 3388
rect 3488 3354 3522 3388
rect 5224 3354 5258 3388
rect 6960 3354 6994 3388
rect 8696 3354 8730 3388
rect 9208 3354 9242 3388
rect 16 3150 50 3184
rect 1752 3150 1786 3184
rect 3488 3150 3522 3184
rect 5224 3150 5258 3184
rect 6960 3150 6994 3184
rect 8696 3150 8730 3184
rect 9208 3150 9242 3184
rect 16 2946 50 2980
rect 1752 2946 1786 2980
rect 3488 2946 3522 2980
rect 5224 2946 5258 2980
rect 6960 2946 6994 2980
rect 8696 2946 8730 2980
rect 9208 2946 9242 2980
rect 16 2742 50 2776
rect 1752 2742 1786 2776
rect 3488 2742 3522 2776
rect 5224 2742 5258 2776
rect 6960 2742 6994 2776
rect 8696 2742 8730 2776
rect 9208 2742 9242 2776
rect 16 2538 50 2572
rect 1752 2538 1786 2572
rect 3488 2538 3522 2572
rect 5224 2538 5258 2572
rect 6960 2538 6994 2572
rect 8696 2538 8730 2572
rect 9208 2538 9242 2572
rect 16 2334 50 2368
rect 1752 2334 1786 2368
rect 3488 2334 3522 2368
rect 5224 2334 5258 2368
rect 6960 2334 6994 2368
rect 8696 2334 8730 2368
rect 9208 2334 9242 2368
rect 16 2130 50 2164
rect 1752 2130 1786 2164
rect 3488 2130 3522 2164
rect 5224 2130 5258 2164
rect 6960 2130 6994 2164
rect 8696 2130 8730 2164
rect 9208 2130 9242 2164
rect 16 1926 50 1960
rect 1752 1926 1786 1960
rect 3488 1926 3522 1960
rect 5224 1926 5258 1960
rect 6960 1926 6994 1960
rect 8696 1926 8730 1960
rect 9208 1926 9242 1960
rect 16 1722 50 1756
rect 1752 1722 1786 1756
rect 3488 1722 3522 1756
rect 5224 1722 5258 1756
rect 6960 1722 6994 1756
rect 8696 1722 8730 1756
rect 9208 1722 9242 1756
rect 16 1518 50 1552
rect 1752 1518 1786 1552
rect 3488 1518 3522 1552
rect 5224 1518 5258 1552
rect 6960 1518 6994 1552
rect 8696 1518 8730 1552
rect 9208 1518 9242 1552
rect 16 1314 50 1348
rect 1752 1314 1786 1348
rect 3488 1314 3522 1348
rect 5224 1314 5258 1348
rect 6960 1314 6994 1348
rect 8696 1314 8730 1348
rect 9208 1314 9242 1348
rect 16 1110 50 1144
rect 1752 1110 1786 1144
rect 3488 1110 3522 1144
rect 5224 1110 5258 1144
rect 6960 1110 6994 1144
rect 8696 1110 8730 1144
rect 9208 1110 9242 1144
rect 16 906 50 940
rect 1752 906 1786 940
rect 3488 906 3522 940
rect 5224 906 5258 940
rect 6960 906 6994 940
rect 8696 906 8730 940
rect 9208 906 9242 940
<< locali >>
rect 16 3388 50 3404
rect 16 3338 50 3354
rect 1752 3388 1786 3404
rect 1752 3338 1786 3354
rect 3488 3388 3522 3404
rect 3488 3338 3522 3354
rect 5224 3388 5258 3404
rect 5224 3338 5258 3354
rect 6960 3388 6994 3404
rect 6960 3338 6994 3354
rect 8696 3388 8730 3404
rect 8696 3338 8730 3354
rect 9208 3388 9242 3404
rect 9208 3338 9242 3354
rect 28 3252 44 3286
rect 78 3252 94 3286
rect 1764 3252 1780 3286
rect 1814 3252 1830 3286
rect 3500 3252 3516 3286
rect 3550 3252 3566 3286
rect 5236 3252 5252 3286
rect 5286 3252 5302 3286
rect 6972 3252 6988 3286
rect 7022 3252 7038 3286
rect 8708 3252 8724 3286
rect 8758 3252 8774 3286
rect 9220 3252 9236 3286
rect 9270 3252 9286 3286
rect 16 3184 50 3200
rect 16 3134 50 3150
rect 1752 3184 1786 3200
rect 1752 3134 1786 3150
rect 3488 3184 3522 3200
rect 3488 3134 3522 3150
rect 5224 3184 5258 3200
rect 5224 3134 5258 3150
rect 6960 3184 6994 3200
rect 6960 3134 6994 3150
rect 8696 3184 8730 3200
rect 8696 3134 8730 3150
rect 9208 3184 9242 3200
rect 9208 3134 9242 3150
rect 28 3048 44 3082
rect 78 3048 94 3082
rect 1764 3048 1780 3082
rect 1814 3048 1830 3082
rect 3500 3048 3516 3082
rect 3550 3048 3566 3082
rect 5236 3048 5252 3082
rect 5286 3048 5302 3082
rect 6972 3048 6988 3082
rect 7022 3048 7038 3082
rect 8708 3048 8724 3082
rect 8758 3048 8774 3082
rect 9220 3048 9236 3082
rect 9270 3048 9286 3082
rect 16 2980 50 2996
rect 16 2930 50 2946
rect 1752 2980 1786 2996
rect 1752 2930 1786 2946
rect 3488 2980 3522 2996
rect 3488 2930 3522 2946
rect 5224 2980 5258 2996
rect 5224 2930 5258 2946
rect 6960 2980 6994 2996
rect 6960 2930 6994 2946
rect 8696 2980 8730 2996
rect 8696 2930 8730 2946
rect 9208 2980 9242 2996
rect 9208 2930 9242 2946
rect 28 2844 44 2878
rect 78 2844 94 2878
rect 1764 2844 1780 2878
rect 1814 2844 1830 2878
rect 3500 2844 3516 2878
rect 3550 2844 3566 2878
rect 5236 2844 5252 2878
rect 5286 2844 5302 2878
rect 6972 2844 6988 2878
rect 7022 2844 7038 2878
rect 8708 2844 8724 2878
rect 8758 2844 8774 2878
rect 9220 2844 9236 2878
rect 9270 2844 9286 2878
rect 16 2776 50 2792
rect 16 2726 50 2742
rect 1752 2776 1786 2792
rect 1752 2726 1786 2742
rect 3488 2776 3522 2792
rect 3488 2726 3522 2742
rect 5224 2776 5258 2792
rect 5224 2726 5258 2742
rect 6960 2776 6994 2792
rect 6960 2726 6994 2742
rect 8696 2776 8730 2792
rect 8696 2726 8730 2742
rect 9208 2776 9242 2792
rect 9208 2726 9242 2742
rect 28 2640 44 2674
rect 78 2640 94 2674
rect 1764 2640 1780 2674
rect 1814 2640 1830 2674
rect 3500 2640 3516 2674
rect 3550 2640 3566 2674
rect 5236 2640 5252 2674
rect 5286 2640 5302 2674
rect 6972 2640 6988 2674
rect 7022 2640 7038 2674
rect 8708 2640 8724 2674
rect 8758 2640 8774 2674
rect 9220 2640 9236 2674
rect 9270 2640 9286 2674
rect 16 2572 50 2588
rect 16 2522 50 2538
rect 1752 2572 1786 2588
rect 1752 2522 1786 2538
rect 3488 2572 3522 2588
rect 3488 2522 3522 2538
rect 5224 2572 5258 2588
rect 5224 2522 5258 2538
rect 6960 2572 6994 2588
rect 6960 2522 6994 2538
rect 8696 2572 8730 2588
rect 8696 2522 8730 2538
rect 9208 2572 9242 2588
rect 9208 2522 9242 2538
rect 28 2436 44 2470
rect 78 2436 94 2470
rect 1764 2436 1780 2470
rect 1814 2436 1830 2470
rect 3500 2436 3516 2470
rect 3550 2436 3566 2470
rect 5236 2436 5252 2470
rect 5286 2436 5302 2470
rect 6972 2436 6988 2470
rect 7022 2436 7038 2470
rect 8708 2436 8724 2470
rect 8758 2436 8774 2470
rect 9220 2436 9236 2470
rect 9270 2436 9286 2470
rect 16 2368 50 2384
rect 16 2318 50 2334
rect 1752 2368 1786 2384
rect 1752 2318 1786 2334
rect 3488 2368 3522 2384
rect 3488 2318 3522 2334
rect 5224 2368 5258 2384
rect 5224 2318 5258 2334
rect 6960 2368 6994 2384
rect 6960 2318 6994 2334
rect 8696 2368 8730 2384
rect 8696 2318 8730 2334
rect 9208 2368 9242 2384
rect 9208 2318 9242 2334
rect 28 2232 44 2266
rect 78 2232 94 2266
rect 1764 2232 1780 2266
rect 1814 2232 1830 2266
rect 3500 2232 3516 2266
rect 3550 2232 3566 2266
rect 5236 2232 5252 2266
rect 5286 2232 5302 2266
rect 6972 2232 6988 2266
rect 7022 2232 7038 2266
rect 8708 2232 8724 2266
rect 8758 2232 8774 2266
rect 9220 2232 9236 2266
rect 9270 2232 9286 2266
rect 16 2164 50 2180
rect 16 2114 50 2130
rect 1752 2164 1786 2180
rect 1752 2114 1786 2130
rect 3488 2164 3522 2180
rect 3488 2114 3522 2130
rect 5224 2164 5258 2180
rect 5224 2114 5258 2130
rect 6960 2164 6994 2180
rect 6960 2114 6994 2130
rect 8696 2164 8730 2180
rect 8696 2114 8730 2130
rect 9208 2164 9242 2180
rect 9208 2114 9242 2130
rect 28 2028 44 2062
rect 78 2028 94 2062
rect 1764 2028 1780 2062
rect 1814 2028 1830 2062
rect 3500 2028 3516 2062
rect 3550 2028 3566 2062
rect 5236 2028 5252 2062
rect 5286 2028 5302 2062
rect 6972 2028 6988 2062
rect 7022 2028 7038 2062
rect 8708 2028 8724 2062
rect 8758 2028 8774 2062
rect 9220 2028 9236 2062
rect 9270 2028 9286 2062
rect 16 1960 50 1976
rect 16 1910 50 1926
rect 1752 1960 1786 1976
rect 1752 1910 1786 1926
rect 3488 1960 3522 1976
rect 3488 1910 3522 1926
rect 5224 1960 5258 1976
rect 5224 1910 5258 1926
rect 6960 1960 6994 1976
rect 6960 1910 6994 1926
rect 8696 1960 8730 1976
rect 8696 1910 8730 1926
rect 9208 1960 9242 1976
rect 9208 1910 9242 1926
rect 28 1824 44 1858
rect 78 1824 94 1858
rect 1764 1824 1780 1858
rect 1814 1824 1830 1858
rect 3500 1824 3516 1858
rect 3550 1824 3566 1858
rect 5236 1824 5252 1858
rect 5286 1824 5302 1858
rect 6972 1824 6988 1858
rect 7022 1824 7038 1858
rect 8708 1824 8724 1858
rect 8758 1824 8774 1858
rect 9220 1824 9236 1858
rect 9270 1824 9286 1858
rect 16 1756 50 1772
rect 16 1706 50 1722
rect 1752 1756 1786 1772
rect 1752 1706 1786 1722
rect 3488 1756 3522 1772
rect 3488 1706 3522 1722
rect 5224 1756 5258 1772
rect 5224 1706 5258 1722
rect 6960 1756 6994 1772
rect 6960 1706 6994 1722
rect 8696 1756 8730 1772
rect 8696 1706 8730 1722
rect 9208 1756 9242 1772
rect 9208 1706 9242 1722
rect 28 1620 44 1654
rect 78 1620 94 1654
rect 1764 1620 1780 1654
rect 1814 1620 1830 1654
rect 3500 1620 3516 1654
rect 3550 1620 3566 1654
rect 5236 1620 5252 1654
rect 5286 1620 5302 1654
rect 6972 1620 6988 1654
rect 7022 1620 7038 1654
rect 8708 1620 8724 1654
rect 8758 1620 8774 1654
rect 9220 1620 9236 1654
rect 9270 1620 9286 1654
rect 16 1552 50 1568
rect 16 1502 50 1518
rect 1752 1552 1786 1568
rect 1752 1502 1786 1518
rect 3488 1552 3522 1568
rect 3488 1502 3522 1518
rect 5224 1552 5258 1568
rect 5224 1502 5258 1518
rect 6960 1552 6994 1568
rect 6960 1502 6994 1518
rect 8696 1552 8730 1568
rect 8696 1502 8730 1518
rect 9208 1552 9242 1568
rect 9208 1502 9242 1518
rect 28 1416 44 1450
rect 78 1416 94 1450
rect 1764 1416 1780 1450
rect 1814 1416 1830 1450
rect 3500 1416 3516 1450
rect 3550 1416 3566 1450
rect 5236 1416 5252 1450
rect 5286 1416 5302 1450
rect 6972 1416 6988 1450
rect 7022 1416 7038 1450
rect 8708 1416 8724 1450
rect 8758 1416 8774 1450
rect 9220 1416 9236 1450
rect 9270 1416 9286 1450
rect 16 1348 50 1364
rect 16 1298 50 1314
rect 1752 1348 1786 1364
rect 1752 1298 1786 1314
rect 3488 1348 3522 1364
rect 3488 1298 3522 1314
rect 5224 1348 5258 1364
rect 5224 1298 5258 1314
rect 6960 1348 6994 1364
rect 6960 1298 6994 1314
rect 8696 1348 8730 1364
rect 8696 1298 8730 1314
rect 9208 1348 9242 1364
rect 9208 1298 9242 1314
rect 28 1212 44 1246
rect 78 1212 94 1246
rect 1764 1212 1780 1246
rect 1814 1212 1830 1246
rect 3500 1212 3516 1246
rect 3550 1212 3566 1246
rect 5236 1212 5252 1246
rect 5286 1212 5302 1246
rect 6972 1212 6988 1246
rect 7022 1212 7038 1246
rect 8708 1212 8724 1246
rect 8758 1212 8774 1246
rect 9220 1212 9236 1246
rect 9270 1212 9286 1246
rect 16 1144 50 1160
rect 16 1094 50 1110
rect 1752 1144 1786 1160
rect 1752 1094 1786 1110
rect 3488 1144 3522 1160
rect 3488 1094 3522 1110
rect 5224 1144 5258 1160
rect 5224 1094 5258 1110
rect 6960 1144 6994 1160
rect 6960 1094 6994 1110
rect 8696 1144 8730 1160
rect 8696 1094 8730 1110
rect 9208 1144 9242 1160
rect 9208 1094 9242 1110
rect 28 1008 44 1042
rect 78 1008 94 1042
rect 1764 1008 1780 1042
rect 1814 1008 1830 1042
rect 3500 1008 3516 1042
rect 3550 1008 3566 1042
rect 5236 1008 5252 1042
rect 5286 1008 5302 1042
rect 6972 1008 6988 1042
rect 7022 1008 7038 1042
rect 8708 1008 8724 1042
rect 8758 1008 8774 1042
rect 9220 1008 9236 1042
rect 9270 1008 9286 1042
rect 16 940 50 956
rect 16 890 50 906
rect 1752 940 1786 956
rect 1752 890 1786 906
rect 3488 940 3522 956
rect 3488 890 3522 906
rect 5224 940 5258 956
rect 5224 890 5258 906
rect 6960 940 6994 956
rect 6960 890 6994 906
rect 8696 940 8730 956
rect 8696 890 8730 906
rect 9208 940 9242 956
rect 9208 890 9242 906
<< viali >>
rect 16 3354 50 3388
rect 1752 3354 1786 3388
rect 3488 3354 3522 3388
rect 5224 3354 5258 3388
rect 6960 3354 6994 3388
rect 8696 3354 8730 3388
rect 9208 3354 9242 3388
rect 44 3252 78 3286
rect 1780 3252 1814 3286
rect 3516 3252 3550 3286
rect 5252 3252 5286 3286
rect 6988 3252 7022 3286
rect 8724 3252 8758 3286
rect 9236 3252 9270 3286
rect 16 3150 50 3184
rect 1752 3150 1786 3184
rect 3488 3150 3522 3184
rect 5224 3150 5258 3184
rect 6960 3150 6994 3184
rect 8696 3150 8730 3184
rect 9208 3150 9242 3184
rect 44 3048 78 3082
rect 1780 3048 1814 3082
rect 3516 3048 3550 3082
rect 5252 3048 5286 3082
rect 6988 3048 7022 3082
rect 8724 3048 8758 3082
rect 9236 3048 9270 3082
rect 16 2946 50 2980
rect 1752 2946 1786 2980
rect 3488 2946 3522 2980
rect 5224 2946 5258 2980
rect 6960 2946 6994 2980
rect 8696 2946 8730 2980
rect 9208 2946 9242 2980
rect 44 2844 78 2878
rect 1780 2844 1814 2878
rect 3516 2844 3550 2878
rect 5252 2844 5286 2878
rect 6988 2844 7022 2878
rect 8724 2844 8758 2878
rect 9236 2844 9270 2878
rect 16 2742 50 2776
rect 1752 2742 1786 2776
rect 3488 2742 3522 2776
rect 5224 2742 5258 2776
rect 6960 2742 6994 2776
rect 8696 2742 8730 2776
rect 9208 2742 9242 2776
rect 44 2640 78 2674
rect 1780 2640 1814 2674
rect 3516 2640 3550 2674
rect 5252 2640 5286 2674
rect 6988 2640 7022 2674
rect 8724 2640 8758 2674
rect 9236 2640 9270 2674
rect 16 2538 50 2572
rect 1752 2538 1786 2572
rect 3488 2538 3522 2572
rect 5224 2538 5258 2572
rect 6960 2538 6994 2572
rect 8696 2538 8730 2572
rect 9208 2538 9242 2572
rect 44 2436 78 2470
rect 1780 2436 1814 2470
rect 3516 2436 3550 2470
rect 5252 2436 5286 2470
rect 6988 2436 7022 2470
rect 8724 2436 8758 2470
rect 9236 2436 9270 2470
rect 16 2334 50 2368
rect 1752 2334 1786 2368
rect 3488 2334 3522 2368
rect 5224 2334 5258 2368
rect 6960 2334 6994 2368
rect 8696 2334 8730 2368
rect 9208 2334 9242 2368
rect 44 2232 78 2266
rect 1780 2232 1814 2266
rect 3516 2232 3550 2266
rect 5252 2232 5286 2266
rect 6988 2232 7022 2266
rect 8724 2232 8758 2266
rect 9236 2232 9270 2266
rect 16 2130 50 2164
rect 1752 2130 1786 2164
rect 3488 2130 3522 2164
rect 5224 2130 5258 2164
rect 6960 2130 6994 2164
rect 8696 2130 8730 2164
rect 9208 2130 9242 2164
rect 44 2028 78 2062
rect 1780 2028 1814 2062
rect 3516 2028 3550 2062
rect 5252 2028 5286 2062
rect 6988 2028 7022 2062
rect 8724 2028 8758 2062
rect 9236 2028 9270 2062
rect 16 1926 50 1960
rect 1752 1926 1786 1960
rect 3488 1926 3522 1960
rect 5224 1926 5258 1960
rect 6960 1926 6994 1960
rect 8696 1926 8730 1960
rect 9208 1926 9242 1960
rect 44 1824 78 1858
rect 1780 1824 1814 1858
rect 3516 1824 3550 1858
rect 5252 1824 5286 1858
rect 6988 1824 7022 1858
rect 8724 1824 8758 1858
rect 9236 1824 9270 1858
rect 16 1722 50 1756
rect 1752 1722 1786 1756
rect 3488 1722 3522 1756
rect 5224 1722 5258 1756
rect 6960 1722 6994 1756
rect 8696 1722 8730 1756
rect 9208 1722 9242 1756
rect 44 1620 78 1654
rect 1780 1620 1814 1654
rect 3516 1620 3550 1654
rect 5252 1620 5286 1654
rect 6988 1620 7022 1654
rect 8724 1620 8758 1654
rect 9236 1620 9270 1654
rect 16 1518 50 1552
rect 1752 1518 1786 1552
rect 3488 1518 3522 1552
rect 5224 1518 5258 1552
rect 6960 1518 6994 1552
rect 8696 1518 8730 1552
rect 9208 1518 9242 1552
rect 44 1416 78 1450
rect 1780 1416 1814 1450
rect 3516 1416 3550 1450
rect 5252 1416 5286 1450
rect 6988 1416 7022 1450
rect 8724 1416 8758 1450
rect 9236 1416 9270 1450
rect 16 1314 50 1348
rect 1752 1314 1786 1348
rect 3488 1314 3522 1348
rect 5224 1314 5258 1348
rect 6960 1314 6994 1348
rect 8696 1314 8730 1348
rect 9208 1314 9242 1348
rect 44 1212 78 1246
rect 1780 1212 1814 1246
rect 3516 1212 3550 1246
rect 5252 1212 5286 1246
rect 6988 1212 7022 1246
rect 8724 1212 8758 1246
rect 9236 1212 9270 1246
rect 16 1110 50 1144
rect 1752 1110 1786 1144
rect 3488 1110 3522 1144
rect 5224 1110 5258 1144
rect 6960 1110 6994 1144
rect 8696 1110 8730 1144
rect 9208 1110 9242 1144
rect 44 1008 78 1042
rect 1780 1008 1814 1042
rect 3516 1008 3550 1042
rect 5252 1008 5286 1042
rect 6988 1008 7022 1042
rect 8724 1008 8758 1042
rect 9236 1008 9270 1042
rect 16 906 50 940
rect 1752 906 1786 940
rect 3488 906 3522 940
rect 5224 906 5258 940
rect 6960 906 6994 940
rect 8696 906 8730 940
rect 9208 906 9242 940
<< metal1 >>
rect 29 3472 35 3524
rect 87 3512 93 3524
rect 1765 3512 1771 3524
rect 87 3484 1771 3512
rect 87 3472 93 3484
rect 1765 3472 1771 3484
rect 1823 3512 1829 3524
rect 3501 3512 3507 3524
rect 1823 3484 3507 3512
rect 1823 3472 1829 3484
rect 3501 3472 3507 3484
rect 3559 3512 3565 3524
rect 5237 3512 5243 3524
rect 3559 3484 5243 3512
rect 3559 3472 3565 3484
rect 5237 3472 5243 3484
rect 5295 3512 5301 3524
rect 6973 3512 6979 3524
rect 5295 3484 6979 3512
rect 5295 3472 5301 3484
rect 6973 3472 6979 3484
rect 7031 3512 7037 3524
rect 8709 3512 8715 3524
rect 7031 3484 8715 3512
rect 7031 3472 7037 3484
rect 8709 3472 8715 3484
rect 8767 3512 8773 3524
rect 9221 3512 9227 3524
rect 8767 3484 9227 3512
rect 8767 3472 8773 3484
rect 9221 3472 9227 3484
rect 9279 3472 9285 3524
rect 8 3397 59 3404
rect 1744 3397 1795 3404
rect 3480 3397 3531 3404
rect 5216 3397 5267 3404
rect 6952 3397 7003 3404
rect 8688 3397 8739 3404
rect 9200 3397 9251 3404
rect 1 3345 7 3397
rect 59 3345 65 3397
rect 1737 3345 1743 3397
rect 1795 3345 1801 3397
rect 3473 3345 3479 3397
rect 3531 3345 3537 3397
rect 5209 3345 5215 3397
rect 5267 3345 5273 3397
rect 6945 3345 6951 3397
rect 7003 3345 7009 3397
rect 8681 3345 8687 3397
rect 8739 3345 8745 3397
rect 9193 3345 9199 3397
rect 9251 3385 9257 3397
rect 9251 3357 9521 3385
rect 9251 3345 9257 3357
rect 8 3338 59 3345
rect 1744 3338 1795 3345
rect 3480 3338 3531 3345
rect 5216 3338 5267 3345
rect 6952 3338 7003 3345
rect 8688 3338 8739 3345
rect 9200 3338 9251 3345
rect 35 3295 87 3301
rect 35 3237 87 3243
rect 1771 3295 1823 3301
rect 1771 3237 1823 3243
rect 3507 3295 3559 3301
rect 3507 3237 3559 3243
rect 5243 3295 5295 3301
rect 5243 3237 5295 3243
rect 6979 3295 7031 3301
rect 6979 3237 7031 3243
rect 8715 3295 8767 3301
rect 8715 3237 8767 3243
rect 9227 3295 9279 3301
rect 9227 3237 9279 3243
rect 8 3193 59 3200
rect 1744 3193 1795 3200
rect 3480 3193 3531 3200
rect 5216 3193 5267 3200
rect 6952 3193 7003 3200
rect 8688 3193 8739 3200
rect 9200 3193 9251 3200
rect 1 3141 7 3193
rect 59 3141 65 3193
rect 1737 3141 1743 3193
rect 1795 3141 1801 3193
rect 3473 3141 3479 3193
rect 3531 3141 3537 3193
rect 5209 3141 5215 3193
rect 5267 3141 5273 3193
rect 6945 3141 6951 3193
rect 7003 3141 7009 3193
rect 8681 3141 8687 3193
rect 8739 3141 8745 3193
rect 9193 3141 9199 3193
rect 9251 3141 9257 3193
rect 8 3134 59 3141
rect 1744 3134 1795 3141
rect 3480 3134 3531 3141
rect 5216 3134 5267 3141
rect 6952 3134 7003 3141
rect 8688 3134 8739 3141
rect 9200 3134 9251 3141
rect 35 3091 87 3097
rect 35 3033 87 3039
rect 1771 3091 1823 3097
rect 1771 3033 1823 3039
rect 3507 3091 3559 3097
rect 3507 3033 3559 3039
rect 5243 3091 5295 3097
rect 5243 3033 5295 3039
rect 6979 3091 7031 3097
rect 6979 3033 7031 3039
rect 8715 3091 8767 3097
rect 8715 3033 8767 3039
rect 9227 3091 9279 3097
rect 9227 3033 9279 3039
rect 8 2989 59 2996
rect 1744 2989 1795 2996
rect 3480 2989 3531 2996
rect 5216 2989 5267 2996
rect 6952 2989 7003 2996
rect 8688 2989 8739 2996
rect 9200 2989 9251 2996
rect 1 2937 7 2989
rect 59 2937 65 2989
rect 1737 2937 1743 2989
rect 1795 2937 1801 2989
rect 3473 2937 3479 2989
rect 3531 2937 3537 2989
rect 5209 2937 5215 2989
rect 5267 2937 5273 2989
rect 6945 2937 6951 2989
rect 7003 2937 7009 2989
rect 8681 2937 8687 2989
rect 8739 2937 8745 2989
rect 9193 2937 9199 2989
rect 9251 2937 9257 2989
rect 8 2930 59 2937
rect 1744 2930 1795 2937
rect 3480 2930 3531 2937
rect 5216 2930 5267 2937
rect 6952 2930 7003 2937
rect 8688 2930 8739 2937
rect 9200 2930 9251 2937
rect 35 2887 87 2893
rect 35 2829 87 2835
rect 1771 2887 1823 2893
rect 1771 2829 1823 2835
rect 3507 2887 3559 2893
rect 3507 2829 3559 2835
rect 5243 2887 5295 2893
rect 5243 2829 5295 2835
rect 6979 2887 7031 2893
rect 6979 2829 7031 2835
rect 8715 2887 8767 2893
rect 8715 2829 8767 2835
rect 9227 2887 9279 2893
rect 9227 2829 9279 2835
rect 8 2785 59 2792
rect 1744 2785 1795 2792
rect 3480 2785 3531 2792
rect 5216 2785 5267 2792
rect 6952 2785 7003 2792
rect 8688 2785 8739 2792
rect 9200 2785 9251 2792
rect 1 2733 7 2785
rect 59 2733 65 2785
rect 1737 2733 1743 2785
rect 1795 2733 1801 2785
rect 3473 2733 3479 2785
rect 3531 2733 3537 2785
rect 5209 2733 5215 2785
rect 5267 2733 5273 2785
rect 6945 2733 6951 2785
rect 7003 2733 7009 2785
rect 8681 2733 8687 2785
rect 8739 2733 8745 2785
rect 9193 2733 9199 2785
rect 9251 2733 9257 2785
rect 8 2726 59 2733
rect 1744 2726 1795 2733
rect 3480 2726 3531 2733
rect 5216 2726 5267 2733
rect 6952 2726 7003 2733
rect 8688 2726 8739 2733
rect 9200 2726 9251 2733
rect 35 2683 87 2689
rect 35 2625 87 2631
rect 1771 2683 1823 2689
rect 1771 2625 1823 2631
rect 3507 2683 3559 2689
rect 3507 2625 3559 2631
rect 5243 2683 5295 2689
rect 5243 2625 5295 2631
rect 6979 2683 7031 2689
rect 6979 2625 7031 2631
rect 8715 2683 8767 2689
rect 8715 2625 8767 2631
rect 9227 2683 9279 2689
rect 9227 2625 9279 2631
rect 8 2581 59 2588
rect 1744 2581 1795 2588
rect 3480 2581 3531 2588
rect 5216 2581 5267 2588
rect 6952 2581 7003 2588
rect 8688 2581 8739 2588
rect 9200 2581 9251 2588
rect 1 2529 7 2581
rect 59 2529 65 2581
rect 1737 2529 1743 2581
rect 1795 2529 1801 2581
rect 3473 2529 3479 2581
rect 3531 2529 3537 2581
rect 5209 2529 5215 2581
rect 5267 2529 5273 2581
rect 6945 2529 6951 2581
rect 7003 2529 7009 2581
rect 8681 2529 8687 2581
rect 8739 2529 8745 2581
rect 9193 2529 9199 2581
rect 9251 2529 9257 2581
rect 8 2522 59 2529
rect 1744 2522 1795 2529
rect 3480 2522 3531 2529
rect 5216 2522 5267 2529
rect 6952 2522 7003 2529
rect 8688 2522 8739 2529
rect 9200 2522 9251 2529
rect 35 2479 87 2485
rect 35 2421 87 2427
rect 1771 2479 1823 2485
rect 1771 2421 1823 2427
rect 3507 2479 3559 2485
rect 3507 2421 3559 2427
rect 5243 2479 5295 2485
rect 5243 2421 5295 2427
rect 6979 2479 7031 2485
rect 6979 2421 7031 2427
rect 8715 2479 8767 2485
rect 8715 2421 8767 2427
rect 9227 2479 9279 2485
rect 9227 2421 9279 2427
rect 8 2377 59 2384
rect 1744 2377 1795 2384
rect 3480 2377 3531 2384
rect 5216 2377 5267 2384
rect 6952 2377 7003 2384
rect 8688 2377 8739 2384
rect 9200 2377 9251 2384
rect 1 2325 7 2377
rect 59 2325 65 2377
rect 1737 2325 1743 2377
rect 1795 2325 1801 2377
rect 3473 2325 3479 2377
rect 3531 2325 3537 2377
rect 5209 2325 5215 2377
rect 5267 2325 5273 2377
rect 6945 2325 6951 2377
rect 7003 2325 7009 2377
rect 8681 2325 8687 2377
rect 8739 2325 8745 2377
rect 9193 2325 9199 2377
rect 9251 2325 9257 2377
rect 8 2318 59 2325
rect 1744 2318 1795 2325
rect 3480 2318 3531 2325
rect 5216 2318 5267 2325
rect 6952 2318 7003 2325
rect 8688 2318 8739 2325
rect 9200 2318 9251 2325
rect 35 2275 87 2281
rect 35 2217 87 2223
rect 1771 2275 1823 2281
rect 1771 2217 1823 2223
rect 3507 2275 3559 2281
rect 3507 2217 3559 2223
rect 5243 2275 5295 2281
rect 5243 2217 5295 2223
rect 6979 2275 7031 2281
rect 6979 2217 7031 2223
rect 8715 2275 8767 2281
rect 8715 2217 8767 2223
rect 9227 2275 9279 2281
rect 9227 2217 9279 2223
rect 8 2173 59 2180
rect 1744 2173 1795 2180
rect 3480 2173 3531 2180
rect 5216 2173 5267 2180
rect 6952 2173 7003 2180
rect 8688 2173 8739 2180
rect 9200 2173 9251 2180
rect 1 2121 7 2173
rect 59 2121 65 2173
rect 1737 2121 1743 2173
rect 1795 2121 1801 2173
rect 3473 2121 3479 2173
rect 3531 2121 3537 2173
rect 5209 2121 5215 2173
rect 5267 2121 5273 2173
rect 6945 2121 6951 2173
rect 7003 2121 7009 2173
rect 8681 2121 8687 2173
rect 8739 2121 8745 2173
rect 9193 2121 9199 2173
rect 9251 2121 9257 2173
rect 8 2114 59 2121
rect 1744 2114 1795 2121
rect 3480 2114 3531 2121
rect 5216 2114 5267 2121
rect 6952 2114 7003 2121
rect 8688 2114 8739 2121
rect 9200 2114 9251 2121
rect 35 2071 87 2077
rect 35 2013 87 2019
rect 1771 2071 1823 2077
rect 1771 2013 1823 2019
rect 3507 2071 3559 2077
rect 3507 2013 3559 2019
rect 5243 2071 5295 2077
rect 5243 2013 5295 2019
rect 6979 2071 7031 2077
rect 6979 2013 7031 2019
rect 8715 2071 8767 2077
rect 8715 2013 8767 2019
rect 9227 2071 9279 2077
rect 9227 2013 9279 2019
rect 8 1969 59 1976
rect 1744 1969 1795 1976
rect 3480 1969 3531 1976
rect 5216 1969 5267 1976
rect 6952 1969 7003 1976
rect 8688 1969 8739 1976
rect 9200 1969 9251 1976
rect 1 1917 7 1969
rect 59 1917 65 1969
rect 1737 1917 1743 1969
rect 1795 1917 1801 1969
rect 3473 1917 3479 1969
rect 3531 1917 3537 1969
rect 5209 1917 5215 1969
rect 5267 1917 5273 1969
rect 6945 1917 6951 1969
rect 7003 1917 7009 1969
rect 8681 1917 8687 1969
rect 8739 1917 8745 1969
rect 9193 1917 9199 1969
rect 9251 1917 9257 1969
rect 8 1910 59 1917
rect 1744 1910 1795 1917
rect 3480 1910 3531 1917
rect 5216 1910 5267 1917
rect 6952 1910 7003 1917
rect 8688 1910 8739 1917
rect 9200 1910 9251 1917
rect 35 1867 87 1873
rect 35 1809 87 1815
rect 1771 1867 1823 1873
rect 1771 1809 1823 1815
rect 3507 1867 3559 1873
rect 3507 1809 3559 1815
rect 5243 1867 5295 1873
rect 5243 1809 5295 1815
rect 6979 1867 7031 1873
rect 6979 1809 7031 1815
rect 8715 1867 8767 1873
rect 8715 1809 8767 1815
rect 9227 1867 9279 1873
rect 9227 1809 9279 1815
rect 8 1765 59 1772
rect 1744 1765 1795 1772
rect 3480 1765 3531 1772
rect 5216 1765 5267 1772
rect 6952 1765 7003 1772
rect 8688 1765 8739 1772
rect 9200 1765 9251 1772
rect 1 1713 7 1765
rect 59 1713 65 1765
rect 1737 1713 1743 1765
rect 1795 1713 1801 1765
rect 3473 1713 3479 1765
rect 3531 1713 3537 1765
rect 5209 1713 5215 1765
rect 5267 1713 5273 1765
rect 6945 1713 6951 1765
rect 7003 1713 7009 1765
rect 8681 1713 8687 1765
rect 8739 1713 8745 1765
rect 9193 1713 9199 1765
rect 9251 1713 9257 1765
rect 8 1706 59 1713
rect 1744 1706 1795 1713
rect 3480 1706 3531 1713
rect 5216 1706 5267 1713
rect 6952 1706 7003 1713
rect 8688 1706 8739 1713
rect 9200 1706 9251 1713
rect 35 1663 87 1669
rect 35 1605 87 1611
rect 1771 1663 1823 1669
rect 1771 1605 1823 1611
rect 3507 1663 3559 1669
rect 3507 1605 3559 1611
rect 5243 1663 5295 1669
rect 5243 1605 5295 1611
rect 6979 1663 7031 1669
rect 6979 1605 7031 1611
rect 8715 1663 8767 1669
rect 8715 1605 8767 1611
rect 9227 1663 9279 1669
rect 9227 1605 9279 1611
rect 8 1561 59 1568
rect 1744 1561 1795 1568
rect 3480 1561 3531 1568
rect 5216 1561 5267 1568
rect 6952 1561 7003 1568
rect 8688 1561 8739 1568
rect 9200 1561 9251 1568
rect 1 1509 7 1561
rect 59 1509 65 1561
rect 1737 1509 1743 1561
rect 1795 1509 1801 1561
rect 3473 1509 3479 1561
rect 3531 1509 3537 1561
rect 5209 1509 5215 1561
rect 5267 1509 5273 1561
rect 6945 1509 6951 1561
rect 7003 1509 7009 1561
rect 8681 1509 8687 1561
rect 8739 1509 8745 1561
rect 9193 1509 9199 1561
rect 9251 1509 9257 1561
rect 8 1502 59 1509
rect 1744 1502 1795 1509
rect 3480 1502 3531 1509
rect 5216 1502 5267 1509
rect 6952 1502 7003 1509
rect 8688 1502 8739 1509
rect 9200 1502 9251 1509
rect 35 1459 87 1465
rect 35 1401 87 1407
rect 1771 1459 1823 1465
rect 1771 1401 1823 1407
rect 3507 1459 3559 1465
rect 3507 1401 3559 1407
rect 5243 1459 5295 1465
rect 5243 1401 5295 1407
rect 6979 1459 7031 1465
rect 6979 1401 7031 1407
rect 8715 1459 8767 1465
rect 8715 1401 8767 1407
rect 9227 1459 9279 1465
rect 9227 1401 9279 1407
rect 8 1357 59 1364
rect 1744 1357 1795 1364
rect 3480 1357 3531 1364
rect 5216 1357 5267 1364
rect 6952 1357 7003 1364
rect 8688 1357 8739 1364
rect 9200 1357 9251 1364
rect 1 1305 7 1357
rect 59 1305 65 1357
rect 1737 1305 1743 1357
rect 1795 1305 1801 1357
rect 3473 1305 3479 1357
rect 3531 1305 3537 1357
rect 5209 1305 5215 1357
rect 5267 1305 5273 1357
rect 6945 1305 6951 1357
rect 7003 1305 7009 1357
rect 8681 1305 8687 1357
rect 8739 1305 8745 1357
rect 9193 1305 9199 1357
rect 9251 1305 9257 1357
rect 8 1298 59 1305
rect 1744 1298 1795 1305
rect 3480 1298 3531 1305
rect 5216 1298 5267 1305
rect 6952 1298 7003 1305
rect 8688 1298 8739 1305
rect 9200 1298 9251 1305
rect 35 1255 87 1261
rect 35 1197 87 1203
rect 1771 1255 1823 1261
rect 1771 1197 1823 1203
rect 3507 1255 3559 1261
rect 3507 1197 3559 1203
rect 5243 1255 5295 1261
rect 5243 1197 5295 1203
rect 6979 1255 7031 1261
rect 6979 1197 7031 1203
rect 8715 1255 8767 1261
rect 8715 1197 8767 1203
rect 9227 1255 9279 1261
rect 9227 1197 9279 1203
rect 8 1153 59 1160
rect 1744 1153 1795 1160
rect 3480 1153 3531 1160
rect 5216 1153 5267 1160
rect 6952 1153 7003 1160
rect 8688 1153 8739 1160
rect 9200 1153 9251 1160
rect 1 1101 7 1153
rect 59 1101 65 1153
rect 1737 1101 1743 1153
rect 1795 1101 1801 1153
rect 3473 1101 3479 1153
rect 3531 1101 3537 1153
rect 5209 1101 5215 1153
rect 5267 1101 5273 1153
rect 6945 1101 6951 1153
rect 7003 1101 7009 1153
rect 8681 1101 8687 1153
rect 8739 1101 8745 1153
rect 9193 1101 9199 1153
rect 9251 1101 9257 1153
rect 8 1094 59 1101
rect 1744 1094 1795 1101
rect 3480 1094 3531 1101
rect 5216 1094 5267 1101
rect 6952 1094 7003 1101
rect 8688 1094 8739 1101
rect 9200 1094 9251 1101
rect 35 1051 87 1057
rect 35 993 87 999
rect 1771 1051 1823 1057
rect 1771 993 1823 999
rect 3507 1051 3559 1057
rect 3507 993 3559 999
rect 5243 1051 5295 1057
rect 5243 993 5295 999
rect 6979 1051 7031 1057
rect 6979 993 7031 999
rect 8715 1051 8767 1057
rect 8715 993 8767 999
rect 9227 1051 9279 1057
rect 9227 993 9279 999
rect 8 949 59 956
rect 1744 949 1795 956
rect 3480 949 3531 956
rect 5216 949 5267 956
rect 6952 949 7003 956
rect 8688 949 8739 956
rect 9200 949 9251 956
rect 1 897 7 949
rect 59 897 65 949
rect 1737 897 1743 949
rect 1795 897 1801 949
rect 3473 897 3479 949
rect 3531 897 3537 949
rect 5209 897 5215 949
rect 5267 897 5273 949
rect 6945 897 6951 949
rect 7003 897 7009 949
rect 8681 897 8687 949
rect 8739 897 8745 949
rect 9193 897 9199 949
rect 9251 897 9257 949
rect 8 890 59 897
rect 1744 890 1795 897
rect 3480 890 3531 897
rect 5216 890 5267 897
rect 6952 890 7003 897
rect 8688 890 8739 897
rect 9200 890 9251 897
rect 232 -14 260 873
rect 436 -14 464 873
rect 640 -14 668 873
rect 844 -14 872 873
rect 1048 -14 1076 873
rect 1252 -14 1280 873
rect 1456 -14 1484 873
rect 1660 -14 1688 873
rect 1968 -14 1996 873
rect 2172 -14 2200 873
rect 2376 -14 2404 873
rect 2580 -14 2608 873
rect 2784 -14 2812 873
rect 2988 -14 3016 873
rect 3192 -14 3220 873
rect 3396 -14 3424 873
rect 3704 -14 3732 873
rect 3908 -14 3936 873
rect 4112 -14 4140 873
rect 4316 -14 4344 873
rect 4520 -14 4548 873
rect 4724 -14 4752 873
rect 4928 -14 4956 873
rect 5132 -14 5160 873
rect 5440 -14 5468 873
rect 5644 -14 5672 873
rect 5848 -14 5876 873
rect 6052 -14 6080 873
rect 6256 -14 6284 873
rect 6460 -14 6488 873
rect 6664 -14 6692 873
rect 6868 -14 6896 873
rect 7176 -14 7204 873
rect 7380 -14 7408 873
rect 7584 -14 7612 873
rect 7788 -14 7816 873
rect 7992 -14 8020 873
rect 8196 -14 8224 873
rect 8400 -14 8428 873
rect 8604 -14 8632 873
rect 8912 -14 8940 873
rect 9116 -14 9144 873
rect 9493 396 9521 3357
rect 9267 368 9521 396
<< via1 >>
rect 35 3472 87 3524
rect 1771 3472 1823 3524
rect 3507 3472 3559 3524
rect 5243 3472 5295 3524
rect 6979 3472 7031 3524
rect 8715 3472 8767 3524
rect 9227 3472 9279 3524
rect 7 3388 59 3397
rect 7 3354 16 3388
rect 16 3354 50 3388
rect 50 3354 59 3388
rect 7 3345 59 3354
rect 1743 3388 1795 3397
rect 1743 3354 1752 3388
rect 1752 3354 1786 3388
rect 1786 3354 1795 3388
rect 1743 3345 1795 3354
rect 3479 3388 3531 3397
rect 3479 3354 3488 3388
rect 3488 3354 3522 3388
rect 3522 3354 3531 3388
rect 3479 3345 3531 3354
rect 5215 3388 5267 3397
rect 5215 3354 5224 3388
rect 5224 3354 5258 3388
rect 5258 3354 5267 3388
rect 5215 3345 5267 3354
rect 6951 3388 7003 3397
rect 6951 3354 6960 3388
rect 6960 3354 6994 3388
rect 6994 3354 7003 3388
rect 6951 3345 7003 3354
rect 8687 3388 8739 3397
rect 8687 3354 8696 3388
rect 8696 3354 8730 3388
rect 8730 3354 8739 3388
rect 8687 3345 8739 3354
rect 9199 3388 9251 3397
rect 9199 3354 9208 3388
rect 9208 3354 9242 3388
rect 9242 3354 9251 3388
rect 9199 3345 9251 3354
rect 35 3286 87 3295
rect 35 3252 44 3286
rect 44 3252 78 3286
rect 78 3252 87 3286
rect 35 3243 87 3252
rect 1771 3286 1823 3295
rect 1771 3252 1780 3286
rect 1780 3252 1814 3286
rect 1814 3252 1823 3286
rect 1771 3243 1823 3252
rect 3507 3286 3559 3295
rect 3507 3252 3516 3286
rect 3516 3252 3550 3286
rect 3550 3252 3559 3286
rect 3507 3243 3559 3252
rect 5243 3286 5295 3295
rect 5243 3252 5252 3286
rect 5252 3252 5286 3286
rect 5286 3252 5295 3286
rect 5243 3243 5295 3252
rect 6979 3286 7031 3295
rect 6979 3252 6988 3286
rect 6988 3252 7022 3286
rect 7022 3252 7031 3286
rect 6979 3243 7031 3252
rect 8715 3286 8767 3295
rect 8715 3252 8724 3286
rect 8724 3252 8758 3286
rect 8758 3252 8767 3286
rect 8715 3243 8767 3252
rect 9227 3286 9279 3295
rect 9227 3252 9236 3286
rect 9236 3252 9270 3286
rect 9270 3252 9279 3286
rect 9227 3243 9279 3252
rect 7 3184 59 3193
rect 7 3150 16 3184
rect 16 3150 50 3184
rect 50 3150 59 3184
rect 7 3141 59 3150
rect 1743 3184 1795 3193
rect 1743 3150 1752 3184
rect 1752 3150 1786 3184
rect 1786 3150 1795 3184
rect 1743 3141 1795 3150
rect 3479 3184 3531 3193
rect 3479 3150 3488 3184
rect 3488 3150 3522 3184
rect 3522 3150 3531 3184
rect 3479 3141 3531 3150
rect 5215 3184 5267 3193
rect 5215 3150 5224 3184
rect 5224 3150 5258 3184
rect 5258 3150 5267 3184
rect 5215 3141 5267 3150
rect 6951 3184 7003 3193
rect 6951 3150 6960 3184
rect 6960 3150 6994 3184
rect 6994 3150 7003 3184
rect 6951 3141 7003 3150
rect 8687 3184 8739 3193
rect 8687 3150 8696 3184
rect 8696 3150 8730 3184
rect 8730 3150 8739 3184
rect 8687 3141 8739 3150
rect 9199 3184 9251 3193
rect 9199 3150 9208 3184
rect 9208 3150 9242 3184
rect 9242 3150 9251 3184
rect 9199 3141 9251 3150
rect 35 3082 87 3091
rect 35 3048 44 3082
rect 44 3048 78 3082
rect 78 3048 87 3082
rect 35 3039 87 3048
rect 1771 3082 1823 3091
rect 1771 3048 1780 3082
rect 1780 3048 1814 3082
rect 1814 3048 1823 3082
rect 1771 3039 1823 3048
rect 3507 3082 3559 3091
rect 3507 3048 3516 3082
rect 3516 3048 3550 3082
rect 3550 3048 3559 3082
rect 3507 3039 3559 3048
rect 5243 3082 5295 3091
rect 5243 3048 5252 3082
rect 5252 3048 5286 3082
rect 5286 3048 5295 3082
rect 5243 3039 5295 3048
rect 6979 3082 7031 3091
rect 6979 3048 6988 3082
rect 6988 3048 7022 3082
rect 7022 3048 7031 3082
rect 6979 3039 7031 3048
rect 8715 3082 8767 3091
rect 8715 3048 8724 3082
rect 8724 3048 8758 3082
rect 8758 3048 8767 3082
rect 8715 3039 8767 3048
rect 9227 3082 9279 3091
rect 9227 3048 9236 3082
rect 9236 3048 9270 3082
rect 9270 3048 9279 3082
rect 9227 3039 9279 3048
rect 7 2980 59 2989
rect 7 2946 16 2980
rect 16 2946 50 2980
rect 50 2946 59 2980
rect 7 2937 59 2946
rect 1743 2980 1795 2989
rect 1743 2946 1752 2980
rect 1752 2946 1786 2980
rect 1786 2946 1795 2980
rect 1743 2937 1795 2946
rect 3479 2980 3531 2989
rect 3479 2946 3488 2980
rect 3488 2946 3522 2980
rect 3522 2946 3531 2980
rect 3479 2937 3531 2946
rect 5215 2980 5267 2989
rect 5215 2946 5224 2980
rect 5224 2946 5258 2980
rect 5258 2946 5267 2980
rect 5215 2937 5267 2946
rect 6951 2980 7003 2989
rect 6951 2946 6960 2980
rect 6960 2946 6994 2980
rect 6994 2946 7003 2980
rect 6951 2937 7003 2946
rect 8687 2980 8739 2989
rect 8687 2946 8696 2980
rect 8696 2946 8730 2980
rect 8730 2946 8739 2980
rect 8687 2937 8739 2946
rect 9199 2980 9251 2989
rect 9199 2946 9208 2980
rect 9208 2946 9242 2980
rect 9242 2946 9251 2980
rect 9199 2937 9251 2946
rect 35 2878 87 2887
rect 35 2844 44 2878
rect 44 2844 78 2878
rect 78 2844 87 2878
rect 35 2835 87 2844
rect 1771 2878 1823 2887
rect 1771 2844 1780 2878
rect 1780 2844 1814 2878
rect 1814 2844 1823 2878
rect 1771 2835 1823 2844
rect 3507 2878 3559 2887
rect 3507 2844 3516 2878
rect 3516 2844 3550 2878
rect 3550 2844 3559 2878
rect 3507 2835 3559 2844
rect 5243 2878 5295 2887
rect 5243 2844 5252 2878
rect 5252 2844 5286 2878
rect 5286 2844 5295 2878
rect 5243 2835 5295 2844
rect 6979 2878 7031 2887
rect 6979 2844 6988 2878
rect 6988 2844 7022 2878
rect 7022 2844 7031 2878
rect 6979 2835 7031 2844
rect 8715 2878 8767 2887
rect 8715 2844 8724 2878
rect 8724 2844 8758 2878
rect 8758 2844 8767 2878
rect 8715 2835 8767 2844
rect 9227 2878 9279 2887
rect 9227 2844 9236 2878
rect 9236 2844 9270 2878
rect 9270 2844 9279 2878
rect 9227 2835 9279 2844
rect 7 2776 59 2785
rect 7 2742 16 2776
rect 16 2742 50 2776
rect 50 2742 59 2776
rect 7 2733 59 2742
rect 1743 2776 1795 2785
rect 1743 2742 1752 2776
rect 1752 2742 1786 2776
rect 1786 2742 1795 2776
rect 1743 2733 1795 2742
rect 3479 2776 3531 2785
rect 3479 2742 3488 2776
rect 3488 2742 3522 2776
rect 3522 2742 3531 2776
rect 3479 2733 3531 2742
rect 5215 2776 5267 2785
rect 5215 2742 5224 2776
rect 5224 2742 5258 2776
rect 5258 2742 5267 2776
rect 5215 2733 5267 2742
rect 6951 2776 7003 2785
rect 6951 2742 6960 2776
rect 6960 2742 6994 2776
rect 6994 2742 7003 2776
rect 6951 2733 7003 2742
rect 8687 2776 8739 2785
rect 8687 2742 8696 2776
rect 8696 2742 8730 2776
rect 8730 2742 8739 2776
rect 8687 2733 8739 2742
rect 9199 2776 9251 2785
rect 9199 2742 9208 2776
rect 9208 2742 9242 2776
rect 9242 2742 9251 2776
rect 9199 2733 9251 2742
rect 35 2674 87 2683
rect 35 2640 44 2674
rect 44 2640 78 2674
rect 78 2640 87 2674
rect 35 2631 87 2640
rect 1771 2674 1823 2683
rect 1771 2640 1780 2674
rect 1780 2640 1814 2674
rect 1814 2640 1823 2674
rect 1771 2631 1823 2640
rect 3507 2674 3559 2683
rect 3507 2640 3516 2674
rect 3516 2640 3550 2674
rect 3550 2640 3559 2674
rect 3507 2631 3559 2640
rect 5243 2674 5295 2683
rect 5243 2640 5252 2674
rect 5252 2640 5286 2674
rect 5286 2640 5295 2674
rect 5243 2631 5295 2640
rect 6979 2674 7031 2683
rect 6979 2640 6988 2674
rect 6988 2640 7022 2674
rect 7022 2640 7031 2674
rect 6979 2631 7031 2640
rect 8715 2674 8767 2683
rect 8715 2640 8724 2674
rect 8724 2640 8758 2674
rect 8758 2640 8767 2674
rect 8715 2631 8767 2640
rect 9227 2674 9279 2683
rect 9227 2640 9236 2674
rect 9236 2640 9270 2674
rect 9270 2640 9279 2674
rect 9227 2631 9279 2640
rect 7 2572 59 2581
rect 7 2538 16 2572
rect 16 2538 50 2572
rect 50 2538 59 2572
rect 7 2529 59 2538
rect 1743 2572 1795 2581
rect 1743 2538 1752 2572
rect 1752 2538 1786 2572
rect 1786 2538 1795 2572
rect 1743 2529 1795 2538
rect 3479 2572 3531 2581
rect 3479 2538 3488 2572
rect 3488 2538 3522 2572
rect 3522 2538 3531 2572
rect 3479 2529 3531 2538
rect 5215 2572 5267 2581
rect 5215 2538 5224 2572
rect 5224 2538 5258 2572
rect 5258 2538 5267 2572
rect 5215 2529 5267 2538
rect 6951 2572 7003 2581
rect 6951 2538 6960 2572
rect 6960 2538 6994 2572
rect 6994 2538 7003 2572
rect 6951 2529 7003 2538
rect 8687 2572 8739 2581
rect 8687 2538 8696 2572
rect 8696 2538 8730 2572
rect 8730 2538 8739 2572
rect 8687 2529 8739 2538
rect 9199 2572 9251 2581
rect 9199 2538 9208 2572
rect 9208 2538 9242 2572
rect 9242 2538 9251 2572
rect 9199 2529 9251 2538
rect 35 2470 87 2479
rect 35 2436 44 2470
rect 44 2436 78 2470
rect 78 2436 87 2470
rect 35 2427 87 2436
rect 1771 2470 1823 2479
rect 1771 2436 1780 2470
rect 1780 2436 1814 2470
rect 1814 2436 1823 2470
rect 1771 2427 1823 2436
rect 3507 2470 3559 2479
rect 3507 2436 3516 2470
rect 3516 2436 3550 2470
rect 3550 2436 3559 2470
rect 3507 2427 3559 2436
rect 5243 2470 5295 2479
rect 5243 2436 5252 2470
rect 5252 2436 5286 2470
rect 5286 2436 5295 2470
rect 5243 2427 5295 2436
rect 6979 2470 7031 2479
rect 6979 2436 6988 2470
rect 6988 2436 7022 2470
rect 7022 2436 7031 2470
rect 6979 2427 7031 2436
rect 8715 2470 8767 2479
rect 8715 2436 8724 2470
rect 8724 2436 8758 2470
rect 8758 2436 8767 2470
rect 8715 2427 8767 2436
rect 9227 2470 9279 2479
rect 9227 2436 9236 2470
rect 9236 2436 9270 2470
rect 9270 2436 9279 2470
rect 9227 2427 9279 2436
rect 7 2368 59 2377
rect 7 2334 16 2368
rect 16 2334 50 2368
rect 50 2334 59 2368
rect 7 2325 59 2334
rect 1743 2368 1795 2377
rect 1743 2334 1752 2368
rect 1752 2334 1786 2368
rect 1786 2334 1795 2368
rect 1743 2325 1795 2334
rect 3479 2368 3531 2377
rect 3479 2334 3488 2368
rect 3488 2334 3522 2368
rect 3522 2334 3531 2368
rect 3479 2325 3531 2334
rect 5215 2368 5267 2377
rect 5215 2334 5224 2368
rect 5224 2334 5258 2368
rect 5258 2334 5267 2368
rect 5215 2325 5267 2334
rect 6951 2368 7003 2377
rect 6951 2334 6960 2368
rect 6960 2334 6994 2368
rect 6994 2334 7003 2368
rect 6951 2325 7003 2334
rect 8687 2368 8739 2377
rect 8687 2334 8696 2368
rect 8696 2334 8730 2368
rect 8730 2334 8739 2368
rect 8687 2325 8739 2334
rect 9199 2368 9251 2377
rect 9199 2334 9208 2368
rect 9208 2334 9242 2368
rect 9242 2334 9251 2368
rect 9199 2325 9251 2334
rect 35 2266 87 2275
rect 35 2232 44 2266
rect 44 2232 78 2266
rect 78 2232 87 2266
rect 35 2223 87 2232
rect 1771 2266 1823 2275
rect 1771 2232 1780 2266
rect 1780 2232 1814 2266
rect 1814 2232 1823 2266
rect 1771 2223 1823 2232
rect 3507 2266 3559 2275
rect 3507 2232 3516 2266
rect 3516 2232 3550 2266
rect 3550 2232 3559 2266
rect 3507 2223 3559 2232
rect 5243 2266 5295 2275
rect 5243 2232 5252 2266
rect 5252 2232 5286 2266
rect 5286 2232 5295 2266
rect 5243 2223 5295 2232
rect 6979 2266 7031 2275
rect 6979 2232 6988 2266
rect 6988 2232 7022 2266
rect 7022 2232 7031 2266
rect 6979 2223 7031 2232
rect 8715 2266 8767 2275
rect 8715 2232 8724 2266
rect 8724 2232 8758 2266
rect 8758 2232 8767 2266
rect 8715 2223 8767 2232
rect 9227 2266 9279 2275
rect 9227 2232 9236 2266
rect 9236 2232 9270 2266
rect 9270 2232 9279 2266
rect 9227 2223 9279 2232
rect 7 2164 59 2173
rect 7 2130 16 2164
rect 16 2130 50 2164
rect 50 2130 59 2164
rect 7 2121 59 2130
rect 1743 2164 1795 2173
rect 1743 2130 1752 2164
rect 1752 2130 1786 2164
rect 1786 2130 1795 2164
rect 1743 2121 1795 2130
rect 3479 2164 3531 2173
rect 3479 2130 3488 2164
rect 3488 2130 3522 2164
rect 3522 2130 3531 2164
rect 3479 2121 3531 2130
rect 5215 2164 5267 2173
rect 5215 2130 5224 2164
rect 5224 2130 5258 2164
rect 5258 2130 5267 2164
rect 5215 2121 5267 2130
rect 6951 2164 7003 2173
rect 6951 2130 6960 2164
rect 6960 2130 6994 2164
rect 6994 2130 7003 2164
rect 6951 2121 7003 2130
rect 8687 2164 8739 2173
rect 8687 2130 8696 2164
rect 8696 2130 8730 2164
rect 8730 2130 8739 2164
rect 8687 2121 8739 2130
rect 9199 2164 9251 2173
rect 9199 2130 9208 2164
rect 9208 2130 9242 2164
rect 9242 2130 9251 2164
rect 9199 2121 9251 2130
rect 35 2062 87 2071
rect 35 2028 44 2062
rect 44 2028 78 2062
rect 78 2028 87 2062
rect 35 2019 87 2028
rect 1771 2062 1823 2071
rect 1771 2028 1780 2062
rect 1780 2028 1814 2062
rect 1814 2028 1823 2062
rect 1771 2019 1823 2028
rect 3507 2062 3559 2071
rect 3507 2028 3516 2062
rect 3516 2028 3550 2062
rect 3550 2028 3559 2062
rect 3507 2019 3559 2028
rect 5243 2062 5295 2071
rect 5243 2028 5252 2062
rect 5252 2028 5286 2062
rect 5286 2028 5295 2062
rect 5243 2019 5295 2028
rect 6979 2062 7031 2071
rect 6979 2028 6988 2062
rect 6988 2028 7022 2062
rect 7022 2028 7031 2062
rect 6979 2019 7031 2028
rect 8715 2062 8767 2071
rect 8715 2028 8724 2062
rect 8724 2028 8758 2062
rect 8758 2028 8767 2062
rect 8715 2019 8767 2028
rect 9227 2062 9279 2071
rect 9227 2028 9236 2062
rect 9236 2028 9270 2062
rect 9270 2028 9279 2062
rect 9227 2019 9279 2028
rect 7 1960 59 1969
rect 7 1926 16 1960
rect 16 1926 50 1960
rect 50 1926 59 1960
rect 7 1917 59 1926
rect 1743 1960 1795 1969
rect 1743 1926 1752 1960
rect 1752 1926 1786 1960
rect 1786 1926 1795 1960
rect 1743 1917 1795 1926
rect 3479 1960 3531 1969
rect 3479 1926 3488 1960
rect 3488 1926 3522 1960
rect 3522 1926 3531 1960
rect 3479 1917 3531 1926
rect 5215 1960 5267 1969
rect 5215 1926 5224 1960
rect 5224 1926 5258 1960
rect 5258 1926 5267 1960
rect 5215 1917 5267 1926
rect 6951 1960 7003 1969
rect 6951 1926 6960 1960
rect 6960 1926 6994 1960
rect 6994 1926 7003 1960
rect 6951 1917 7003 1926
rect 8687 1960 8739 1969
rect 8687 1926 8696 1960
rect 8696 1926 8730 1960
rect 8730 1926 8739 1960
rect 8687 1917 8739 1926
rect 9199 1960 9251 1969
rect 9199 1926 9208 1960
rect 9208 1926 9242 1960
rect 9242 1926 9251 1960
rect 9199 1917 9251 1926
rect 35 1858 87 1867
rect 35 1824 44 1858
rect 44 1824 78 1858
rect 78 1824 87 1858
rect 35 1815 87 1824
rect 1771 1858 1823 1867
rect 1771 1824 1780 1858
rect 1780 1824 1814 1858
rect 1814 1824 1823 1858
rect 1771 1815 1823 1824
rect 3507 1858 3559 1867
rect 3507 1824 3516 1858
rect 3516 1824 3550 1858
rect 3550 1824 3559 1858
rect 3507 1815 3559 1824
rect 5243 1858 5295 1867
rect 5243 1824 5252 1858
rect 5252 1824 5286 1858
rect 5286 1824 5295 1858
rect 5243 1815 5295 1824
rect 6979 1858 7031 1867
rect 6979 1824 6988 1858
rect 6988 1824 7022 1858
rect 7022 1824 7031 1858
rect 6979 1815 7031 1824
rect 8715 1858 8767 1867
rect 8715 1824 8724 1858
rect 8724 1824 8758 1858
rect 8758 1824 8767 1858
rect 8715 1815 8767 1824
rect 9227 1858 9279 1867
rect 9227 1824 9236 1858
rect 9236 1824 9270 1858
rect 9270 1824 9279 1858
rect 9227 1815 9279 1824
rect 7 1756 59 1765
rect 7 1722 16 1756
rect 16 1722 50 1756
rect 50 1722 59 1756
rect 7 1713 59 1722
rect 1743 1756 1795 1765
rect 1743 1722 1752 1756
rect 1752 1722 1786 1756
rect 1786 1722 1795 1756
rect 1743 1713 1795 1722
rect 3479 1756 3531 1765
rect 3479 1722 3488 1756
rect 3488 1722 3522 1756
rect 3522 1722 3531 1756
rect 3479 1713 3531 1722
rect 5215 1756 5267 1765
rect 5215 1722 5224 1756
rect 5224 1722 5258 1756
rect 5258 1722 5267 1756
rect 5215 1713 5267 1722
rect 6951 1756 7003 1765
rect 6951 1722 6960 1756
rect 6960 1722 6994 1756
rect 6994 1722 7003 1756
rect 6951 1713 7003 1722
rect 8687 1756 8739 1765
rect 8687 1722 8696 1756
rect 8696 1722 8730 1756
rect 8730 1722 8739 1756
rect 8687 1713 8739 1722
rect 9199 1756 9251 1765
rect 9199 1722 9208 1756
rect 9208 1722 9242 1756
rect 9242 1722 9251 1756
rect 9199 1713 9251 1722
rect 35 1654 87 1663
rect 35 1620 44 1654
rect 44 1620 78 1654
rect 78 1620 87 1654
rect 35 1611 87 1620
rect 1771 1654 1823 1663
rect 1771 1620 1780 1654
rect 1780 1620 1814 1654
rect 1814 1620 1823 1654
rect 1771 1611 1823 1620
rect 3507 1654 3559 1663
rect 3507 1620 3516 1654
rect 3516 1620 3550 1654
rect 3550 1620 3559 1654
rect 3507 1611 3559 1620
rect 5243 1654 5295 1663
rect 5243 1620 5252 1654
rect 5252 1620 5286 1654
rect 5286 1620 5295 1654
rect 5243 1611 5295 1620
rect 6979 1654 7031 1663
rect 6979 1620 6988 1654
rect 6988 1620 7022 1654
rect 7022 1620 7031 1654
rect 6979 1611 7031 1620
rect 8715 1654 8767 1663
rect 8715 1620 8724 1654
rect 8724 1620 8758 1654
rect 8758 1620 8767 1654
rect 8715 1611 8767 1620
rect 9227 1654 9279 1663
rect 9227 1620 9236 1654
rect 9236 1620 9270 1654
rect 9270 1620 9279 1654
rect 9227 1611 9279 1620
rect 7 1552 59 1561
rect 7 1518 16 1552
rect 16 1518 50 1552
rect 50 1518 59 1552
rect 7 1509 59 1518
rect 1743 1552 1795 1561
rect 1743 1518 1752 1552
rect 1752 1518 1786 1552
rect 1786 1518 1795 1552
rect 1743 1509 1795 1518
rect 3479 1552 3531 1561
rect 3479 1518 3488 1552
rect 3488 1518 3522 1552
rect 3522 1518 3531 1552
rect 3479 1509 3531 1518
rect 5215 1552 5267 1561
rect 5215 1518 5224 1552
rect 5224 1518 5258 1552
rect 5258 1518 5267 1552
rect 5215 1509 5267 1518
rect 6951 1552 7003 1561
rect 6951 1518 6960 1552
rect 6960 1518 6994 1552
rect 6994 1518 7003 1552
rect 6951 1509 7003 1518
rect 8687 1552 8739 1561
rect 8687 1518 8696 1552
rect 8696 1518 8730 1552
rect 8730 1518 8739 1552
rect 8687 1509 8739 1518
rect 9199 1552 9251 1561
rect 9199 1518 9208 1552
rect 9208 1518 9242 1552
rect 9242 1518 9251 1552
rect 9199 1509 9251 1518
rect 35 1450 87 1459
rect 35 1416 44 1450
rect 44 1416 78 1450
rect 78 1416 87 1450
rect 35 1407 87 1416
rect 1771 1450 1823 1459
rect 1771 1416 1780 1450
rect 1780 1416 1814 1450
rect 1814 1416 1823 1450
rect 1771 1407 1823 1416
rect 3507 1450 3559 1459
rect 3507 1416 3516 1450
rect 3516 1416 3550 1450
rect 3550 1416 3559 1450
rect 3507 1407 3559 1416
rect 5243 1450 5295 1459
rect 5243 1416 5252 1450
rect 5252 1416 5286 1450
rect 5286 1416 5295 1450
rect 5243 1407 5295 1416
rect 6979 1450 7031 1459
rect 6979 1416 6988 1450
rect 6988 1416 7022 1450
rect 7022 1416 7031 1450
rect 6979 1407 7031 1416
rect 8715 1450 8767 1459
rect 8715 1416 8724 1450
rect 8724 1416 8758 1450
rect 8758 1416 8767 1450
rect 8715 1407 8767 1416
rect 9227 1450 9279 1459
rect 9227 1416 9236 1450
rect 9236 1416 9270 1450
rect 9270 1416 9279 1450
rect 9227 1407 9279 1416
rect 7 1348 59 1357
rect 7 1314 16 1348
rect 16 1314 50 1348
rect 50 1314 59 1348
rect 7 1305 59 1314
rect 1743 1348 1795 1357
rect 1743 1314 1752 1348
rect 1752 1314 1786 1348
rect 1786 1314 1795 1348
rect 1743 1305 1795 1314
rect 3479 1348 3531 1357
rect 3479 1314 3488 1348
rect 3488 1314 3522 1348
rect 3522 1314 3531 1348
rect 3479 1305 3531 1314
rect 5215 1348 5267 1357
rect 5215 1314 5224 1348
rect 5224 1314 5258 1348
rect 5258 1314 5267 1348
rect 5215 1305 5267 1314
rect 6951 1348 7003 1357
rect 6951 1314 6960 1348
rect 6960 1314 6994 1348
rect 6994 1314 7003 1348
rect 6951 1305 7003 1314
rect 8687 1348 8739 1357
rect 8687 1314 8696 1348
rect 8696 1314 8730 1348
rect 8730 1314 8739 1348
rect 8687 1305 8739 1314
rect 9199 1348 9251 1357
rect 9199 1314 9208 1348
rect 9208 1314 9242 1348
rect 9242 1314 9251 1348
rect 9199 1305 9251 1314
rect 35 1246 87 1255
rect 35 1212 44 1246
rect 44 1212 78 1246
rect 78 1212 87 1246
rect 35 1203 87 1212
rect 1771 1246 1823 1255
rect 1771 1212 1780 1246
rect 1780 1212 1814 1246
rect 1814 1212 1823 1246
rect 1771 1203 1823 1212
rect 3507 1246 3559 1255
rect 3507 1212 3516 1246
rect 3516 1212 3550 1246
rect 3550 1212 3559 1246
rect 3507 1203 3559 1212
rect 5243 1246 5295 1255
rect 5243 1212 5252 1246
rect 5252 1212 5286 1246
rect 5286 1212 5295 1246
rect 5243 1203 5295 1212
rect 6979 1246 7031 1255
rect 6979 1212 6988 1246
rect 6988 1212 7022 1246
rect 7022 1212 7031 1246
rect 6979 1203 7031 1212
rect 8715 1246 8767 1255
rect 8715 1212 8724 1246
rect 8724 1212 8758 1246
rect 8758 1212 8767 1246
rect 8715 1203 8767 1212
rect 9227 1246 9279 1255
rect 9227 1212 9236 1246
rect 9236 1212 9270 1246
rect 9270 1212 9279 1246
rect 9227 1203 9279 1212
rect 7 1144 59 1153
rect 7 1110 16 1144
rect 16 1110 50 1144
rect 50 1110 59 1144
rect 7 1101 59 1110
rect 1743 1144 1795 1153
rect 1743 1110 1752 1144
rect 1752 1110 1786 1144
rect 1786 1110 1795 1144
rect 1743 1101 1795 1110
rect 3479 1144 3531 1153
rect 3479 1110 3488 1144
rect 3488 1110 3522 1144
rect 3522 1110 3531 1144
rect 3479 1101 3531 1110
rect 5215 1144 5267 1153
rect 5215 1110 5224 1144
rect 5224 1110 5258 1144
rect 5258 1110 5267 1144
rect 5215 1101 5267 1110
rect 6951 1144 7003 1153
rect 6951 1110 6960 1144
rect 6960 1110 6994 1144
rect 6994 1110 7003 1144
rect 6951 1101 7003 1110
rect 8687 1144 8739 1153
rect 8687 1110 8696 1144
rect 8696 1110 8730 1144
rect 8730 1110 8739 1144
rect 8687 1101 8739 1110
rect 9199 1144 9251 1153
rect 9199 1110 9208 1144
rect 9208 1110 9242 1144
rect 9242 1110 9251 1144
rect 9199 1101 9251 1110
rect 35 1042 87 1051
rect 35 1008 44 1042
rect 44 1008 78 1042
rect 78 1008 87 1042
rect 35 999 87 1008
rect 1771 1042 1823 1051
rect 1771 1008 1780 1042
rect 1780 1008 1814 1042
rect 1814 1008 1823 1042
rect 1771 999 1823 1008
rect 3507 1042 3559 1051
rect 3507 1008 3516 1042
rect 3516 1008 3550 1042
rect 3550 1008 3559 1042
rect 3507 999 3559 1008
rect 5243 1042 5295 1051
rect 5243 1008 5252 1042
rect 5252 1008 5286 1042
rect 5286 1008 5295 1042
rect 5243 999 5295 1008
rect 6979 1042 7031 1051
rect 6979 1008 6988 1042
rect 6988 1008 7022 1042
rect 7022 1008 7031 1042
rect 6979 999 7031 1008
rect 8715 1042 8767 1051
rect 8715 1008 8724 1042
rect 8724 1008 8758 1042
rect 8758 1008 8767 1042
rect 8715 999 8767 1008
rect 9227 1042 9279 1051
rect 9227 1008 9236 1042
rect 9236 1008 9270 1042
rect 9270 1008 9279 1042
rect 9227 999 9279 1008
rect 7 940 59 949
rect 7 906 16 940
rect 16 906 50 940
rect 50 906 59 940
rect 7 897 59 906
rect 1743 940 1795 949
rect 1743 906 1752 940
rect 1752 906 1786 940
rect 1786 906 1795 940
rect 1743 897 1795 906
rect 3479 940 3531 949
rect 3479 906 3488 940
rect 3488 906 3522 940
rect 3522 906 3531 940
rect 3479 897 3531 906
rect 5215 940 5267 949
rect 5215 906 5224 940
rect 5224 906 5258 940
rect 5258 906 5267 940
rect 5215 897 5267 906
rect 6951 940 7003 949
rect 6951 906 6960 940
rect 6960 906 6994 940
rect 6994 906 7003 940
rect 6951 897 7003 906
rect 8687 940 8739 949
rect 8687 906 8696 940
rect 8696 906 8730 940
rect 8730 906 8739 940
rect 8687 897 8739 906
rect 9199 940 9251 949
rect 9199 906 9208 940
rect 9208 906 9242 940
rect 9242 906 9251 940
rect 9199 897 9251 906
<< metal2 >>
rect 33 3527 89 3536
rect 33 3462 89 3471
rect 1769 3527 1825 3536
rect 1769 3462 1825 3471
rect 3505 3527 3561 3536
rect 3505 3462 3561 3471
rect 5241 3527 5297 3536
rect 5241 3462 5297 3471
rect 6977 3527 7033 3536
rect 6977 3462 7033 3471
rect 8713 3527 8769 3536
rect 8713 3462 8769 3471
rect 9225 3527 9281 3536
rect 9225 3462 9281 3471
rect 7 3397 59 3403
rect 1 3350 7 3393
rect 1743 3397 1795 3403
rect 59 3385 65 3393
rect 1737 3385 1743 3393
rect 59 3357 1743 3385
rect 59 3350 65 3357
rect 1737 3350 1743 3357
rect 7 3339 59 3345
rect 3479 3397 3531 3403
rect 1795 3385 1801 3393
rect 3473 3385 3479 3393
rect 1795 3357 3479 3385
rect 1795 3350 1801 3357
rect 3473 3350 3479 3357
rect 1743 3339 1795 3345
rect 5215 3397 5267 3403
rect 3531 3385 3537 3393
rect 5209 3385 5215 3393
rect 3531 3357 5215 3385
rect 3531 3350 3537 3357
rect 5209 3350 5215 3357
rect 3479 3339 3531 3345
rect 6951 3397 7003 3403
rect 5267 3385 5273 3393
rect 6945 3385 6951 3393
rect 5267 3357 6951 3385
rect 5267 3350 5273 3357
rect 6945 3350 6951 3357
rect 5215 3339 5267 3345
rect 8687 3397 8739 3403
rect 7003 3385 7009 3393
rect 8681 3385 8687 3393
rect 7003 3357 8687 3385
rect 7003 3350 7009 3357
rect 8681 3350 8687 3357
rect 6951 3339 7003 3345
rect 9199 3397 9251 3403
rect 8739 3385 8745 3393
rect 9193 3385 9199 3393
rect 8739 3357 9199 3385
rect 8739 3350 8745 3357
rect 9193 3350 9199 3357
rect 8687 3339 8739 3345
rect 9251 3350 9257 3393
rect 9199 3339 9251 3345
rect 24 3241 33 3297
rect 89 3241 98 3297
rect 1760 3241 1769 3297
rect 1825 3241 1834 3297
rect 3496 3241 3505 3297
rect 3561 3241 3570 3297
rect 5232 3241 5241 3297
rect 5297 3241 5306 3297
rect 6968 3241 6977 3297
rect 7033 3241 7042 3297
rect 8704 3241 8713 3297
rect 8769 3241 8778 3297
rect 9216 3241 9225 3297
rect 9281 3241 9290 3297
rect 7 3193 59 3199
rect 1 3146 7 3189
rect 1743 3193 1795 3199
rect 59 3181 65 3189
rect 1737 3181 1743 3189
rect 59 3153 1743 3181
rect 59 3146 65 3153
rect 1737 3146 1743 3153
rect 7 3135 59 3141
rect 3479 3193 3531 3199
rect 1795 3181 1801 3189
rect 3473 3181 3479 3189
rect 1795 3153 3479 3181
rect 1795 3146 1801 3153
rect 3473 3146 3479 3153
rect 1743 3135 1795 3141
rect 5215 3193 5267 3199
rect 3531 3181 3537 3189
rect 5209 3181 5215 3189
rect 3531 3153 5215 3181
rect 3531 3146 3537 3153
rect 5209 3146 5215 3153
rect 3479 3135 3531 3141
rect 6951 3193 7003 3199
rect 5267 3181 5273 3189
rect 6945 3181 6951 3189
rect 5267 3153 6951 3181
rect 5267 3146 5273 3153
rect 6945 3146 6951 3153
rect 5215 3135 5267 3141
rect 8687 3193 8739 3199
rect 7003 3181 7009 3189
rect 8681 3181 8687 3189
rect 7003 3153 8687 3181
rect 7003 3146 7009 3153
rect 8681 3146 8687 3153
rect 6951 3135 7003 3141
rect 9199 3193 9251 3199
rect 8739 3181 8745 3189
rect 9193 3181 9199 3189
rect 8739 3153 9199 3181
rect 8739 3146 8745 3153
rect 9193 3146 9199 3153
rect 8687 3135 8739 3141
rect 9251 3146 9257 3189
rect 9199 3135 9251 3141
rect 24 3037 33 3093
rect 89 3037 98 3093
rect 1760 3037 1769 3093
rect 1825 3037 1834 3093
rect 3496 3037 3505 3093
rect 3561 3037 3570 3093
rect 5232 3037 5241 3093
rect 5297 3037 5306 3093
rect 6968 3037 6977 3093
rect 7033 3037 7042 3093
rect 8704 3037 8713 3093
rect 8769 3037 8778 3093
rect 9216 3037 9225 3093
rect 9281 3037 9290 3093
rect 7 2989 59 2995
rect 1 2942 7 2985
rect 1743 2989 1795 2995
rect 59 2977 65 2985
rect 1737 2977 1743 2985
rect 59 2949 1743 2977
rect 59 2942 65 2949
rect 1737 2942 1743 2949
rect 7 2931 59 2937
rect 3479 2989 3531 2995
rect 1795 2977 1801 2985
rect 3473 2977 3479 2985
rect 1795 2949 3479 2977
rect 1795 2942 1801 2949
rect 3473 2942 3479 2949
rect 1743 2931 1795 2937
rect 5215 2989 5267 2995
rect 3531 2977 3537 2985
rect 5209 2977 5215 2985
rect 3531 2949 5215 2977
rect 3531 2942 3537 2949
rect 5209 2942 5215 2949
rect 3479 2931 3531 2937
rect 6951 2989 7003 2995
rect 5267 2977 5273 2985
rect 6945 2977 6951 2985
rect 5267 2949 6951 2977
rect 5267 2942 5273 2949
rect 6945 2942 6951 2949
rect 5215 2931 5267 2937
rect 8687 2989 8739 2995
rect 7003 2977 7009 2985
rect 8681 2977 8687 2985
rect 7003 2949 8687 2977
rect 7003 2942 7009 2949
rect 8681 2942 8687 2949
rect 6951 2931 7003 2937
rect 9199 2989 9251 2995
rect 8739 2977 8745 2985
rect 9193 2977 9199 2985
rect 8739 2949 9199 2977
rect 8739 2942 8745 2949
rect 9193 2942 9199 2949
rect 8687 2931 8739 2937
rect 9251 2942 9257 2985
rect 9199 2931 9251 2937
rect 24 2833 33 2889
rect 89 2833 98 2889
rect 1760 2833 1769 2889
rect 1825 2833 1834 2889
rect 3496 2833 3505 2889
rect 3561 2833 3570 2889
rect 5232 2833 5241 2889
rect 5297 2833 5306 2889
rect 6968 2833 6977 2889
rect 7033 2833 7042 2889
rect 8704 2833 8713 2889
rect 8769 2833 8778 2889
rect 9216 2833 9225 2889
rect 9281 2833 9290 2889
rect 7 2785 59 2791
rect 1 2738 7 2781
rect 1743 2785 1795 2791
rect 59 2773 65 2781
rect 1737 2773 1743 2781
rect 59 2745 1743 2773
rect 59 2738 65 2745
rect 1737 2738 1743 2745
rect 7 2727 59 2733
rect 3479 2785 3531 2791
rect 1795 2773 1801 2781
rect 3473 2773 3479 2781
rect 1795 2745 3479 2773
rect 1795 2738 1801 2745
rect 3473 2738 3479 2745
rect 1743 2727 1795 2733
rect 5215 2785 5267 2791
rect 3531 2773 3537 2781
rect 5209 2773 5215 2781
rect 3531 2745 5215 2773
rect 3531 2738 3537 2745
rect 5209 2738 5215 2745
rect 3479 2727 3531 2733
rect 6951 2785 7003 2791
rect 5267 2773 5273 2781
rect 6945 2773 6951 2781
rect 5267 2745 6951 2773
rect 5267 2738 5273 2745
rect 6945 2738 6951 2745
rect 5215 2727 5267 2733
rect 8687 2785 8739 2791
rect 7003 2773 7009 2781
rect 8681 2773 8687 2781
rect 7003 2745 8687 2773
rect 7003 2738 7009 2745
rect 8681 2738 8687 2745
rect 6951 2727 7003 2733
rect 9199 2785 9251 2791
rect 8739 2773 8745 2781
rect 9193 2773 9199 2781
rect 8739 2745 9199 2773
rect 8739 2738 8745 2745
rect 9193 2738 9199 2745
rect 8687 2727 8739 2733
rect 9251 2738 9257 2781
rect 9199 2727 9251 2733
rect 24 2629 33 2685
rect 89 2629 98 2685
rect 1760 2629 1769 2685
rect 1825 2629 1834 2685
rect 3496 2629 3505 2685
rect 3561 2629 3570 2685
rect 5232 2629 5241 2685
rect 5297 2629 5306 2685
rect 6968 2629 6977 2685
rect 7033 2629 7042 2685
rect 8704 2629 8713 2685
rect 8769 2629 8778 2685
rect 9216 2629 9225 2685
rect 9281 2629 9290 2685
rect 7 2581 59 2587
rect 1 2534 7 2577
rect 1743 2581 1795 2587
rect 59 2569 65 2577
rect 1737 2569 1743 2577
rect 59 2541 1743 2569
rect 59 2534 65 2541
rect 1737 2534 1743 2541
rect 7 2523 59 2529
rect 3479 2581 3531 2587
rect 1795 2569 1801 2577
rect 3473 2569 3479 2577
rect 1795 2541 3479 2569
rect 1795 2534 1801 2541
rect 3473 2534 3479 2541
rect 1743 2523 1795 2529
rect 5215 2581 5267 2587
rect 3531 2569 3537 2577
rect 5209 2569 5215 2577
rect 3531 2541 5215 2569
rect 3531 2534 3537 2541
rect 5209 2534 5215 2541
rect 3479 2523 3531 2529
rect 6951 2581 7003 2587
rect 5267 2569 5273 2577
rect 6945 2569 6951 2577
rect 5267 2541 6951 2569
rect 5267 2534 5273 2541
rect 6945 2534 6951 2541
rect 5215 2523 5267 2529
rect 8687 2581 8739 2587
rect 7003 2569 7009 2577
rect 8681 2569 8687 2577
rect 7003 2541 8687 2569
rect 7003 2534 7009 2541
rect 8681 2534 8687 2541
rect 6951 2523 7003 2529
rect 9199 2581 9251 2587
rect 8739 2569 8745 2577
rect 9193 2569 9199 2577
rect 8739 2541 9199 2569
rect 8739 2534 8745 2541
rect 9193 2534 9199 2541
rect 8687 2523 8739 2529
rect 9251 2534 9257 2577
rect 9199 2523 9251 2529
rect 24 2425 33 2481
rect 89 2425 98 2481
rect 1760 2425 1769 2481
rect 1825 2425 1834 2481
rect 3496 2425 3505 2481
rect 3561 2425 3570 2481
rect 5232 2425 5241 2481
rect 5297 2425 5306 2481
rect 6968 2425 6977 2481
rect 7033 2425 7042 2481
rect 8704 2425 8713 2481
rect 8769 2425 8778 2481
rect 9216 2425 9225 2481
rect 9281 2425 9290 2481
rect 7 2377 59 2383
rect 1 2330 7 2373
rect 1743 2377 1795 2383
rect 59 2365 65 2373
rect 1737 2365 1743 2373
rect 59 2337 1743 2365
rect 59 2330 65 2337
rect 1737 2330 1743 2337
rect 7 2319 59 2325
rect 3479 2377 3531 2383
rect 1795 2365 1801 2373
rect 3473 2365 3479 2373
rect 1795 2337 3479 2365
rect 1795 2330 1801 2337
rect 3473 2330 3479 2337
rect 1743 2319 1795 2325
rect 5215 2377 5267 2383
rect 3531 2365 3537 2373
rect 5209 2365 5215 2373
rect 3531 2337 5215 2365
rect 3531 2330 3537 2337
rect 5209 2330 5215 2337
rect 3479 2319 3531 2325
rect 6951 2377 7003 2383
rect 5267 2365 5273 2373
rect 6945 2365 6951 2373
rect 5267 2337 6951 2365
rect 5267 2330 5273 2337
rect 6945 2330 6951 2337
rect 5215 2319 5267 2325
rect 8687 2377 8739 2383
rect 7003 2365 7009 2373
rect 8681 2365 8687 2373
rect 7003 2337 8687 2365
rect 7003 2330 7009 2337
rect 8681 2330 8687 2337
rect 6951 2319 7003 2325
rect 9199 2377 9251 2383
rect 8739 2365 8745 2373
rect 9193 2365 9199 2373
rect 8739 2337 9199 2365
rect 8739 2330 8745 2337
rect 9193 2330 9199 2337
rect 8687 2319 8739 2325
rect 9251 2330 9257 2373
rect 9199 2319 9251 2325
rect 24 2221 33 2277
rect 89 2221 98 2277
rect 1760 2221 1769 2277
rect 1825 2221 1834 2277
rect 3496 2221 3505 2277
rect 3561 2221 3570 2277
rect 5232 2221 5241 2277
rect 5297 2221 5306 2277
rect 6968 2221 6977 2277
rect 7033 2221 7042 2277
rect 8704 2221 8713 2277
rect 8769 2221 8778 2277
rect 9216 2221 9225 2277
rect 9281 2221 9290 2277
rect 7 2173 59 2179
rect 1 2126 7 2169
rect 1743 2173 1795 2179
rect 59 2161 65 2169
rect 1737 2161 1743 2169
rect 59 2133 1743 2161
rect 59 2126 65 2133
rect 1737 2126 1743 2133
rect 7 2115 59 2121
rect 3479 2173 3531 2179
rect 1795 2161 1801 2169
rect 3473 2161 3479 2169
rect 1795 2133 3479 2161
rect 1795 2126 1801 2133
rect 3473 2126 3479 2133
rect 1743 2115 1795 2121
rect 5215 2173 5267 2179
rect 3531 2161 3537 2169
rect 5209 2161 5215 2169
rect 3531 2133 5215 2161
rect 3531 2126 3537 2133
rect 5209 2126 5215 2133
rect 3479 2115 3531 2121
rect 6951 2173 7003 2179
rect 5267 2161 5273 2169
rect 6945 2161 6951 2169
rect 5267 2133 6951 2161
rect 5267 2126 5273 2133
rect 6945 2126 6951 2133
rect 5215 2115 5267 2121
rect 8687 2173 8739 2179
rect 7003 2161 7009 2169
rect 8681 2161 8687 2169
rect 7003 2133 8687 2161
rect 7003 2126 7009 2133
rect 8681 2126 8687 2133
rect 6951 2115 7003 2121
rect 9199 2173 9251 2179
rect 8739 2161 8745 2169
rect 9193 2161 9199 2169
rect 8739 2133 9199 2161
rect 8739 2126 8745 2133
rect 9193 2126 9199 2133
rect 8687 2115 8739 2121
rect 9251 2126 9257 2169
rect 9199 2115 9251 2121
rect 24 2017 33 2073
rect 89 2017 98 2073
rect 1760 2017 1769 2073
rect 1825 2017 1834 2073
rect 3496 2017 3505 2073
rect 3561 2017 3570 2073
rect 5232 2017 5241 2073
rect 5297 2017 5306 2073
rect 6968 2017 6977 2073
rect 7033 2017 7042 2073
rect 8704 2017 8713 2073
rect 8769 2017 8778 2073
rect 9216 2017 9225 2073
rect 9281 2017 9290 2073
rect 7 1969 59 1975
rect 1 1922 7 1965
rect 1743 1969 1795 1975
rect 59 1957 65 1965
rect 1737 1957 1743 1965
rect 59 1929 1743 1957
rect 59 1922 65 1929
rect 1737 1922 1743 1929
rect 7 1911 59 1917
rect 3479 1969 3531 1975
rect 1795 1957 1801 1965
rect 3473 1957 3479 1965
rect 1795 1929 3479 1957
rect 1795 1922 1801 1929
rect 3473 1922 3479 1929
rect 1743 1911 1795 1917
rect 5215 1969 5267 1975
rect 3531 1957 3537 1965
rect 5209 1957 5215 1965
rect 3531 1929 5215 1957
rect 3531 1922 3537 1929
rect 5209 1922 5215 1929
rect 3479 1911 3531 1917
rect 6951 1969 7003 1975
rect 5267 1957 5273 1965
rect 6945 1957 6951 1965
rect 5267 1929 6951 1957
rect 5267 1922 5273 1929
rect 6945 1922 6951 1929
rect 5215 1911 5267 1917
rect 8687 1969 8739 1975
rect 7003 1957 7009 1965
rect 8681 1957 8687 1965
rect 7003 1929 8687 1957
rect 7003 1922 7009 1929
rect 8681 1922 8687 1929
rect 6951 1911 7003 1917
rect 9199 1969 9251 1975
rect 8739 1957 8745 1965
rect 9193 1957 9199 1965
rect 8739 1929 9199 1957
rect 8739 1922 8745 1929
rect 9193 1922 9199 1929
rect 8687 1911 8739 1917
rect 9251 1922 9257 1965
rect 9199 1911 9251 1917
rect 24 1813 33 1869
rect 89 1813 98 1869
rect 1760 1813 1769 1869
rect 1825 1813 1834 1869
rect 3496 1813 3505 1869
rect 3561 1813 3570 1869
rect 5232 1813 5241 1869
rect 5297 1813 5306 1869
rect 6968 1813 6977 1869
rect 7033 1813 7042 1869
rect 8704 1813 8713 1869
rect 8769 1813 8778 1869
rect 9216 1813 9225 1869
rect 9281 1813 9290 1869
rect 7 1765 59 1771
rect 1 1718 7 1761
rect 1743 1765 1795 1771
rect 59 1753 65 1761
rect 1737 1753 1743 1761
rect 59 1725 1743 1753
rect 59 1718 65 1725
rect 1737 1718 1743 1725
rect 7 1707 59 1713
rect 3479 1765 3531 1771
rect 1795 1753 1801 1761
rect 3473 1753 3479 1761
rect 1795 1725 3479 1753
rect 1795 1718 1801 1725
rect 3473 1718 3479 1725
rect 1743 1707 1795 1713
rect 5215 1765 5267 1771
rect 3531 1753 3537 1761
rect 5209 1753 5215 1761
rect 3531 1725 5215 1753
rect 3531 1718 3537 1725
rect 5209 1718 5215 1725
rect 3479 1707 3531 1713
rect 6951 1765 7003 1771
rect 5267 1753 5273 1761
rect 6945 1753 6951 1761
rect 5267 1725 6951 1753
rect 5267 1718 5273 1725
rect 6945 1718 6951 1725
rect 5215 1707 5267 1713
rect 8687 1765 8739 1771
rect 7003 1753 7009 1761
rect 8681 1753 8687 1761
rect 7003 1725 8687 1753
rect 7003 1718 7009 1725
rect 8681 1718 8687 1725
rect 6951 1707 7003 1713
rect 9199 1765 9251 1771
rect 8739 1753 8745 1761
rect 9193 1753 9199 1761
rect 8739 1725 9199 1753
rect 8739 1718 8745 1725
rect 9193 1718 9199 1725
rect 8687 1707 8739 1713
rect 9251 1718 9257 1761
rect 9199 1707 9251 1713
rect 24 1609 33 1665
rect 89 1609 98 1665
rect 1760 1609 1769 1665
rect 1825 1609 1834 1665
rect 3496 1609 3505 1665
rect 3561 1609 3570 1665
rect 5232 1609 5241 1665
rect 5297 1609 5306 1665
rect 6968 1609 6977 1665
rect 7033 1609 7042 1665
rect 8704 1609 8713 1665
rect 8769 1609 8778 1665
rect 9216 1609 9225 1665
rect 9281 1609 9290 1665
rect 7 1561 59 1567
rect 1 1514 7 1557
rect 1743 1561 1795 1567
rect 59 1549 65 1557
rect 1737 1549 1743 1557
rect 59 1521 1743 1549
rect 59 1514 65 1521
rect 1737 1514 1743 1521
rect 7 1503 59 1509
rect 3479 1561 3531 1567
rect 1795 1549 1801 1557
rect 3473 1549 3479 1557
rect 1795 1521 3479 1549
rect 1795 1514 1801 1521
rect 3473 1514 3479 1521
rect 1743 1503 1795 1509
rect 5215 1561 5267 1567
rect 3531 1549 3537 1557
rect 5209 1549 5215 1557
rect 3531 1521 5215 1549
rect 3531 1514 3537 1521
rect 5209 1514 5215 1521
rect 3479 1503 3531 1509
rect 6951 1561 7003 1567
rect 5267 1549 5273 1557
rect 6945 1549 6951 1557
rect 5267 1521 6951 1549
rect 5267 1514 5273 1521
rect 6945 1514 6951 1521
rect 5215 1503 5267 1509
rect 8687 1561 8739 1567
rect 7003 1549 7009 1557
rect 8681 1549 8687 1557
rect 7003 1521 8687 1549
rect 7003 1514 7009 1521
rect 8681 1514 8687 1521
rect 6951 1503 7003 1509
rect 9199 1561 9251 1567
rect 8739 1549 8745 1557
rect 9193 1549 9199 1557
rect 8739 1521 9199 1549
rect 8739 1514 8745 1521
rect 9193 1514 9199 1521
rect 8687 1503 8739 1509
rect 9251 1514 9257 1557
rect 9199 1503 9251 1509
rect 24 1405 33 1461
rect 89 1405 98 1461
rect 1760 1405 1769 1461
rect 1825 1405 1834 1461
rect 3496 1405 3505 1461
rect 3561 1405 3570 1461
rect 5232 1405 5241 1461
rect 5297 1405 5306 1461
rect 6968 1405 6977 1461
rect 7033 1405 7042 1461
rect 8704 1405 8713 1461
rect 8769 1405 8778 1461
rect 9216 1405 9225 1461
rect 9281 1405 9290 1461
rect 7 1357 59 1363
rect 1 1310 7 1353
rect 1743 1357 1795 1363
rect 59 1345 65 1353
rect 1737 1345 1743 1353
rect 59 1317 1743 1345
rect 59 1310 65 1317
rect 1737 1310 1743 1317
rect 7 1299 59 1305
rect 3479 1357 3531 1363
rect 1795 1345 1801 1353
rect 3473 1345 3479 1353
rect 1795 1317 3479 1345
rect 1795 1310 1801 1317
rect 3473 1310 3479 1317
rect 1743 1299 1795 1305
rect 5215 1357 5267 1363
rect 3531 1345 3537 1353
rect 5209 1345 5215 1353
rect 3531 1317 5215 1345
rect 3531 1310 3537 1317
rect 5209 1310 5215 1317
rect 3479 1299 3531 1305
rect 6951 1357 7003 1363
rect 5267 1345 5273 1353
rect 6945 1345 6951 1353
rect 5267 1317 6951 1345
rect 5267 1310 5273 1317
rect 6945 1310 6951 1317
rect 5215 1299 5267 1305
rect 8687 1357 8739 1363
rect 7003 1345 7009 1353
rect 8681 1345 8687 1353
rect 7003 1317 8687 1345
rect 7003 1310 7009 1317
rect 8681 1310 8687 1317
rect 6951 1299 7003 1305
rect 9199 1357 9251 1363
rect 8739 1345 8745 1353
rect 9193 1345 9199 1353
rect 8739 1317 9199 1345
rect 8739 1310 8745 1317
rect 9193 1310 9199 1317
rect 8687 1299 8739 1305
rect 9251 1310 9257 1353
rect 9199 1299 9251 1305
rect 24 1201 33 1257
rect 89 1201 98 1257
rect 1760 1201 1769 1257
rect 1825 1201 1834 1257
rect 3496 1201 3505 1257
rect 3561 1201 3570 1257
rect 5232 1201 5241 1257
rect 5297 1201 5306 1257
rect 6968 1201 6977 1257
rect 7033 1201 7042 1257
rect 8704 1201 8713 1257
rect 8769 1201 8778 1257
rect 9216 1201 9225 1257
rect 9281 1201 9290 1257
rect 7 1153 59 1159
rect 1 1106 7 1149
rect 1743 1153 1795 1159
rect 59 1141 65 1149
rect 1737 1141 1743 1149
rect 59 1113 1743 1141
rect 59 1106 65 1113
rect 1737 1106 1743 1113
rect 7 1095 59 1101
rect 3479 1153 3531 1159
rect 1795 1141 1801 1149
rect 3473 1141 3479 1149
rect 1795 1113 3479 1141
rect 1795 1106 1801 1113
rect 3473 1106 3479 1113
rect 1743 1095 1795 1101
rect 5215 1153 5267 1159
rect 3531 1141 3537 1149
rect 5209 1141 5215 1149
rect 3531 1113 5215 1141
rect 3531 1106 3537 1113
rect 5209 1106 5215 1113
rect 3479 1095 3531 1101
rect 6951 1153 7003 1159
rect 5267 1141 5273 1149
rect 6945 1141 6951 1149
rect 5267 1113 6951 1141
rect 5267 1106 5273 1113
rect 6945 1106 6951 1113
rect 5215 1095 5267 1101
rect 8687 1153 8739 1159
rect 7003 1141 7009 1149
rect 8681 1141 8687 1149
rect 7003 1113 8687 1141
rect 7003 1106 7009 1113
rect 8681 1106 8687 1113
rect 6951 1095 7003 1101
rect 9199 1153 9251 1159
rect 8739 1141 8745 1149
rect 9193 1141 9199 1149
rect 8739 1113 9199 1141
rect 8739 1106 8745 1113
rect 9193 1106 9199 1113
rect 8687 1095 8739 1101
rect 9251 1106 9257 1149
rect 9199 1095 9251 1101
rect 24 997 33 1053
rect 89 997 98 1053
rect 1760 997 1769 1053
rect 1825 997 1834 1053
rect 3496 997 3505 1053
rect 3561 997 3570 1053
rect 5232 997 5241 1053
rect 5297 997 5306 1053
rect 6968 997 6977 1053
rect 7033 997 7042 1053
rect 8704 997 8713 1053
rect 8769 997 8778 1053
rect 9216 997 9225 1053
rect 9281 997 9290 1053
rect 7 949 59 955
rect 1 902 7 945
rect 1743 949 1795 955
rect 59 937 65 945
rect 1737 937 1743 945
rect 59 909 1743 937
rect 59 902 65 909
rect 1737 902 1743 909
rect 7 891 59 897
rect 3479 949 3531 955
rect 1795 937 1801 945
rect 3473 937 3479 945
rect 1795 909 3479 937
rect 1795 902 1801 909
rect 3473 902 3479 909
rect 1743 891 1795 897
rect 5215 949 5267 955
rect 3531 937 3537 945
rect 5209 937 5215 945
rect 3531 909 5215 937
rect 3531 902 3537 909
rect 5209 902 5215 909
rect 3479 891 3531 897
rect 6951 949 7003 955
rect 5267 937 5273 945
rect 6945 937 6951 945
rect 5267 909 6951 937
rect 5267 902 5273 909
rect 6945 902 6951 909
rect 5215 891 5267 897
rect 8687 949 8739 955
rect 7003 937 7009 945
rect 8681 937 8687 945
rect 7003 909 8687 937
rect 7003 902 7009 909
rect 8681 902 8687 909
rect 6951 891 7003 897
rect 9199 949 9251 955
rect 8739 937 8745 945
rect 9193 937 9199 945
rect 8739 909 9199 937
rect 8739 902 8745 909
rect 9193 902 9199 909
rect 8687 891 8739 897
rect 9251 902 9257 945
rect 9199 891 9251 897
rect 61 368 89 396
rect 12 -32 40 32
<< via2 >>
rect 33 3524 89 3527
rect 33 3472 35 3524
rect 35 3472 87 3524
rect 87 3472 89 3524
rect 33 3471 89 3472
rect 1769 3524 1825 3527
rect 1769 3472 1771 3524
rect 1771 3472 1823 3524
rect 1823 3472 1825 3524
rect 1769 3471 1825 3472
rect 3505 3524 3561 3527
rect 3505 3472 3507 3524
rect 3507 3472 3559 3524
rect 3559 3472 3561 3524
rect 3505 3471 3561 3472
rect 5241 3524 5297 3527
rect 5241 3472 5243 3524
rect 5243 3472 5295 3524
rect 5295 3472 5297 3524
rect 5241 3471 5297 3472
rect 6977 3524 7033 3527
rect 6977 3472 6979 3524
rect 6979 3472 7031 3524
rect 7031 3472 7033 3524
rect 6977 3471 7033 3472
rect 8713 3524 8769 3527
rect 8713 3472 8715 3524
rect 8715 3472 8767 3524
rect 8767 3472 8769 3524
rect 8713 3471 8769 3472
rect 9225 3524 9281 3527
rect 9225 3472 9227 3524
rect 9227 3472 9279 3524
rect 9279 3472 9281 3524
rect 9225 3471 9281 3472
rect 33 3295 89 3297
rect 33 3243 35 3295
rect 35 3243 87 3295
rect 87 3243 89 3295
rect 33 3241 89 3243
rect 1769 3295 1825 3297
rect 1769 3243 1771 3295
rect 1771 3243 1823 3295
rect 1823 3243 1825 3295
rect 1769 3241 1825 3243
rect 3505 3295 3561 3297
rect 3505 3243 3507 3295
rect 3507 3243 3559 3295
rect 3559 3243 3561 3295
rect 3505 3241 3561 3243
rect 5241 3295 5297 3297
rect 5241 3243 5243 3295
rect 5243 3243 5295 3295
rect 5295 3243 5297 3295
rect 5241 3241 5297 3243
rect 6977 3295 7033 3297
rect 6977 3243 6979 3295
rect 6979 3243 7031 3295
rect 7031 3243 7033 3295
rect 6977 3241 7033 3243
rect 8713 3295 8769 3297
rect 8713 3243 8715 3295
rect 8715 3243 8767 3295
rect 8767 3243 8769 3295
rect 8713 3241 8769 3243
rect 9225 3295 9281 3297
rect 9225 3243 9227 3295
rect 9227 3243 9279 3295
rect 9279 3243 9281 3295
rect 9225 3241 9281 3243
rect 33 3091 89 3093
rect 33 3039 35 3091
rect 35 3039 87 3091
rect 87 3039 89 3091
rect 33 3037 89 3039
rect 1769 3091 1825 3093
rect 1769 3039 1771 3091
rect 1771 3039 1823 3091
rect 1823 3039 1825 3091
rect 1769 3037 1825 3039
rect 3505 3091 3561 3093
rect 3505 3039 3507 3091
rect 3507 3039 3559 3091
rect 3559 3039 3561 3091
rect 3505 3037 3561 3039
rect 5241 3091 5297 3093
rect 5241 3039 5243 3091
rect 5243 3039 5295 3091
rect 5295 3039 5297 3091
rect 5241 3037 5297 3039
rect 6977 3091 7033 3093
rect 6977 3039 6979 3091
rect 6979 3039 7031 3091
rect 7031 3039 7033 3091
rect 6977 3037 7033 3039
rect 8713 3091 8769 3093
rect 8713 3039 8715 3091
rect 8715 3039 8767 3091
rect 8767 3039 8769 3091
rect 8713 3037 8769 3039
rect 9225 3091 9281 3093
rect 9225 3039 9227 3091
rect 9227 3039 9279 3091
rect 9279 3039 9281 3091
rect 9225 3037 9281 3039
rect 33 2887 89 2889
rect 33 2835 35 2887
rect 35 2835 87 2887
rect 87 2835 89 2887
rect 33 2833 89 2835
rect 1769 2887 1825 2889
rect 1769 2835 1771 2887
rect 1771 2835 1823 2887
rect 1823 2835 1825 2887
rect 1769 2833 1825 2835
rect 3505 2887 3561 2889
rect 3505 2835 3507 2887
rect 3507 2835 3559 2887
rect 3559 2835 3561 2887
rect 3505 2833 3561 2835
rect 5241 2887 5297 2889
rect 5241 2835 5243 2887
rect 5243 2835 5295 2887
rect 5295 2835 5297 2887
rect 5241 2833 5297 2835
rect 6977 2887 7033 2889
rect 6977 2835 6979 2887
rect 6979 2835 7031 2887
rect 7031 2835 7033 2887
rect 6977 2833 7033 2835
rect 8713 2887 8769 2889
rect 8713 2835 8715 2887
rect 8715 2835 8767 2887
rect 8767 2835 8769 2887
rect 8713 2833 8769 2835
rect 9225 2887 9281 2889
rect 9225 2835 9227 2887
rect 9227 2835 9279 2887
rect 9279 2835 9281 2887
rect 9225 2833 9281 2835
rect 33 2683 89 2685
rect 33 2631 35 2683
rect 35 2631 87 2683
rect 87 2631 89 2683
rect 33 2629 89 2631
rect 1769 2683 1825 2685
rect 1769 2631 1771 2683
rect 1771 2631 1823 2683
rect 1823 2631 1825 2683
rect 1769 2629 1825 2631
rect 3505 2683 3561 2685
rect 3505 2631 3507 2683
rect 3507 2631 3559 2683
rect 3559 2631 3561 2683
rect 3505 2629 3561 2631
rect 5241 2683 5297 2685
rect 5241 2631 5243 2683
rect 5243 2631 5295 2683
rect 5295 2631 5297 2683
rect 5241 2629 5297 2631
rect 6977 2683 7033 2685
rect 6977 2631 6979 2683
rect 6979 2631 7031 2683
rect 7031 2631 7033 2683
rect 6977 2629 7033 2631
rect 8713 2683 8769 2685
rect 8713 2631 8715 2683
rect 8715 2631 8767 2683
rect 8767 2631 8769 2683
rect 8713 2629 8769 2631
rect 9225 2683 9281 2685
rect 9225 2631 9227 2683
rect 9227 2631 9279 2683
rect 9279 2631 9281 2683
rect 9225 2629 9281 2631
rect 33 2479 89 2481
rect 33 2427 35 2479
rect 35 2427 87 2479
rect 87 2427 89 2479
rect 33 2425 89 2427
rect 1769 2479 1825 2481
rect 1769 2427 1771 2479
rect 1771 2427 1823 2479
rect 1823 2427 1825 2479
rect 1769 2425 1825 2427
rect 3505 2479 3561 2481
rect 3505 2427 3507 2479
rect 3507 2427 3559 2479
rect 3559 2427 3561 2479
rect 3505 2425 3561 2427
rect 5241 2479 5297 2481
rect 5241 2427 5243 2479
rect 5243 2427 5295 2479
rect 5295 2427 5297 2479
rect 5241 2425 5297 2427
rect 6977 2479 7033 2481
rect 6977 2427 6979 2479
rect 6979 2427 7031 2479
rect 7031 2427 7033 2479
rect 6977 2425 7033 2427
rect 8713 2479 8769 2481
rect 8713 2427 8715 2479
rect 8715 2427 8767 2479
rect 8767 2427 8769 2479
rect 8713 2425 8769 2427
rect 9225 2479 9281 2481
rect 9225 2427 9227 2479
rect 9227 2427 9279 2479
rect 9279 2427 9281 2479
rect 9225 2425 9281 2427
rect 33 2275 89 2277
rect 33 2223 35 2275
rect 35 2223 87 2275
rect 87 2223 89 2275
rect 33 2221 89 2223
rect 1769 2275 1825 2277
rect 1769 2223 1771 2275
rect 1771 2223 1823 2275
rect 1823 2223 1825 2275
rect 1769 2221 1825 2223
rect 3505 2275 3561 2277
rect 3505 2223 3507 2275
rect 3507 2223 3559 2275
rect 3559 2223 3561 2275
rect 3505 2221 3561 2223
rect 5241 2275 5297 2277
rect 5241 2223 5243 2275
rect 5243 2223 5295 2275
rect 5295 2223 5297 2275
rect 5241 2221 5297 2223
rect 6977 2275 7033 2277
rect 6977 2223 6979 2275
rect 6979 2223 7031 2275
rect 7031 2223 7033 2275
rect 6977 2221 7033 2223
rect 8713 2275 8769 2277
rect 8713 2223 8715 2275
rect 8715 2223 8767 2275
rect 8767 2223 8769 2275
rect 8713 2221 8769 2223
rect 9225 2275 9281 2277
rect 9225 2223 9227 2275
rect 9227 2223 9279 2275
rect 9279 2223 9281 2275
rect 9225 2221 9281 2223
rect 33 2071 89 2073
rect 33 2019 35 2071
rect 35 2019 87 2071
rect 87 2019 89 2071
rect 33 2017 89 2019
rect 1769 2071 1825 2073
rect 1769 2019 1771 2071
rect 1771 2019 1823 2071
rect 1823 2019 1825 2071
rect 1769 2017 1825 2019
rect 3505 2071 3561 2073
rect 3505 2019 3507 2071
rect 3507 2019 3559 2071
rect 3559 2019 3561 2071
rect 3505 2017 3561 2019
rect 5241 2071 5297 2073
rect 5241 2019 5243 2071
rect 5243 2019 5295 2071
rect 5295 2019 5297 2071
rect 5241 2017 5297 2019
rect 6977 2071 7033 2073
rect 6977 2019 6979 2071
rect 6979 2019 7031 2071
rect 7031 2019 7033 2071
rect 6977 2017 7033 2019
rect 8713 2071 8769 2073
rect 8713 2019 8715 2071
rect 8715 2019 8767 2071
rect 8767 2019 8769 2071
rect 8713 2017 8769 2019
rect 9225 2071 9281 2073
rect 9225 2019 9227 2071
rect 9227 2019 9279 2071
rect 9279 2019 9281 2071
rect 9225 2017 9281 2019
rect 33 1867 89 1869
rect 33 1815 35 1867
rect 35 1815 87 1867
rect 87 1815 89 1867
rect 33 1813 89 1815
rect 1769 1867 1825 1869
rect 1769 1815 1771 1867
rect 1771 1815 1823 1867
rect 1823 1815 1825 1867
rect 1769 1813 1825 1815
rect 3505 1867 3561 1869
rect 3505 1815 3507 1867
rect 3507 1815 3559 1867
rect 3559 1815 3561 1867
rect 3505 1813 3561 1815
rect 5241 1867 5297 1869
rect 5241 1815 5243 1867
rect 5243 1815 5295 1867
rect 5295 1815 5297 1867
rect 5241 1813 5297 1815
rect 6977 1867 7033 1869
rect 6977 1815 6979 1867
rect 6979 1815 7031 1867
rect 7031 1815 7033 1867
rect 6977 1813 7033 1815
rect 8713 1867 8769 1869
rect 8713 1815 8715 1867
rect 8715 1815 8767 1867
rect 8767 1815 8769 1867
rect 8713 1813 8769 1815
rect 9225 1867 9281 1869
rect 9225 1815 9227 1867
rect 9227 1815 9279 1867
rect 9279 1815 9281 1867
rect 9225 1813 9281 1815
rect 33 1663 89 1665
rect 33 1611 35 1663
rect 35 1611 87 1663
rect 87 1611 89 1663
rect 33 1609 89 1611
rect 1769 1663 1825 1665
rect 1769 1611 1771 1663
rect 1771 1611 1823 1663
rect 1823 1611 1825 1663
rect 1769 1609 1825 1611
rect 3505 1663 3561 1665
rect 3505 1611 3507 1663
rect 3507 1611 3559 1663
rect 3559 1611 3561 1663
rect 3505 1609 3561 1611
rect 5241 1663 5297 1665
rect 5241 1611 5243 1663
rect 5243 1611 5295 1663
rect 5295 1611 5297 1663
rect 5241 1609 5297 1611
rect 6977 1663 7033 1665
rect 6977 1611 6979 1663
rect 6979 1611 7031 1663
rect 7031 1611 7033 1663
rect 6977 1609 7033 1611
rect 8713 1663 8769 1665
rect 8713 1611 8715 1663
rect 8715 1611 8767 1663
rect 8767 1611 8769 1663
rect 8713 1609 8769 1611
rect 9225 1663 9281 1665
rect 9225 1611 9227 1663
rect 9227 1611 9279 1663
rect 9279 1611 9281 1663
rect 9225 1609 9281 1611
rect 33 1459 89 1461
rect 33 1407 35 1459
rect 35 1407 87 1459
rect 87 1407 89 1459
rect 33 1405 89 1407
rect 1769 1459 1825 1461
rect 1769 1407 1771 1459
rect 1771 1407 1823 1459
rect 1823 1407 1825 1459
rect 1769 1405 1825 1407
rect 3505 1459 3561 1461
rect 3505 1407 3507 1459
rect 3507 1407 3559 1459
rect 3559 1407 3561 1459
rect 3505 1405 3561 1407
rect 5241 1459 5297 1461
rect 5241 1407 5243 1459
rect 5243 1407 5295 1459
rect 5295 1407 5297 1459
rect 5241 1405 5297 1407
rect 6977 1459 7033 1461
rect 6977 1407 6979 1459
rect 6979 1407 7031 1459
rect 7031 1407 7033 1459
rect 6977 1405 7033 1407
rect 8713 1459 8769 1461
rect 8713 1407 8715 1459
rect 8715 1407 8767 1459
rect 8767 1407 8769 1459
rect 8713 1405 8769 1407
rect 9225 1459 9281 1461
rect 9225 1407 9227 1459
rect 9227 1407 9279 1459
rect 9279 1407 9281 1459
rect 9225 1405 9281 1407
rect 33 1255 89 1257
rect 33 1203 35 1255
rect 35 1203 87 1255
rect 87 1203 89 1255
rect 33 1201 89 1203
rect 1769 1255 1825 1257
rect 1769 1203 1771 1255
rect 1771 1203 1823 1255
rect 1823 1203 1825 1255
rect 1769 1201 1825 1203
rect 3505 1255 3561 1257
rect 3505 1203 3507 1255
rect 3507 1203 3559 1255
rect 3559 1203 3561 1255
rect 3505 1201 3561 1203
rect 5241 1255 5297 1257
rect 5241 1203 5243 1255
rect 5243 1203 5295 1255
rect 5295 1203 5297 1255
rect 5241 1201 5297 1203
rect 6977 1255 7033 1257
rect 6977 1203 6979 1255
rect 6979 1203 7031 1255
rect 7031 1203 7033 1255
rect 6977 1201 7033 1203
rect 8713 1255 8769 1257
rect 8713 1203 8715 1255
rect 8715 1203 8767 1255
rect 8767 1203 8769 1255
rect 8713 1201 8769 1203
rect 9225 1255 9281 1257
rect 9225 1203 9227 1255
rect 9227 1203 9279 1255
rect 9279 1203 9281 1255
rect 9225 1201 9281 1203
rect 33 1051 89 1053
rect 33 999 35 1051
rect 35 999 87 1051
rect 87 999 89 1051
rect 33 997 89 999
rect 1769 1051 1825 1053
rect 1769 999 1771 1051
rect 1771 999 1823 1051
rect 1823 999 1825 1051
rect 1769 997 1825 999
rect 3505 1051 3561 1053
rect 3505 999 3507 1051
rect 3507 999 3559 1051
rect 3559 999 3561 1051
rect 3505 997 3561 999
rect 5241 1051 5297 1053
rect 5241 999 5243 1051
rect 5243 999 5295 1051
rect 5295 999 5297 1051
rect 5241 997 5297 999
rect 6977 1051 7033 1053
rect 6977 999 6979 1051
rect 6979 999 7031 1051
rect 7031 999 7033 1051
rect 6977 997 7033 999
rect 8713 1051 8769 1053
rect 8713 999 8715 1051
rect 8715 999 8767 1051
rect 8767 999 8769 1051
rect 8713 997 8769 999
rect 9225 1051 9281 1053
rect 9225 999 9227 1051
rect 9227 999 9279 1051
rect 9279 999 9281 1051
rect 9225 997 9281 999
<< metal3 >>
rect 28 3527 94 3532
rect 28 3471 33 3527
rect 89 3471 94 3527
rect 28 3466 94 3471
rect 1764 3527 1830 3532
rect 1764 3471 1769 3527
rect 1825 3471 1830 3527
rect 1764 3466 1830 3471
rect 3500 3527 3566 3532
rect 3500 3471 3505 3527
rect 3561 3471 3566 3527
rect 3500 3466 3566 3471
rect 5236 3527 5302 3532
rect 5236 3471 5241 3527
rect 5297 3471 5302 3527
rect 5236 3466 5302 3471
rect 6972 3527 7038 3532
rect 6972 3471 6977 3527
rect 7033 3471 7038 3527
rect 6972 3466 7038 3471
rect 8708 3527 8774 3532
rect 8708 3471 8713 3527
rect 8769 3471 8774 3527
rect 8708 3466 8774 3471
rect 9220 3527 9286 3532
rect 9220 3471 9225 3527
rect 9281 3471 9286 3527
rect 9220 3466 9286 3471
rect 31 3302 91 3466
rect 1767 3302 1827 3466
rect 3503 3302 3563 3466
rect 5239 3302 5299 3466
rect 6975 3302 7035 3466
rect 8711 3302 8771 3466
rect 9223 3302 9283 3466
rect 28 3297 94 3302
rect 28 3241 33 3297
rect 89 3241 94 3297
rect 28 3236 94 3241
rect 1764 3297 1830 3302
rect 1764 3241 1769 3297
rect 1825 3241 1830 3297
rect 1764 3236 1830 3241
rect 3500 3297 3566 3302
rect 3500 3241 3505 3297
rect 3561 3241 3566 3297
rect 3500 3236 3566 3241
rect 5236 3297 5302 3302
rect 5236 3241 5241 3297
rect 5297 3241 5302 3297
rect 5236 3236 5302 3241
rect 6972 3297 7038 3302
rect 6972 3241 6977 3297
rect 7033 3241 7038 3297
rect 6972 3236 7038 3241
rect 8708 3297 8774 3302
rect 8708 3241 8713 3297
rect 8769 3241 8774 3297
rect 8708 3236 8774 3241
rect 9220 3297 9286 3302
rect 9220 3241 9225 3297
rect 9281 3241 9286 3297
rect 9220 3236 9286 3241
rect 31 3098 91 3236
rect 1767 3098 1827 3236
rect 3503 3098 3563 3236
rect 5239 3098 5299 3236
rect 6975 3098 7035 3236
rect 8711 3098 8771 3236
rect 9223 3098 9283 3236
rect 28 3093 94 3098
rect 28 3037 33 3093
rect 89 3037 94 3093
rect 28 3032 94 3037
rect 1764 3093 1830 3098
rect 1764 3037 1769 3093
rect 1825 3037 1830 3093
rect 1764 3032 1830 3037
rect 3500 3093 3566 3098
rect 3500 3037 3505 3093
rect 3561 3037 3566 3093
rect 3500 3032 3566 3037
rect 5236 3093 5302 3098
rect 5236 3037 5241 3093
rect 5297 3037 5302 3093
rect 5236 3032 5302 3037
rect 6972 3093 7038 3098
rect 6972 3037 6977 3093
rect 7033 3037 7038 3093
rect 6972 3032 7038 3037
rect 8708 3093 8774 3098
rect 8708 3037 8713 3093
rect 8769 3037 8774 3093
rect 8708 3032 8774 3037
rect 9220 3093 9286 3098
rect 9220 3037 9225 3093
rect 9281 3037 9286 3093
rect 9220 3032 9286 3037
rect 31 2894 91 3032
rect 1767 2894 1827 3032
rect 3503 2894 3563 3032
rect 5239 2894 5299 3032
rect 6975 2894 7035 3032
rect 8711 2894 8771 3032
rect 9223 2894 9283 3032
rect 28 2889 94 2894
rect 28 2833 33 2889
rect 89 2833 94 2889
rect 28 2828 94 2833
rect 1764 2889 1830 2894
rect 1764 2833 1769 2889
rect 1825 2833 1830 2889
rect 1764 2828 1830 2833
rect 3500 2889 3566 2894
rect 3500 2833 3505 2889
rect 3561 2833 3566 2889
rect 3500 2828 3566 2833
rect 5236 2889 5302 2894
rect 5236 2833 5241 2889
rect 5297 2833 5302 2889
rect 5236 2828 5302 2833
rect 6972 2889 7038 2894
rect 6972 2833 6977 2889
rect 7033 2833 7038 2889
rect 6972 2828 7038 2833
rect 8708 2889 8774 2894
rect 8708 2833 8713 2889
rect 8769 2833 8774 2889
rect 8708 2828 8774 2833
rect 9220 2889 9286 2894
rect 9220 2833 9225 2889
rect 9281 2833 9286 2889
rect 9220 2828 9286 2833
rect 31 2690 91 2828
rect 1767 2690 1827 2828
rect 3503 2690 3563 2828
rect 5239 2690 5299 2828
rect 6975 2690 7035 2828
rect 8711 2690 8771 2828
rect 9223 2690 9283 2828
rect 28 2685 94 2690
rect 28 2629 33 2685
rect 89 2629 94 2685
rect 28 2624 94 2629
rect 1764 2685 1830 2690
rect 1764 2629 1769 2685
rect 1825 2629 1830 2685
rect 1764 2624 1830 2629
rect 3500 2685 3566 2690
rect 3500 2629 3505 2685
rect 3561 2629 3566 2685
rect 3500 2624 3566 2629
rect 5236 2685 5302 2690
rect 5236 2629 5241 2685
rect 5297 2629 5302 2685
rect 5236 2624 5302 2629
rect 6972 2685 7038 2690
rect 6972 2629 6977 2685
rect 7033 2629 7038 2685
rect 6972 2624 7038 2629
rect 8708 2685 8774 2690
rect 8708 2629 8713 2685
rect 8769 2629 8774 2685
rect 8708 2624 8774 2629
rect 9220 2685 9286 2690
rect 9220 2629 9225 2685
rect 9281 2629 9286 2685
rect 9220 2624 9286 2629
rect 31 2486 91 2624
rect 1767 2486 1827 2624
rect 3503 2486 3563 2624
rect 5239 2486 5299 2624
rect 6975 2486 7035 2624
rect 8711 2486 8771 2624
rect 9223 2486 9283 2624
rect 28 2481 94 2486
rect 28 2425 33 2481
rect 89 2425 94 2481
rect 28 2420 94 2425
rect 1764 2481 1830 2486
rect 1764 2425 1769 2481
rect 1825 2425 1830 2481
rect 1764 2420 1830 2425
rect 3500 2481 3566 2486
rect 3500 2425 3505 2481
rect 3561 2425 3566 2481
rect 3500 2420 3566 2425
rect 5236 2481 5302 2486
rect 5236 2425 5241 2481
rect 5297 2425 5302 2481
rect 5236 2420 5302 2425
rect 6972 2481 7038 2486
rect 6972 2425 6977 2481
rect 7033 2425 7038 2481
rect 6972 2420 7038 2425
rect 8708 2481 8774 2486
rect 8708 2425 8713 2481
rect 8769 2425 8774 2481
rect 8708 2420 8774 2425
rect 9220 2481 9286 2486
rect 9220 2425 9225 2481
rect 9281 2425 9286 2481
rect 9220 2420 9286 2425
rect 31 2282 91 2420
rect 1767 2282 1827 2420
rect 3503 2282 3563 2420
rect 5239 2282 5299 2420
rect 6975 2282 7035 2420
rect 8711 2282 8771 2420
rect 9223 2282 9283 2420
rect 28 2277 94 2282
rect 28 2221 33 2277
rect 89 2221 94 2277
rect 28 2216 94 2221
rect 1764 2277 1830 2282
rect 1764 2221 1769 2277
rect 1825 2221 1830 2277
rect 1764 2216 1830 2221
rect 3500 2277 3566 2282
rect 3500 2221 3505 2277
rect 3561 2221 3566 2277
rect 3500 2216 3566 2221
rect 5236 2277 5302 2282
rect 5236 2221 5241 2277
rect 5297 2221 5302 2277
rect 5236 2216 5302 2221
rect 6972 2277 7038 2282
rect 6972 2221 6977 2277
rect 7033 2221 7038 2277
rect 6972 2216 7038 2221
rect 8708 2277 8774 2282
rect 8708 2221 8713 2277
rect 8769 2221 8774 2277
rect 8708 2216 8774 2221
rect 9220 2277 9286 2282
rect 9220 2221 9225 2277
rect 9281 2221 9286 2277
rect 9220 2216 9286 2221
rect 31 2078 91 2216
rect 1767 2078 1827 2216
rect 3503 2078 3563 2216
rect 5239 2078 5299 2216
rect 6975 2078 7035 2216
rect 8711 2078 8771 2216
rect 9223 2078 9283 2216
rect 28 2073 94 2078
rect 28 2017 33 2073
rect 89 2017 94 2073
rect 28 2012 94 2017
rect 1764 2073 1830 2078
rect 1764 2017 1769 2073
rect 1825 2017 1830 2073
rect 1764 2012 1830 2017
rect 3500 2073 3566 2078
rect 3500 2017 3505 2073
rect 3561 2017 3566 2073
rect 3500 2012 3566 2017
rect 5236 2073 5302 2078
rect 5236 2017 5241 2073
rect 5297 2017 5302 2073
rect 5236 2012 5302 2017
rect 6972 2073 7038 2078
rect 6972 2017 6977 2073
rect 7033 2017 7038 2073
rect 6972 2012 7038 2017
rect 8708 2073 8774 2078
rect 8708 2017 8713 2073
rect 8769 2017 8774 2073
rect 8708 2012 8774 2017
rect 9220 2073 9286 2078
rect 9220 2017 9225 2073
rect 9281 2017 9286 2073
rect 9220 2012 9286 2017
rect 31 1874 91 2012
rect 1767 1874 1827 2012
rect 3503 1874 3563 2012
rect 5239 1874 5299 2012
rect 6975 1874 7035 2012
rect 8711 1874 8771 2012
rect 9223 1874 9283 2012
rect 28 1869 94 1874
rect 28 1813 33 1869
rect 89 1813 94 1869
rect 28 1808 94 1813
rect 1764 1869 1830 1874
rect 1764 1813 1769 1869
rect 1825 1813 1830 1869
rect 1764 1808 1830 1813
rect 3500 1869 3566 1874
rect 3500 1813 3505 1869
rect 3561 1813 3566 1869
rect 3500 1808 3566 1813
rect 5236 1869 5302 1874
rect 5236 1813 5241 1869
rect 5297 1813 5302 1869
rect 5236 1808 5302 1813
rect 6972 1869 7038 1874
rect 6972 1813 6977 1869
rect 7033 1813 7038 1869
rect 6972 1808 7038 1813
rect 8708 1869 8774 1874
rect 8708 1813 8713 1869
rect 8769 1813 8774 1869
rect 8708 1808 8774 1813
rect 9220 1869 9286 1874
rect 9220 1813 9225 1869
rect 9281 1813 9286 1869
rect 9220 1808 9286 1813
rect 31 1670 91 1808
rect 1767 1670 1827 1808
rect 3503 1670 3563 1808
rect 5239 1670 5299 1808
rect 6975 1670 7035 1808
rect 8711 1670 8771 1808
rect 9223 1670 9283 1808
rect 28 1665 94 1670
rect 28 1609 33 1665
rect 89 1609 94 1665
rect 28 1604 94 1609
rect 1764 1665 1830 1670
rect 1764 1609 1769 1665
rect 1825 1609 1830 1665
rect 1764 1604 1830 1609
rect 3500 1665 3566 1670
rect 3500 1609 3505 1665
rect 3561 1609 3566 1665
rect 3500 1604 3566 1609
rect 5236 1665 5302 1670
rect 5236 1609 5241 1665
rect 5297 1609 5302 1665
rect 5236 1604 5302 1609
rect 6972 1665 7038 1670
rect 6972 1609 6977 1665
rect 7033 1609 7038 1665
rect 6972 1604 7038 1609
rect 8708 1665 8774 1670
rect 8708 1609 8713 1665
rect 8769 1609 8774 1665
rect 8708 1604 8774 1609
rect 9220 1665 9286 1670
rect 9220 1609 9225 1665
rect 9281 1609 9286 1665
rect 9220 1604 9286 1609
rect 31 1466 91 1604
rect 1767 1466 1827 1604
rect 3503 1466 3563 1604
rect 5239 1466 5299 1604
rect 6975 1466 7035 1604
rect 8711 1466 8771 1604
rect 9223 1466 9283 1604
rect 28 1461 94 1466
rect 28 1405 33 1461
rect 89 1405 94 1461
rect 28 1400 94 1405
rect 1764 1461 1830 1466
rect 1764 1405 1769 1461
rect 1825 1405 1830 1461
rect 1764 1400 1830 1405
rect 3500 1461 3566 1466
rect 3500 1405 3505 1461
rect 3561 1405 3566 1461
rect 3500 1400 3566 1405
rect 5236 1461 5302 1466
rect 5236 1405 5241 1461
rect 5297 1405 5302 1461
rect 5236 1400 5302 1405
rect 6972 1461 7038 1466
rect 6972 1405 6977 1461
rect 7033 1405 7038 1461
rect 6972 1400 7038 1405
rect 8708 1461 8774 1466
rect 8708 1405 8713 1461
rect 8769 1405 8774 1461
rect 8708 1400 8774 1405
rect 9220 1461 9286 1466
rect 9220 1405 9225 1461
rect 9281 1405 9286 1461
rect 9220 1400 9286 1405
rect 31 1262 91 1400
rect 1767 1262 1827 1400
rect 3503 1262 3563 1400
rect 5239 1262 5299 1400
rect 6975 1262 7035 1400
rect 8711 1262 8771 1400
rect 9223 1262 9283 1400
rect 28 1257 94 1262
rect 28 1201 33 1257
rect 89 1201 94 1257
rect 28 1196 94 1201
rect 1764 1257 1830 1262
rect 1764 1201 1769 1257
rect 1825 1201 1830 1257
rect 1764 1196 1830 1201
rect 3500 1257 3566 1262
rect 3500 1201 3505 1257
rect 3561 1201 3566 1257
rect 3500 1196 3566 1201
rect 5236 1257 5302 1262
rect 5236 1201 5241 1257
rect 5297 1201 5302 1257
rect 5236 1196 5302 1201
rect 6972 1257 7038 1262
rect 6972 1201 6977 1257
rect 7033 1201 7038 1257
rect 6972 1196 7038 1201
rect 8708 1257 8774 1262
rect 8708 1201 8713 1257
rect 8769 1201 8774 1257
rect 8708 1196 8774 1201
rect 9220 1257 9286 1262
rect 9220 1201 9225 1257
rect 9281 1201 9286 1257
rect 9220 1196 9286 1201
rect 31 1058 91 1196
rect 1767 1058 1827 1196
rect 3503 1058 3563 1196
rect 5239 1058 5299 1196
rect 6975 1058 7035 1196
rect 8711 1058 8771 1196
rect 9223 1058 9283 1196
rect 28 1053 94 1058
rect 28 997 33 1053
rect 89 997 94 1053
rect 28 992 94 997
rect 1764 1053 1830 1058
rect 1764 997 1769 1053
rect 1825 997 1830 1053
rect 1764 992 1830 997
rect 3500 1053 3566 1058
rect 3500 997 3505 1053
rect 3561 997 3566 1053
rect 3500 992 3566 997
rect 5236 1053 5302 1058
rect 5236 997 5241 1053
rect 5297 997 5302 1053
rect 5236 992 5302 997
rect 6972 1053 7038 1058
rect 6972 997 6977 1053
rect 7033 997 7038 1053
rect 6972 992 7038 997
rect 8708 1053 8774 1058
rect 8708 997 8713 1053
rect 8769 997 8774 1053
rect 8708 992 8774 997
rect 9220 1053 9286 1058
rect 9220 997 9225 1053
rect 9281 997 9286 1053
rect 9220 992 9286 997
rect 31 978 91 992
rect 1767 978 1827 992
rect 3503 978 3563 992
rect 5239 978 5299 992
rect 6975 978 7035 992
rect 8711 978 8771 992
rect 9223 978 9283 992
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_0
timestamp 1581321262
transform 1 0 8988 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1
timestamp 1581321262
transform 1 0 8784 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_2
timestamp 1581321262
transform 1 0 8476 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_3
timestamp 1581321262
transform 1 0 8272 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_4
timestamp 1581321262
transform 1 0 8068 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_5
timestamp 1581321262
transform 1 0 7864 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_6
timestamp 1581321262
transform 1 0 7660 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_7
timestamp 1581321262
transform 1 0 7456 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_8
timestamp 1581321262
transform 1 0 7252 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_9
timestamp 1581321262
transform 1 0 7048 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_10
timestamp 1581321262
transform 1 0 6740 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_11
timestamp 1581321262
transform 1 0 6536 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_12
timestamp 1581321262
transform 1 0 6332 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_13
timestamp 1581321262
transform 1 0 6128 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_14
timestamp 1581321262
transform 1 0 5924 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_15
timestamp 1581321262
transform 1 0 5720 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_16
timestamp 1581321262
transform 1 0 5516 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_17
timestamp 1581321262
transform 1 0 5312 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_18
timestamp 1581321262
transform 1 0 5004 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_19
timestamp 1581321262
transform 1 0 4800 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_20
timestamp 1581321262
transform 1 0 4596 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_21
timestamp 1581321262
transform 1 0 4392 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_22
timestamp 1581321262
transform 1 0 4188 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_23
timestamp 1581321262
transform 1 0 3984 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_24
timestamp 1581321262
transform 1 0 3780 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_25
timestamp 1581321262
transform 1 0 3576 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_26
timestamp 1581321262
transform 1 0 3268 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_27
timestamp 1581321262
transform 1 0 3064 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_28
timestamp 1581321262
transform 1 0 2860 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_29
timestamp 1581321262
transform 1 0 2656 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_30
timestamp 1581321262
transform 1 0 2452 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_31
timestamp 1581321262
transform 1 0 2248 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_32
timestamp 1581321262
transform 1 0 2044 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_33
timestamp 1581321262
transform 1 0 1840 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_34
timestamp 1581321262
transform 1 0 1532 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_35
timestamp 1581321262
transform 1 0 1328 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_36
timestamp 1581321262
transform 1 0 1124 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_37
timestamp 1581321262
transform 1 0 920 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_38
timestamp 1581321262
transform 1 0 716 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_39
timestamp 1581321262
transform 1 0 512 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_40
timestamp 1581321262
transform 1 0 308 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_41
timestamp 1581321262
transform 1 0 104 0 1 3321
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_42
timestamp 1581321262
transform 1 0 8988 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_43
timestamp 1581321262
transform 1 0 8476 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_44
timestamp 1581321262
transform 1 0 8068 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_45
timestamp 1581321262
transform 1 0 7660 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_46
timestamp 1581321262
transform 1 0 7252 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_47
timestamp 1581321262
transform 1 0 6740 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_48
timestamp 1581321262
transform 1 0 6332 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_49
timestamp 1581321262
transform 1 0 5924 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_50
timestamp 1581321262
transform 1 0 5516 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_51
timestamp 1581321262
transform 1 0 5004 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_52
timestamp 1581321262
transform 1 0 4596 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_53
timestamp 1581321262
transform 1 0 4188 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_54
timestamp 1581321262
transform 1 0 3780 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_55
timestamp 1581321262
transform 1 0 3268 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_56
timestamp 1581321262
transform 1 0 2860 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_57
timestamp 1581321262
transform 1 0 2452 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_58
timestamp 1581321262
transform 1 0 2044 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_59
timestamp 1581321262
transform 1 0 1532 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_60
timestamp 1581321262
transform 1 0 1124 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_61
timestamp 1581321262
transform 1 0 716 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_62
timestamp 1581321262
transform 1 0 308 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_63
timestamp 1581321262
transform 1 0 8784 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_64
timestamp 1581321262
transform 1 0 8272 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_65
timestamp 1581321262
transform 1 0 7864 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_66
timestamp 1581321262
transform 1 0 7456 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_67
timestamp 1581321262
transform 1 0 7048 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_68
timestamp 1581321262
transform 1 0 6536 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_69
timestamp 1581321262
transform 1 0 6128 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_70
timestamp 1581321262
transform 1 0 5720 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_71
timestamp 1581321262
transform 1 0 5312 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_72
timestamp 1581321262
transform 1 0 4800 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_73
timestamp 1581321262
transform 1 0 4392 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_74
timestamp 1581321262
transform 1 0 3984 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_75
timestamp 1581321262
transform 1 0 3576 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_76
timestamp 1581321262
transform 1 0 3064 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_77
timestamp 1581321262
transform 1 0 2656 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_78
timestamp 1581321262
transform 1 0 2248 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_79
timestamp 1581321262
transform 1 0 1840 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_80
timestamp 1581321262
transform 1 0 1328 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_81
timestamp 1581321262
transform 1 0 920 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_82
timestamp 1581321262
transform 1 0 512 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_83
timestamp 1581321262
transform 1 0 104 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_84
timestamp 1581321262
transform 1 0 8476 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_85
timestamp 1581321262
transform 1 0 8272 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_86
timestamp 1581321262
transform 1 0 7660 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_87
timestamp 1581321262
transform 1 0 7456 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_88
timestamp 1581321262
transform 1 0 6740 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_89
timestamp 1581321262
transform 1 0 6536 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_90
timestamp 1581321262
transform 1 0 5924 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_91
timestamp 1581321262
transform 1 0 5720 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_92
timestamp 1581321262
transform 1 0 5004 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_93
timestamp 1581321262
transform 1 0 4800 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_94
timestamp 1581321262
transform 1 0 4188 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_95
timestamp 1581321262
transform 1 0 3984 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_96
timestamp 1581321262
transform 1 0 3268 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_97
timestamp 1581321262
transform 1 0 3064 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_98
timestamp 1581321262
transform 1 0 2452 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_99
timestamp 1581321262
transform 1 0 2248 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_100
timestamp 1581321262
transform 1 0 1532 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_101
timestamp 1581321262
transform 1 0 1328 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_102
timestamp 1581321262
transform 1 0 716 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_103
timestamp 1581321262
transform 1 0 512 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_104
timestamp 1581321262
transform 1 0 8988 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_105
timestamp 1581321262
transform 1 0 8784 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_106
timestamp 1581321262
transform 1 0 8068 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_107
timestamp 1581321262
transform 1 0 7864 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_108
timestamp 1581321262
transform 1 0 7252 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_109
timestamp 1581321262
transform 1 0 7048 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_110
timestamp 1581321262
transform 1 0 6332 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_111
timestamp 1581321262
transform 1 0 6128 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_112
timestamp 1581321262
transform 1 0 5516 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_113
timestamp 1581321262
transform 1 0 5312 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_114
timestamp 1581321262
transform 1 0 4596 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_115
timestamp 1581321262
transform 1 0 4392 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_116
timestamp 1581321262
transform 1 0 3780 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_117
timestamp 1581321262
transform 1 0 3576 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_118
timestamp 1581321262
transform 1 0 2860 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_119
timestamp 1581321262
transform 1 0 2656 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_120
timestamp 1581321262
transform 1 0 2044 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_121
timestamp 1581321262
transform 1 0 1840 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_122
timestamp 1581321262
transform 1 0 1124 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_123
timestamp 1581321262
transform 1 0 920 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_124
timestamp 1581321262
transform 1 0 308 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_125
timestamp 1581321262
transform 1 0 104 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_126
timestamp 1581321262
transform 1 0 8476 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_127
timestamp 1581321262
transform 1 0 8272 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_128
timestamp 1581321262
transform 1 0 8068 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_129
timestamp 1581321262
transform 1 0 7864 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_130
timestamp 1581321262
transform 1 0 6740 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_131
timestamp 1581321262
transform 1 0 6536 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_132
timestamp 1581321262
transform 1 0 6332 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_133
timestamp 1581321262
transform 1 0 6128 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_134
timestamp 1581321262
transform 1 0 5004 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_135
timestamp 1581321262
transform 1 0 4800 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_136
timestamp 1581321262
transform 1 0 4596 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_137
timestamp 1581321262
transform 1 0 4392 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_138
timestamp 1581321262
transform 1 0 3268 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_139
timestamp 1581321262
transform 1 0 3064 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_140
timestamp 1581321262
transform 1 0 2860 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_141
timestamp 1581321262
transform 1 0 2656 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_142
timestamp 1581321262
transform 1 0 1532 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_143
timestamp 1581321262
transform 1 0 1328 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_144
timestamp 1581321262
transform 1 0 1124 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_145
timestamp 1581321262
transform 1 0 920 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_146
timestamp 1581321262
transform 1 0 8988 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_147
timestamp 1581321262
transform 1 0 8784 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_148
timestamp 1581321262
transform 1 0 7660 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_149
timestamp 1581321262
transform 1 0 7456 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_150
timestamp 1581321262
transform 1 0 7252 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_151
timestamp 1581321262
transform 1 0 7048 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_152
timestamp 1581321262
transform 1 0 5924 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_153
timestamp 1581321262
transform 1 0 5720 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_154
timestamp 1581321262
transform 1 0 5516 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_155
timestamp 1581321262
transform 1 0 5312 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_156
timestamp 1581321262
transform 1 0 4188 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_157
timestamp 1581321262
transform 1 0 3984 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_158
timestamp 1581321262
transform 1 0 3780 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_159
timestamp 1581321262
transform 1 0 3576 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_160
timestamp 1581321262
transform 1 0 2452 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_161
timestamp 1581321262
transform 1 0 2248 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_162
timestamp 1581321262
transform 1 0 2044 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_163
timestamp 1581321262
transform 1 0 1840 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_164
timestamp 1581321262
transform 1 0 716 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_165
timestamp 1581321262
transform 1 0 512 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_166
timestamp 1581321262
transform 1 0 308 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_167
timestamp 1581321262
transform 1 0 104 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_168
timestamp 1581321262
transform 1 0 8988 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_169
timestamp 1581321262
transform 1 0 8784 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_170
timestamp 1581321262
transform 1 0 6740 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_171
timestamp 1581321262
transform 1 0 6536 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_172
timestamp 1581321262
transform 1 0 6332 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_173
timestamp 1581321262
transform 1 0 6128 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_174
timestamp 1581321262
transform 1 0 5924 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_175
timestamp 1581321262
transform 1 0 5720 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_176
timestamp 1581321262
transform 1 0 5516 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_177
timestamp 1581321262
transform 1 0 5312 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_178
timestamp 1581321262
transform 1 0 3268 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_179
timestamp 1581321262
transform 1 0 3064 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_180
timestamp 1581321262
transform 1 0 2860 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_181
timestamp 1581321262
transform 1 0 2656 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_182
timestamp 1581321262
transform 1 0 2452 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_183
timestamp 1581321262
transform 1 0 2248 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_184
timestamp 1581321262
transform 1 0 2044 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_185
timestamp 1581321262
transform 1 0 1840 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_186
timestamp 1581321262
transform 1 0 8476 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_187
timestamp 1581321262
transform 1 0 8272 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_188
timestamp 1581321262
transform 1 0 8068 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_189
timestamp 1581321262
transform 1 0 7864 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_190
timestamp 1581321262
transform 1 0 7660 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_191
timestamp 1581321262
transform 1 0 7456 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_192
timestamp 1581321262
transform 1 0 7252 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_193
timestamp 1581321262
transform 1 0 7048 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_194
timestamp 1581321262
transform 1 0 5004 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_195
timestamp 1581321262
transform 1 0 4800 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_196
timestamp 1581321262
transform 1 0 4596 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_197
timestamp 1581321262
transform 1 0 4392 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_198
timestamp 1581321262
transform 1 0 4188 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_199
timestamp 1581321262
transform 1 0 3984 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_200
timestamp 1581321262
transform 1 0 3780 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_201
timestamp 1581321262
transform 1 0 3576 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_202
timestamp 1581321262
transform 1 0 1532 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_203
timestamp 1581321262
transform 1 0 1328 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_204
timestamp 1581321262
transform 1 0 1124 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_205
timestamp 1581321262
transform 1 0 920 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_206
timestamp 1581321262
transform 1 0 716 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_207
timestamp 1581321262
transform 1 0 512 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_208
timestamp 1581321262
transform 1 0 308 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_209
timestamp 1581321262
transform 1 0 104 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_210
timestamp 1581321262
transform 1 0 6740 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_211
timestamp 1581321262
transform 1 0 6536 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_212
timestamp 1581321262
transform 1 0 6332 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_213
timestamp 1581321262
transform 1 0 6128 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_214
timestamp 1581321262
transform 1 0 5924 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_215
timestamp 1581321262
transform 1 0 5720 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_216
timestamp 1581321262
transform 1 0 5516 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_217
timestamp 1581321262
transform 1 0 5312 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_218
timestamp 1581321262
transform 1 0 5004 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_219
timestamp 1581321262
transform 1 0 4800 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_220
timestamp 1581321262
transform 1 0 4596 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_221
timestamp 1581321262
transform 1 0 4392 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_222
timestamp 1581321262
transform 1 0 4188 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_223
timestamp 1581321262
transform 1 0 3984 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_224
timestamp 1581321262
transform 1 0 3780 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_225
timestamp 1581321262
transform 1 0 3576 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_226
timestamp 1581321262
transform 1 0 8988 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_227
timestamp 1581321262
transform 1 0 8784 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_228
timestamp 1581321262
transform 1 0 8476 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_229
timestamp 1581321262
transform 1 0 8272 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_230
timestamp 1581321262
transform 1 0 8068 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_231
timestamp 1581321262
transform 1 0 7864 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_232
timestamp 1581321262
transform 1 0 7660 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_233
timestamp 1581321262
transform 1 0 7456 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_234
timestamp 1581321262
transform 1 0 7252 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_235
timestamp 1581321262
transform 1 0 7048 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_236
timestamp 1581321262
transform 1 0 3268 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_237
timestamp 1581321262
transform 1 0 3064 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_238
timestamp 1581321262
transform 1 0 2860 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_239
timestamp 1581321262
transform 1 0 2656 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_240
timestamp 1581321262
transform 1 0 2452 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_241
timestamp 1581321262
transform 1 0 2248 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_242
timestamp 1581321262
transform 1 0 2044 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_243
timestamp 1581321262
transform 1 0 1840 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_244
timestamp 1581321262
transform 1 0 1532 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_245
timestamp 1581321262
transform 1 0 1328 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_246
timestamp 1581321262
transform 1 0 1124 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_247
timestamp 1581321262
transform 1 0 920 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_248
timestamp 1581321262
transform 1 0 716 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_249
timestamp 1581321262
transform 1 0 512 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_250
timestamp 1581321262
transform 1 0 308 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_251
timestamp 1581321262
transform 1 0 104 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_252
timestamp 1581321262
transform 1 0 8988 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_253
timestamp 1581321262
transform 1 0 8784 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_254
timestamp 1581321262
transform 1 0 8476 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_255
timestamp 1581321262
transform 1 0 8272 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_256
timestamp 1581321262
transform 1 0 8068 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_257
timestamp 1581321262
transform 1 0 7864 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_258
timestamp 1581321262
transform 1 0 7660 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_259
timestamp 1581321262
transform 1 0 7456 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_260
timestamp 1581321262
transform 1 0 7252 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_261
timestamp 1581321262
transform 1 0 7048 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_262
timestamp 1581321262
transform 1 0 6740 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_263
timestamp 1581321262
transform 1 0 6536 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_264
timestamp 1581321262
transform 1 0 6332 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_265
timestamp 1581321262
transform 1 0 6128 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_266
timestamp 1581321262
transform 1 0 5924 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_267
timestamp 1581321262
transform 1 0 5720 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_268
timestamp 1581321262
transform 1 0 5516 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_269
timestamp 1581321262
transform 1 0 5312 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_270
timestamp 1581321262
transform 1 0 5004 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_271
timestamp 1581321262
transform 1 0 4800 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_272
timestamp 1581321262
transform 1 0 4596 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_273
timestamp 1581321262
transform 1 0 4392 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_274
timestamp 1581321262
transform 1 0 4188 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_275
timestamp 1581321262
transform 1 0 3984 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_276
timestamp 1581321262
transform 1 0 3780 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_277
timestamp 1581321262
transform 1 0 3576 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_278
timestamp 1581321262
transform 1 0 3268 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_279
timestamp 1581321262
transform 1 0 3064 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_280
timestamp 1581321262
transform 1 0 2860 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_281
timestamp 1581321262
transform 1 0 2656 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_282
timestamp 1581321262
transform 1 0 2452 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_283
timestamp 1581321262
transform 1 0 2248 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_284
timestamp 1581321262
transform 1 0 2044 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_285
timestamp 1581321262
transform 1 0 1840 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_286
timestamp 1581321262
transform 1 0 1532 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_287
timestamp 1581321262
transform 1 0 1328 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_288
timestamp 1581321262
transform 1 0 1124 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_289
timestamp 1581321262
transform 1 0 920 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_290
timestamp 1581321262
transform 1 0 716 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_291
timestamp 1581321262
transform 1 0 512 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_292
timestamp 1581321262
transform 1 0 308 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_293
timestamp 1581321262
transform 1 0 104 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_0
timestamp 1581321262
transform 1 0 8784 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1
timestamp 1581321262
transform 1 0 8272 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_2
timestamp 1581321262
transform 1 0 7864 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_3
timestamp 1581321262
transform 1 0 7456 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_4
timestamp 1581321262
transform 1 0 7048 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_5
timestamp 1581321262
transform 1 0 6536 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_6
timestamp 1581321262
transform 1 0 6128 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_7
timestamp 1581321262
transform 1 0 5720 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_8
timestamp 1581321262
transform 1 0 5312 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_9
timestamp 1581321262
transform 1 0 4800 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_10
timestamp 1581321262
transform 1 0 4392 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_11
timestamp 1581321262
transform 1 0 3984 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_12
timestamp 1581321262
transform 1 0 3576 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_13
timestamp 1581321262
transform 1 0 3064 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_14
timestamp 1581321262
transform 1 0 2656 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_15
timestamp 1581321262
transform 1 0 2248 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_16
timestamp 1581321262
transform 1 0 1840 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_17
timestamp 1581321262
transform 1 0 1328 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_18
timestamp 1581321262
transform 1 0 920 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_19
timestamp 1581321262
transform 1 0 512 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_20
timestamp 1581321262
transform 1 0 104 0 1 3117
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_21
timestamp 1581321262
transform 1 0 8988 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_22
timestamp 1581321262
transform 1 0 8476 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_23
timestamp 1581321262
transform 1 0 8068 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_24
timestamp 1581321262
transform 1 0 7660 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_25
timestamp 1581321262
transform 1 0 7252 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_26
timestamp 1581321262
transform 1 0 6740 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_27
timestamp 1581321262
transform 1 0 6332 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_28
timestamp 1581321262
transform 1 0 5924 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_29
timestamp 1581321262
transform 1 0 5516 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_30
timestamp 1581321262
transform 1 0 5004 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_31
timestamp 1581321262
transform 1 0 4596 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_32
timestamp 1581321262
transform 1 0 4188 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_33
timestamp 1581321262
transform 1 0 3780 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_34
timestamp 1581321262
transform 1 0 3268 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_35
timestamp 1581321262
transform 1 0 2860 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_36
timestamp 1581321262
transform 1 0 2452 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_37
timestamp 1581321262
transform 1 0 2044 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_38
timestamp 1581321262
transform 1 0 1532 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_39
timestamp 1581321262
transform 1 0 1124 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_40
timestamp 1581321262
transform 1 0 716 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_41
timestamp 1581321262
transform 1 0 308 0 1 2913
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_42
timestamp 1581321262
transform 1 0 8988 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_43
timestamp 1581321262
transform 1 0 8784 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_44
timestamp 1581321262
transform 1 0 8068 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_45
timestamp 1581321262
transform 1 0 7864 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_46
timestamp 1581321262
transform 1 0 7252 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_47
timestamp 1581321262
transform 1 0 7048 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_48
timestamp 1581321262
transform 1 0 6332 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_49
timestamp 1581321262
transform 1 0 6128 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_50
timestamp 1581321262
transform 1 0 5516 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_51
timestamp 1581321262
transform 1 0 5312 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_52
timestamp 1581321262
transform 1 0 4596 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_53
timestamp 1581321262
transform 1 0 4392 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_54
timestamp 1581321262
transform 1 0 3780 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_55
timestamp 1581321262
transform 1 0 3576 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_56
timestamp 1581321262
transform 1 0 2860 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_57
timestamp 1581321262
transform 1 0 2656 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_58
timestamp 1581321262
transform 1 0 2044 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_59
timestamp 1581321262
transform 1 0 1840 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_60
timestamp 1581321262
transform 1 0 1124 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_61
timestamp 1581321262
transform 1 0 920 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_62
timestamp 1581321262
transform 1 0 308 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_63
timestamp 1581321262
transform 1 0 104 0 1 2709
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_64
timestamp 1581321262
transform 1 0 8476 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_65
timestamp 1581321262
transform 1 0 8272 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_66
timestamp 1581321262
transform 1 0 7660 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_67
timestamp 1581321262
transform 1 0 7456 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_68
timestamp 1581321262
transform 1 0 6740 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_69
timestamp 1581321262
transform 1 0 6536 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_70
timestamp 1581321262
transform 1 0 5924 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_71
timestamp 1581321262
transform 1 0 5720 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_72
timestamp 1581321262
transform 1 0 5004 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_73
timestamp 1581321262
transform 1 0 4800 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_74
timestamp 1581321262
transform 1 0 4188 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_75
timestamp 1581321262
transform 1 0 3984 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_76
timestamp 1581321262
transform 1 0 3268 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_77
timestamp 1581321262
transform 1 0 3064 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_78
timestamp 1581321262
transform 1 0 2452 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_79
timestamp 1581321262
transform 1 0 2248 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_80
timestamp 1581321262
transform 1 0 1532 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_81
timestamp 1581321262
transform 1 0 1328 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_82
timestamp 1581321262
transform 1 0 716 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_83
timestamp 1581321262
transform 1 0 512 0 1 2505
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_84
timestamp 1581321262
transform 1 0 8988 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_85
timestamp 1581321262
transform 1 0 8784 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_86
timestamp 1581321262
transform 1 0 7660 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_87
timestamp 1581321262
transform 1 0 7456 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_88
timestamp 1581321262
transform 1 0 7252 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_89
timestamp 1581321262
transform 1 0 7048 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_90
timestamp 1581321262
transform 1 0 5924 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_91
timestamp 1581321262
transform 1 0 5720 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_92
timestamp 1581321262
transform 1 0 5516 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_93
timestamp 1581321262
transform 1 0 5312 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_94
timestamp 1581321262
transform 1 0 4188 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_95
timestamp 1581321262
transform 1 0 3984 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_96
timestamp 1581321262
transform 1 0 3780 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_97
timestamp 1581321262
transform 1 0 3576 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_98
timestamp 1581321262
transform 1 0 2452 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_99
timestamp 1581321262
transform 1 0 2248 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_100
timestamp 1581321262
transform 1 0 2044 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_101
timestamp 1581321262
transform 1 0 1840 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_102
timestamp 1581321262
transform 1 0 716 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_103
timestamp 1581321262
transform 1 0 512 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_104
timestamp 1581321262
transform 1 0 308 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_105
timestamp 1581321262
transform 1 0 104 0 1 2301
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_106
timestamp 1581321262
transform 1 0 8476 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_107
timestamp 1581321262
transform 1 0 8272 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_108
timestamp 1581321262
transform 1 0 8068 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_109
timestamp 1581321262
transform 1 0 7864 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_110
timestamp 1581321262
transform 1 0 6740 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_111
timestamp 1581321262
transform 1 0 6536 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_112
timestamp 1581321262
transform 1 0 6332 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_113
timestamp 1581321262
transform 1 0 6128 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_114
timestamp 1581321262
transform 1 0 5004 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_115
timestamp 1581321262
transform 1 0 4800 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_116
timestamp 1581321262
transform 1 0 4596 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_117
timestamp 1581321262
transform 1 0 4392 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_118
timestamp 1581321262
transform 1 0 3268 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_119
timestamp 1581321262
transform 1 0 3064 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_120
timestamp 1581321262
transform 1 0 2860 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_121
timestamp 1581321262
transform 1 0 2656 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_122
timestamp 1581321262
transform 1 0 1532 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_123
timestamp 1581321262
transform 1 0 1328 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_124
timestamp 1581321262
transform 1 0 1124 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_125
timestamp 1581321262
transform 1 0 920 0 1 2097
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_126
timestamp 1581321262
transform 1 0 8476 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_127
timestamp 1581321262
transform 1 0 8272 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_128
timestamp 1581321262
transform 1 0 8068 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_129
timestamp 1581321262
transform 1 0 7864 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_130
timestamp 1581321262
transform 1 0 7660 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_131
timestamp 1581321262
transform 1 0 7456 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_132
timestamp 1581321262
transform 1 0 7252 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_133
timestamp 1581321262
transform 1 0 7048 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_134
timestamp 1581321262
transform 1 0 5004 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_135
timestamp 1581321262
transform 1 0 4800 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_136
timestamp 1581321262
transform 1 0 4596 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_137
timestamp 1581321262
transform 1 0 4392 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_138
timestamp 1581321262
transform 1 0 4188 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_139
timestamp 1581321262
transform 1 0 3984 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_140
timestamp 1581321262
transform 1 0 3780 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_141
timestamp 1581321262
transform 1 0 3576 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_142
timestamp 1581321262
transform 1 0 1532 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_143
timestamp 1581321262
transform 1 0 1328 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_144
timestamp 1581321262
transform 1 0 1124 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_145
timestamp 1581321262
transform 1 0 920 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_146
timestamp 1581321262
transform 1 0 716 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_147
timestamp 1581321262
transform 1 0 512 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_148
timestamp 1581321262
transform 1 0 308 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_149
timestamp 1581321262
transform 1 0 104 0 1 1893
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_150
timestamp 1581321262
transform 1 0 8988 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_151
timestamp 1581321262
transform 1 0 8784 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_152
timestamp 1581321262
transform 1 0 6740 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_153
timestamp 1581321262
transform 1 0 6536 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_154
timestamp 1581321262
transform 1 0 6332 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_155
timestamp 1581321262
transform 1 0 6128 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_156
timestamp 1581321262
transform 1 0 5924 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_157
timestamp 1581321262
transform 1 0 5720 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_158
timestamp 1581321262
transform 1 0 5516 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_159
timestamp 1581321262
transform 1 0 5312 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_160
timestamp 1581321262
transform 1 0 3268 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_161
timestamp 1581321262
transform 1 0 3064 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_162
timestamp 1581321262
transform 1 0 2860 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_163
timestamp 1581321262
transform 1 0 2656 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_164
timestamp 1581321262
transform 1 0 2452 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_165
timestamp 1581321262
transform 1 0 2248 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_166
timestamp 1581321262
transform 1 0 2044 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_167
timestamp 1581321262
transform 1 0 1840 0 1 1689
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_168
timestamp 1581321262
transform 1 0 8988 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_169
timestamp 1581321262
transform 1 0 8784 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_170
timestamp 1581321262
transform 1 0 8476 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_171
timestamp 1581321262
transform 1 0 8272 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_172
timestamp 1581321262
transform 1 0 8068 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_173
timestamp 1581321262
transform 1 0 7864 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_174
timestamp 1581321262
transform 1 0 7660 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_175
timestamp 1581321262
transform 1 0 7456 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_176
timestamp 1581321262
transform 1 0 7252 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_177
timestamp 1581321262
transform 1 0 7048 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_178
timestamp 1581321262
transform 1 0 3268 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_179
timestamp 1581321262
transform 1 0 3064 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_180
timestamp 1581321262
transform 1 0 2860 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_181
timestamp 1581321262
transform 1 0 2656 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_182
timestamp 1581321262
transform 1 0 2452 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_183
timestamp 1581321262
transform 1 0 2248 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_184
timestamp 1581321262
transform 1 0 2044 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_185
timestamp 1581321262
transform 1 0 1840 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_186
timestamp 1581321262
transform 1 0 1532 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_187
timestamp 1581321262
transform 1 0 1328 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_188
timestamp 1581321262
transform 1 0 1124 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_189
timestamp 1581321262
transform 1 0 920 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_190
timestamp 1581321262
transform 1 0 716 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_191
timestamp 1581321262
transform 1 0 512 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_192
timestamp 1581321262
transform 1 0 308 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_193
timestamp 1581321262
transform 1 0 104 0 1 1485
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_194
timestamp 1581321262
transform 1 0 6740 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_195
timestamp 1581321262
transform 1 0 6536 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_196
timestamp 1581321262
transform 1 0 6332 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_197
timestamp 1581321262
transform 1 0 6128 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_198
timestamp 1581321262
transform 1 0 5924 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_199
timestamp 1581321262
transform 1 0 5720 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_200
timestamp 1581321262
transform 1 0 5516 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_201
timestamp 1581321262
transform 1 0 5312 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_202
timestamp 1581321262
transform 1 0 5004 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_203
timestamp 1581321262
transform 1 0 4800 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_204
timestamp 1581321262
transform 1 0 4596 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_205
timestamp 1581321262
transform 1 0 4392 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_206
timestamp 1581321262
transform 1 0 4188 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_207
timestamp 1581321262
transform 1 0 3984 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_208
timestamp 1581321262
transform 1 0 3780 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_209
timestamp 1581321262
transform 1 0 3576 0 1 1281
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_210
timestamp 1581321262
transform 1 0 6740 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_211
timestamp 1581321262
transform 1 0 6536 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_212
timestamp 1581321262
transform 1 0 6332 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_213
timestamp 1581321262
transform 1 0 6128 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_214
timestamp 1581321262
transform 1 0 5924 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_215
timestamp 1581321262
transform 1 0 5720 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_216
timestamp 1581321262
transform 1 0 5516 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_217
timestamp 1581321262
transform 1 0 5312 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_218
timestamp 1581321262
transform 1 0 5004 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_219
timestamp 1581321262
transform 1 0 4800 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_220
timestamp 1581321262
transform 1 0 4596 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_221
timestamp 1581321262
transform 1 0 4392 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_222
timestamp 1581321262
transform 1 0 4188 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_223
timestamp 1581321262
transform 1 0 3984 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_224
timestamp 1581321262
transform 1 0 3780 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_225
timestamp 1581321262
transform 1 0 3576 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_226
timestamp 1581321262
transform 1 0 3268 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_227
timestamp 1581321262
transform 1 0 3064 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_228
timestamp 1581321262
transform 1 0 2860 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_229
timestamp 1581321262
transform 1 0 2656 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_230
timestamp 1581321262
transform 1 0 2452 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_231
timestamp 1581321262
transform 1 0 2248 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_232
timestamp 1581321262
transform 1 0 2044 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_233
timestamp 1581321262
transform 1 0 1840 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_234
timestamp 1581321262
transform 1 0 1532 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_235
timestamp 1581321262
transform 1 0 1328 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_236
timestamp 1581321262
transform 1 0 1124 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_237
timestamp 1581321262
transform 1 0 920 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_238
timestamp 1581321262
transform 1 0 716 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_239
timestamp 1581321262
transform 1 0 512 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_240
timestamp 1581321262
transform 1 0 308 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_241
timestamp 1581321262
transform 1 0 104 0 1 1077
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_242
timestamp 1581321262
transform 1 0 8988 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_243
timestamp 1581321262
transform 1 0 8784 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_244
timestamp 1581321262
transform 1 0 8476 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_245
timestamp 1581321262
transform 1 0 8272 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_246
timestamp 1581321262
transform 1 0 8068 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_247
timestamp 1581321262
transform 1 0 7864 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_248
timestamp 1581321262
transform 1 0 7660 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_249
timestamp 1581321262
transform 1 0 7456 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_250
timestamp 1581321262
transform 1 0 7252 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_251
timestamp 1581321262
transform 1 0 7048 0 1 873
box 0 -51 204 204
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_0
timestamp 1581321264
transform 1 0 9192 0 1 3117
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_1
timestamp 1581321264
transform 1 0 8680 0 1 3117
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_2
timestamp 1581321264
transform 1 0 6944 0 1 3117
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_3
timestamp 1581321264
transform 1 0 5208 0 1 3117
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_4
timestamp 1581321264
transform 1 0 3472 0 1 3117
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_5
timestamp 1581321264
transform 1 0 1736 0 1 3117
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_6
timestamp 1581321264
transform 1 0 0 0 1 3117
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_7
timestamp 1581321264
transform 1 0 9192 0 1 2913
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_8
timestamp 1581321264
transform 1 0 8680 0 1 2913
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_9
timestamp 1581321264
transform 1 0 6944 0 1 2913
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_10
timestamp 1581321264
transform 1 0 5208 0 1 2913
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_11
timestamp 1581321264
transform 1 0 3472 0 1 2913
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_12
timestamp 1581321264
transform 1 0 1736 0 1 2913
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_13
timestamp 1581321264
transform 1 0 0 0 1 2913
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_14
timestamp 1581321264
transform 1 0 9192 0 1 2709
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_15
timestamp 1581321264
transform 1 0 8680 0 1 2709
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_16
timestamp 1581321264
transform 1 0 6944 0 1 2709
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_17
timestamp 1581321264
transform 1 0 5208 0 1 2709
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_18
timestamp 1581321264
transform 1 0 3472 0 1 2709
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_19
timestamp 1581321264
transform 1 0 1736 0 1 2709
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_20
timestamp 1581321264
transform 1 0 0 0 1 2709
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_21
timestamp 1581321264
transform 1 0 9192 0 1 2505
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_22
timestamp 1581321264
transform 1 0 8680 0 1 2505
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_23
timestamp 1581321264
transform 1 0 6944 0 1 2505
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_24
timestamp 1581321264
transform 1 0 5208 0 1 2505
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_25
timestamp 1581321264
transform 1 0 3472 0 1 2505
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_26
timestamp 1581321264
transform 1 0 1736 0 1 2505
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_27
timestamp 1581321264
transform 1 0 0 0 1 2505
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_28
timestamp 1581321264
transform 1 0 9192 0 1 2301
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_29
timestamp 1581321264
transform 1 0 8680 0 1 2301
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_30
timestamp 1581321264
transform 1 0 6944 0 1 2301
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_31
timestamp 1581321264
transform 1 0 5208 0 1 2301
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_32
timestamp 1581321264
transform 1 0 3472 0 1 2301
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_33
timestamp 1581321264
transform 1 0 1736 0 1 2301
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_34
timestamp 1581321264
transform 1 0 0 0 1 2301
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_35
timestamp 1581321264
transform 1 0 9192 0 1 2097
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_36
timestamp 1581321264
transform 1 0 8680 0 1 2097
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_37
timestamp 1581321264
transform 1 0 6944 0 1 2097
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_38
timestamp 1581321264
transform 1 0 5208 0 1 2097
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_39
timestamp 1581321264
transform 1 0 3472 0 1 2097
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_40
timestamp 1581321264
transform 1 0 1736 0 1 2097
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_41
timestamp 1581321264
transform 1 0 0 0 1 2097
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_42
timestamp 1581321264
transform 1 0 9192 0 1 1893
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_43
timestamp 1581321264
transform 1 0 8680 0 1 1893
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_44
timestamp 1581321264
transform 1 0 6944 0 1 1893
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_45
timestamp 1581321264
transform 1 0 5208 0 1 1893
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_46
timestamp 1581321264
transform 1 0 3472 0 1 1893
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_47
timestamp 1581321264
transform 1 0 1736 0 1 1893
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_48
timestamp 1581321264
transform 1 0 0 0 1 1893
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_49
timestamp 1581321264
transform 1 0 9192 0 1 1689
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_50
timestamp 1581321264
transform 1 0 8680 0 1 1689
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_51
timestamp 1581321264
transform 1 0 6944 0 1 1689
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_52
timestamp 1581321264
transform 1 0 5208 0 1 1689
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_53
timestamp 1581321264
transform 1 0 3472 0 1 1689
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_54
timestamp 1581321264
transform 1 0 1736 0 1 1689
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_55
timestamp 1581321264
transform 1 0 0 0 1 1689
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_56
timestamp 1581321264
transform 1 0 9192 0 1 1485
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_57
timestamp 1581321264
transform 1 0 8680 0 1 1485
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_58
timestamp 1581321264
transform 1 0 6944 0 1 1485
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_59
timestamp 1581321264
transform 1 0 5208 0 1 1485
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_60
timestamp 1581321264
transform 1 0 3472 0 1 1485
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_61
timestamp 1581321264
transform 1 0 1736 0 1 1485
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_62
timestamp 1581321264
transform 1 0 0 0 1 1485
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_63
timestamp 1581321264
transform 1 0 9192 0 1 1281
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_64
timestamp 1581321264
transform 1 0 8680 0 1 1281
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_65
timestamp 1581321264
transform 1 0 6944 0 1 1281
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_66
timestamp 1581321264
transform 1 0 5208 0 1 1281
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_67
timestamp 1581321264
transform 1 0 3472 0 1 1281
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_68
timestamp 1581321264
transform 1 0 1736 0 1 1281
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_69
timestamp 1581321264
transform 1 0 0 0 1 1281
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_70
timestamp 1581321264
transform 1 0 9192 0 1 1077
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_71
timestamp 1581321264
transform 1 0 8680 0 1 1077
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_72
timestamp 1581321264
transform 1 0 6944 0 1 1077
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_73
timestamp 1581321264
transform 1 0 5208 0 1 1077
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_74
timestamp 1581321264
transform 1 0 3472 0 1 1077
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_75
timestamp 1581321264
transform 1 0 1736 0 1 1077
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_76
timestamp 1581321264
transform 1 0 0 0 1 1077
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_77
timestamp 1581321264
transform 1 0 9192 0 1 873
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_78
timestamp 1581321264
transform 1 0 8680 0 1 873
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_79
timestamp 1581321264
transform 1 0 6944 0 1 873
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_80
timestamp 1581321264
transform 1 0 5208 0 1 873
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_81
timestamp 1581321264
transform 1 0 3472 0 1 873
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_82
timestamp 1581321264
transform 1 0 1736 0 1 873
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_1  sky130_rom_krom_rom_poly_tap_1_83
timestamp 1581321264
transform 1 0 0 0 1 873
box -6 17 128 203
use sky130_rom_krom_rom_poly_tap_2  sky130_rom_krom_rom_poly_tap_2_0
timestamp 1581321264
transform 1 0 9192 0 1 3321
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_2  sky130_rom_krom_rom_poly_tap_2_1
timestamp 1581321264
transform 1 0 8680 0 1 3321
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_2  sky130_rom_krom_rom_poly_tap_2_2
timestamp 1581321264
transform 1 0 6944 0 1 3321
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_2  sky130_rom_krom_rom_poly_tap_2_3
timestamp 1581321264
transform 1 0 5208 0 1 3321
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_2  sky130_rom_krom_rom_poly_tap_2_4
timestamp 1581321264
transform 1 0 3472 0 1 3321
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_2  sky130_rom_krom_rom_poly_tap_2_5
timestamp 1581321264
transform 1 0 1736 0 1 3321
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap_2  sky130_rom_krom_rom_poly_tap_2_6
timestamp 1581321264
transform 1 0 0 0 1 3321
box 0 17 66 83
use sky130_rom_krom_rom_precharge_array_0  sky130_rom_krom_rom_precharge_array_0_0
timestamp 1581321264
transform 1 0 0 0 1 128
box 0 -212 9404 408
<< labels >>
rlabel metal2 s 61 368 89 396 4 precharge
port 3 nsew
rlabel metal2 s 19 909 47 937 4 wl_0_0
port 5 nsew
rlabel metal2 s 19 1113 47 1141 4 wl_0_1
port 7 nsew
rlabel metal2 s 19 1317 47 1345 4 wl_0_2
port 9 nsew
rlabel metal2 s 19 1521 47 1549 4 wl_0_3
port 11 nsew
rlabel metal2 s 19 1725 47 1753 4 wl_0_4
port 13 nsew
rlabel metal2 s 19 1929 47 1957 4 wl_0_5
port 15 nsew
rlabel metal2 s 19 2133 47 2161 4 wl_0_6
port 17 nsew
rlabel metal2 s 19 2337 47 2365 4 wl_0_7
port 19 nsew
rlabel metal2 s 19 2541 47 2569 4 wl_0_8
port 21 nsew
rlabel metal2 s 19 2745 47 2773 4 wl_0_9
port 23 nsew
rlabel metal2 s 19 2949 47 2977 4 wl_0_10
port 25 nsew
rlabel metal2 s 19 3153 47 3181 4 wl_0_11
port 27 nsew
rlabel metal1 s 232 -14 260 14 4 bl_0_0
port 29 nsew
rlabel metal1 s 436 -14 464 14 4 bl_0_1
port 31 nsew
rlabel metal1 s 640 -14 668 14 4 bl_0_2
port 33 nsew
rlabel metal1 s 844 -14 872 14 4 bl_0_3
port 35 nsew
rlabel metal1 s 1048 -14 1076 14 4 bl_0_4
port 37 nsew
rlabel metal1 s 1252 -14 1280 14 4 bl_0_5
port 39 nsew
rlabel metal1 s 1456 -14 1484 14 4 bl_0_6
port 41 nsew
rlabel metal1 s 1660 -14 1688 14 4 bl_0_7
port 43 nsew
rlabel metal1 s 1968 -14 1996 14 4 bl_0_8
port 45 nsew
rlabel metal1 s 2172 -14 2200 14 4 bl_0_9
port 47 nsew
rlabel metal1 s 2376 -14 2404 14 4 bl_0_10
port 49 nsew
rlabel metal1 s 2580 -14 2608 14 4 bl_0_11
port 51 nsew
rlabel metal1 s 2784 -14 2812 14 4 bl_0_12
port 53 nsew
rlabel metal1 s 2988 -14 3016 14 4 bl_0_13
port 55 nsew
rlabel metal1 s 3192 -14 3220 14 4 bl_0_14
port 57 nsew
rlabel metal1 s 3396 -14 3424 14 4 bl_0_15
port 59 nsew
rlabel metal1 s 3704 -14 3732 14 4 bl_0_16
port 61 nsew
rlabel metal1 s 3908 -14 3936 14 4 bl_0_17
port 63 nsew
rlabel metal1 s 4112 -14 4140 14 4 bl_0_18
port 65 nsew
rlabel metal1 s 4316 -14 4344 14 4 bl_0_19
port 67 nsew
rlabel metal1 s 4520 -14 4548 14 4 bl_0_20
port 69 nsew
rlabel metal1 s 4724 -14 4752 14 4 bl_0_21
port 71 nsew
rlabel metal1 s 4928 -14 4956 14 4 bl_0_22
port 73 nsew
rlabel metal1 s 5132 -14 5160 14 4 bl_0_23
port 75 nsew
rlabel metal1 s 5440 -14 5468 14 4 bl_0_24
port 77 nsew
rlabel metal1 s 5644 -14 5672 14 4 bl_0_25
port 79 nsew
rlabel metal1 s 5848 -14 5876 14 4 bl_0_26
port 81 nsew
rlabel metal1 s 6052 -14 6080 14 4 bl_0_27
port 83 nsew
rlabel metal1 s 6256 -14 6284 14 4 bl_0_28
port 85 nsew
rlabel metal1 s 6460 -14 6488 14 4 bl_0_29
port 87 nsew
rlabel metal1 s 6664 -14 6692 14 4 bl_0_30
port 89 nsew
rlabel metal1 s 6868 -14 6896 14 4 bl_0_31
port 91 nsew
rlabel metal1 s 7176 -14 7204 14 4 bl_0_32
port 93 nsew
rlabel metal1 s 7380 -14 7408 14 4 bl_0_33
port 95 nsew
rlabel metal1 s 7584 -14 7612 14 4 bl_0_34
port 97 nsew
rlabel metal1 s 7788 -14 7816 14 4 bl_0_35
port 99 nsew
rlabel metal1 s 7992 -14 8020 14 4 bl_0_36
port 101 nsew
rlabel metal1 s 8196 -14 8224 14 4 bl_0_37
port 103 nsew
rlabel metal1 s 8400 -14 8428 14 4 bl_0_38
port 105 nsew
rlabel metal1 s 8604 -14 8632 14 4 bl_0_39
port 107 nsew
rlabel metal1 s 8912 -14 8940 14 4 bl_0_40
port 109 nsew
rlabel metal1 s 9116 -14 9144 14 4 bl_0_41
port 111 nsew
rlabel metal1 s 9493 368 9521 396 4 precharge_r
port 113 nsew
rlabel metal3 s 3503 3468 3563 3528 4 gnd
port 115 nsew
rlabel metal3 s 6975 3468 7035 3528 4 gnd
port 115 nsew
rlabel metal3 s 31 3468 91 3528 4 gnd
port 115 nsew
rlabel metal3 s 5239 978 5299 1038 4 gnd
port 115 nsew
rlabel metal3 s 9223 3468 9283 3528 4 gnd
port 115 nsew
rlabel metal3 s 9223 978 9283 1038 4 gnd
port 115 nsew
rlabel metal3 s 3503 978 3563 1038 4 gnd
port 115 nsew
rlabel metal3 s 8711 978 8771 1038 4 gnd
port 115 nsew
rlabel metal3 s 5239 3468 5299 3528 4 gnd
port 115 nsew
rlabel metal3 s 6975 978 7035 1038 4 gnd
port 115 nsew
rlabel metal3 s 1767 3468 1827 3528 4 gnd
port 115 nsew
rlabel metal3 s 31 978 91 1038 4 gnd
port 115 nsew
rlabel metal3 s 8711 3468 8771 3528 4 gnd
port 115 nsew
rlabel metal3 s 1767 978 1827 1038 4 gnd
port 115 nsew
rlabel metal2 s 12 -32 40 32 4 vdd
port 117 nsew
<< properties >>
string FIXED_BBOX 0 0 9521 870
<< end >>
