magic
tech sky130A
magscale 1 2
timestamp 1581320207
<< checkpaint >>
rect -1296 -1277 3308 3946
<< nwell >>
rect -36 1261 2048 2686
<< locali >>
rect 0 2611 2012 2645
rect 64 1244 98 1310
rect 179 1272 449 1306
rect 551 1282 585 1289
rect 551 1248 925 1282
rect 1027 1232 1061 1265
rect 1027 1198 1401 1232
rect 1611 1198 1645 1232
rect 0 -17 2012 17
use sky130_rom_krom_pinv  sky130_rom_krom_pinv_0
timestamp 1581320207
transform 1 0 0 0 1 0
box -36 -17 404 2686
use sky130_rom_krom_pinv_0  sky130_rom_krom_pinv_0_0
timestamp 1581320207
transform 1 0 368 0 1 0
box -36 -17 512 2686
use sky130_rom_krom_pinv_1  sky130_rom_krom_pinv_1_0
timestamp 1581320207
transform 1 0 844 0 1 0
box -36 -17 512 2686
use sky130_rom_krom_pinv_2  sky130_rom_krom_pinv_2_0
timestamp 1581320207
transform 1 0 1320 0 1 0
box -36 -17 728 2686
<< labels >>
rlabel locali s 1628 1215 1628 1215 4 Z
port 1 nsew
rlabel locali s 81 1277 81 1277 4 A
port 2 nsew
rlabel locali s 1006 0 1006 0 4 gnd
port 3 nsew
rlabel locali s 1006 2628 1006 2628 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2012 2628
<< end >>
