magic
tech sky130A
magscale 1 2
timestamp 1581365163
<< checkpaint >>
rect -1260 -1260 1261 1261
<< end >>
