VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_rom_krom
   CLASS BLOCK ;
   SIZE 100.87 BY 79.67 ;
   SYMMETRY X Y R90 ;
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 6.86 -7.1 7.24 ;
      END
   END clk0
   PIN cs0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  12.645 -7.48 13.025 -7.1 ;
      END
   END cs0
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  17.825 -7.48 18.205 -7.1 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  19.93 -7.48 20.31 -7.1 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  21.97 -7.48 22.35 -7.1 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 27.54 -7.1 27.92 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 28.285 -7.1 28.665 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 28.975 -7.1 29.355 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 26.07 -7.1 26.45 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 29.665 -7.1 30.045 ;
      END
   END addr0[7]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  42.695 -7.48 43.075 -7.1 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  44.235 -7.48 44.615 -7.1 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  45.775 -7.48 46.155 -7.1 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  47.315 -7.48 47.695 -7.1 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  48.855 -7.48 49.235 -7.1 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  50.395 -7.48 50.775 -7.1 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  51.935 -7.48 52.315 -7.1 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  53.475 -7.48 53.855 -7.1 ;
      END
   END dout0[7]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  -7.48 -7.48 108.35 -5.74 ;
         LAYER met3 ;
         RECT  -7.48 85.41 108.35 87.15 ;
         LAYER met4 ;
         RECT  106.61 -7.48 108.35 87.15 ;
         LAYER met4 ;
         RECT  -7.48 -7.48 -5.74 87.15 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  -4.0 -4.0 -2.26 83.67 ;
         LAYER met3 ;
         RECT  -4.0 81.93 104.87 83.67 ;
         LAYER met3 ;
         RECT  -4.0 -4.0 104.87 -2.26 ;
         LAYER met4 ;
         RECT  103.13 -4.0 104.87 83.67 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 100.25 79.05 ;
   LAYER  met2 ;
      RECT  0.62 0.62 100.25 79.05 ;
   LAYER  met3 ;
      RECT  0.62 0.62 100.25 79.05 ;
   LAYER  met4 ;
      RECT  0.62 0.62 100.25 79.05 ;
   END
END    sky130_rom_krom
END    LIBRARY
