magic
tech sky130A
magscale 1 2
timestamp 1581320207
<< checkpaint >>
rect -1216 -1310 4918 1559
<< locali >>
rect 60 51 94 117
rect 1254 51 1288 101
rect 1194 17 1288 51
rect 1623 17 3640 51
<< metal1 >>
rect 222 0 250 204
rect 844 0 872 204
rect 1642 0 1670 204
rect 2890 0 2918 204
use sky130_rom_krom_pinv_dec_0  sky130_rom_krom_pinv_dec_0_0
timestamp 1581320207
transform 1 0 0 0 1 0
box 44 -50 1212 299
use sky130_rom_krom_pinv_dec_1  sky130_rom_krom_pinv_dec_1_0
timestamp 1581320207
transform 1 0 1194 0 1 0
box 44 -50 2464 299
<< labels >>
rlabel locali s 2631 34 2631 34 4 Z
port 2 nsew
rlabel locali s 77 84 77 84 4 A
port 3 nsew
rlabel metal1 s 2890 0 2918 204 4 vdd
port 5 nsew
rlabel metal1 s 844 0 872 204 4 vdd
port 5 nsew
rlabel metal1 s 1642 0 1670 204 4 gnd
port 7 nsew
rlabel metal1 s 222 0 250 204 4 gnd
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 3640 204
<< end >>
