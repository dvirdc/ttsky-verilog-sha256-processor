magic
tech sky130A
magscale 1 2
timestamp 1581398725
<< checkpaint >>
rect -1296 -1277 3716 3946
<< nwell >>
rect -36 1262 2456 2686
<< pwell >>
rect 28 159 2282 1077
rect 28 25 2386 159
<< scnmos >>
rect 114 51 144 1051
rect 222 51 252 1051
rect 330 51 360 1051
rect 438 51 468 1051
rect 546 51 576 1051
rect 654 51 684 1051
rect 762 51 792 1051
rect 870 51 900 1051
rect 978 51 1008 1051
rect 1086 51 1116 1051
rect 1194 51 1224 1051
rect 1302 51 1332 1051
rect 1410 51 1440 1051
rect 1518 51 1548 1051
rect 1626 51 1656 1051
rect 1734 51 1764 1051
rect 1842 51 1872 1051
rect 1950 51 1980 1051
rect 2058 51 2088 1051
rect 2166 51 2196 1051
<< scpmos >>
rect 114 1578 144 2578
rect 222 1578 252 2578
rect 330 1578 360 2578
rect 438 1578 468 2578
rect 546 1578 576 2578
rect 654 1578 684 2578
rect 762 1578 792 2578
rect 870 1578 900 2578
rect 978 1578 1008 2578
rect 1086 1578 1116 2578
rect 1194 1578 1224 2578
rect 1302 1578 1332 2578
rect 1410 1578 1440 2578
rect 1518 1578 1548 2578
rect 1626 1578 1656 2578
rect 1734 1578 1764 2578
rect 1842 1578 1872 2578
rect 1950 1578 1980 2578
rect 2058 1578 2088 2578
rect 2166 1578 2196 2578
<< ndiff >>
rect 54 568 114 1051
rect 54 534 62 568
rect 96 534 114 568
rect 54 51 114 534
rect 144 568 222 1051
rect 144 534 166 568
rect 200 534 222 568
rect 144 51 222 534
rect 252 568 330 1051
rect 252 534 274 568
rect 308 534 330 568
rect 252 51 330 534
rect 360 568 438 1051
rect 360 534 382 568
rect 416 534 438 568
rect 360 51 438 534
rect 468 568 546 1051
rect 468 534 490 568
rect 524 534 546 568
rect 468 51 546 534
rect 576 568 654 1051
rect 576 534 598 568
rect 632 534 654 568
rect 576 51 654 534
rect 684 568 762 1051
rect 684 534 706 568
rect 740 534 762 568
rect 684 51 762 534
rect 792 568 870 1051
rect 792 534 814 568
rect 848 534 870 568
rect 792 51 870 534
rect 900 568 978 1051
rect 900 534 922 568
rect 956 534 978 568
rect 900 51 978 534
rect 1008 568 1086 1051
rect 1008 534 1030 568
rect 1064 534 1086 568
rect 1008 51 1086 534
rect 1116 568 1194 1051
rect 1116 534 1138 568
rect 1172 534 1194 568
rect 1116 51 1194 534
rect 1224 568 1302 1051
rect 1224 534 1246 568
rect 1280 534 1302 568
rect 1224 51 1302 534
rect 1332 568 1410 1051
rect 1332 534 1354 568
rect 1388 534 1410 568
rect 1332 51 1410 534
rect 1440 568 1518 1051
rect 1440 534 1462 568
rect 1496 534 1518 568
rect 1440 51 1518 534
rect 1548 568 1626 1051
rect 1548 534 1570 568
rect 1604 534 1626 568
rect 1548 51 1626 534
rect 1656 568 1734 1051
rect 1656 534 1678 568
rect 1712 534 1734 568
rect 1656 51 1734 534
rect 1764 568 1842 1051
rect 1764 534 1786 568
rect 1820 534 1842 568
rect 1764 51 1842 534
rect 1872 568 1950 1051
rect 1872 534 1894 568
rect 1928 534 1950 568
rect 1872 51 1950 534
rect 1980 568 2058 1051
rect 1980 534 2002 568
rect 2036 534 2058 568
rect 1980 51 2058 534
rect 2088 568 2166 1051
rect 2088 534 2110 568
rect 2144 534 2166 568
rect 2088 51 2166 534
rect 2196 568 2256 1051
rect 2196 534 2214 568
rect 2248 534 2256 568
rect 2196 51 2256 534
<< pdiff >>
rect 54 2095 114 2578
rect 54 2061 62 2095
rect 96 2061 114 2095
rect 54 1578 114 2061
rect 144 2095 222 2578
rect 144 2061 166 2095
rect 200 2061 222 2095
rect 144 1578 222 2061
rect 252 2095 330 2578
rect 252 2061 274 2095
rect 308 2061 330 2095
rect 252 1578 330 2061
rect 360 2095 438 2578
rect 360 2061 382 2095
rect 416 2061 438 2095
rect 360 1578 438 2061
rect 468 2095 546 2578
rect 468 2061 490 2095
rect 524 2061 546 2095
rect 468 1578 546 2061
rect 576 2095 654 2578
rect 576 2061 598 2095
rect 632 2061 654 2095
rect 576 1578 654 2061
rect 684 2095 762 2578
rect 684 2061 706 2095
rect 740 2061 762 2095
rect 684 1578 762 2061
rect 792 2095 870 2578
rect 792 2061 814 2095
rect 848 2061 870 2095
rect 792 1578 870 2061
rect 900 2095 978 2578
rect 900 2061 922 2095
rect 956 2061 978 2095
rect 900 1578 978 2061
rect 1008 2095 1086 2578
rect 1008 2061 1030 2095
rect 1064 2061 1086 2095
rect 1008 1578 1086 2061
rect 1116 2095 1194 2578
rect 1116 2061 1138 2095
rect 1172 2061 1194 2095
rect 1116 1578 1194 2061
rect 1224 2095 1302 2578
rect 1224 2061 1246 2095
rect 1280 2061 1302 2095
rect 1224 1578 1302 2061
rect 1332 2095 1410 2578
rect 1332 2061 1354 2095
rect 1388 2061 1410 2095
rect 1332 1578 1410 2061
rect 1440 2095 1518 2578
rect 1440 2061 1462 2095
rect 1496 2061 1518 2095
rect 1440 1578 1518 2061
rect 1548 2095 1626 2578
rect 1548 2061 1570 2095
rect 1604 2061 1626 2095
rect 1548 1578 1626 2061
rect 1656 2095 1734 2578
rect 1656 2061 1678 2095
rect 1712 2061 1734 2095
rect 1656 1578 1734 2061
rect 1764 2095 1842 2578
rect 1764 2061 1786 2095
rect 1820 2061 1842 2095
rect 1764 1578 1842 2061
rect 1872 2095 1950 2578
rect 1872 2061 1894 2095
rect 1928 2061 1950 2095
rect 1872 1578 1950 2061
rect 1980 2095 2058 2578
rect 1980 2061 2002 2095
rect 2036 2061 2058 2095
rect 1980 1578 2058 2061
rect 2088 2095 2166 2578
rect 2088 2061 2110 2095
rect 2144 2061 2166 2095
rect 2088 1578 2166 2061
rect 2196 2095 2256 2578
rect 2196 2061 2214 2095
rect 2248 2061 2256 2095
rect 2196 1578 2256 2061
<< ndiffc >>
rect 62 534 96 568
rect 166 534 200 568
rect 274 534 308 568
rect 382 534 416 568
rect 490 534 524 568
rect 598 534 632 568
rect 706 534 740 568
rect 814 534 848 568
rect 922 534 956 568
rect 1030 534 1064 568
rect 1138 534 1172 568
rect 1246 534 1280 568
rect 1354 534 1388 568
rect 1462 534 1496 568
rect 1570 534 1604 568
rect 1678 534 1712 568
rect 1786 534 1820 568
rect 1894 534 1928 568
rect 2002 534 2036 568
rect 2110 534 2144 568
rect 2214 534 2248 568
<< pdiffc >>
rect 62 2061 96 2095
rect 166 2061 200 2095
rect 274 2061 308 2095
rect 382 2061 416 2095
rect 490 2061 524 2095
rect 598 2061 632 2095
rect 706 2061 740 2095
rect 814 2061 848 2095
rect 922 2061 956 2095
rect 1030 2061 1064 2095
rect 1138 2061 1172 2095
rect 1246 2061 1280 2095
rect 1354 2061 1388 2095
rect 1462 2061 1496 2095
rect 1570 2061 1604 2095
rect 1678 2061 1712 2095
rect 1786 2061 1820 2095
rect 1894 2061 1928 2095
rect 2002 2061 2036 2095
rect 2110 2061 2144 2095
rect 2214 2061 2248 2095
<< psubdiff >>
rect 2310 109 2360 133
rect 2310 75 2318 109
rect 2352 75 2360 109
rect 2310 51 2360 75
<< nsubdiff >>
rect 2310 2541 2360 2565
rect 2310 2507 2318 2541
rect 2352 2507 2360 2541
rect 2310 2483 2360 2507
<< psubdiffcont >>
rect 2318 75 2352 109
<< nsubdiffcont >>
rect 2318 2507 2352 2541
<< poly >>
rect 114 2578 144 2604
rect 222 2578 252 2604
rect 330 2578 360 2604
rect 438 2578 468 2604
rect 546 2578 576 2604
rect 654 2578 684 2604
rect 762 2578 792 2604
rect 870 2578 900 2604
rect 978 2578 1008 2604
rect 1086 2578 1116 2604
rect 1194 2578 1224 2604
rect 1302 2578 1332 2604
rect 1410 2578 1440 2604
rect 1518 2578 1548 2604
rect 1626 2578 1656 2604
rect 1734 2578 1764 2604
rect 1842 2578 1872 2604
rect 1950 2578 1980 2604
rect 2058 2578 2088 2604
rect 2166 2578 2196 2604
rect 114 1552 144 1578
rect 222 1552 252 1578
rect 330 1552 360 1578
rect 438 1552 468 1578
rect 546 1552 576 1578
rect 654 1552 684 1578
rect 762 1552 792 1578
rect 870 1552 900 1578
rect 978 1552 1008 1578
rect 1086 1552 1116 1578
rect 1194 1552 1224 1578
rect 1302 1552 1332 1578
rect 1410 1552 1440 1578
rect 1518 1552 1548 1578
rect 1626 1552 1656 1578
rect 1734 1552 1764 1578
rect 1842 1552 1872 1578
rect 1950 1552 1980 1578
rect 2058 1552 2088 1578
rect 2166 1552 2196 1578
rect 114 1522 2196 1552
rect 114 1348 144 1522
rect 48 1332 144 1348
rect 48 1298 64 1332
rect 98 1298 144 1332
rect 48 1282 144 1298
rect 114 1107 144 1282
rect 114 1077 2196 1107
rect 114 1051 144 1077
rect 222 1051 252 1077
rect 330 1051 360 1077
rect 438 1051 468 1077
rect 546 1051 576 1077
rect 654 1051 684 1077
rect 762 1051 792 1077
rect 870 1051 900 1077
rect 978 1051 1008 1077
rect 1086 1051 1116 1077
rect 1194 1051 1224 1077
rect 1302 1051 1332 1077
rect 1410 1051 1440 1077
rect 1518 1051 1548 1077
rect 1626 1051 1656 1077
rect 1734 1051 1764 1077
rect 1842 1051 1872 1077
rect 1950 1051 1980 1077
rect 2058 1051 2088 1077
rect 2166 1051 2196 1077
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
rect 438 25 468 51
rect 546 25 576 51
rect 654 25 684 51
rect 762 25 792 51
rect 870 25 900 51
rect 978 25 1008 51
rect 1086 25 1116 51
rect 1194 25 1224 51
rect 1302 25 1332 51
rect 1410 25 1440 51
rect 1518 25 1548 51
rect 1626 25 1656 51
rect 1734 25 1764 51
rect 1842 25 1872 51
rect 1950 25 1980 51
rect 2058 25 2088 51
rect 2166 25 2196 51
<< polycont >>
rect 64 1298 98 1332
<< locali >>
rect 0 2612 2420 2646
rect 62 2095 96 2612
rect 62 2045 96 2061
rect 166 2095 200 2111
rect 166 2011 200 2061
rect 274 2095 308 2612
rect 274 2045 308 2061
rect 382 2095 416 2111
rect 382 2011 416 2061
rect 490 2095 524 2612
rect 490 2045 524 2061
rect 598 2095 632 2111
rect 598 2011 632 2061
rect 706 2095 740 2612
rect 706 2045 740 2061
rect 814 2095 848 2111
rect 814 2011 848 2061
rect 922 2095 956 2612
rect 922 2045 956 2061
rect 1030 2095 1064 2111
rect 1030 2011 1064 2061
rect 1138 2095 1172 2612
rect 1138 2045 1172 2061
rect 1246 2095 1280 2111
rect 1246 2011 1280 2061
rect 1354 2095 1388 2612
rect 1354 2045 1388 2061
rect 1462 2095 1496 2111
rect 1462 2011 1496 2061
rect 1570 2095 1604 2612
rect 1570 2045 1604 2061
rect 1678 2095 1712 2111
rect 1678 2011 1712 2061
rect 1786 2095 1820 2612
rect 1786 2045 1820 2061
rect 1894 2095 1928 2111
rect 1894 2011 1928 2061
rect 2002 2095 2036 2612
rect 2002 2045 2036 2061
rect 2110 2095 2144 2111
rect 2110 2011 2144 2061
rect 2214 2095 2248 2612
rect 2318 2541 2352 2612
rect 2318 2491 2352 2507
rect 2214 2045 2248 2061
rect 166 1977 2144 2011
rect 64 1332 98 1348
rect 64 1282 98 1298
rect 1138 1332 1172 1977
rect 1138 1298 1189 1332
rect 1138 652 1172 1298
rect 166 618 2144 652
rect 62 568 96 584
rect 62 17 96 534
rect 166 568 200 618
rect 166 518 200 534
rect 274 568 308 584
rect 274 17 308 534
rect 382 568 416 618
rect 382 518 416 534
rect 490 568 524 584
rect 490 17 524 534
rect 598 568 632 618
rect 598 518 632 534
rect 706 568 740 584
rect 706 17 740 534
rect 814 568 848 618
rect 814 518 848 534
rect 922 568 956 584
rect 922 17 956 534
rect 1030 568 1064 618
rect 1030 518 1064 534
rect 1138 568 1172 584
rect 1138 17 1172 534
rect 1246 568 1280 618
rect 1246 518 1280 534
rect 1354 568 1388 584
rect 1354 17 1388 534
rect 1462 568 1496 618
rect 1462 518 1496 534
rect 1570 568 1604 584
rect 1570 17 1604 534
rect 1678 568 1712 618
rect 1678 518 1712 534
rect 1786 568 1820 584
rect 1786 17 1820 534
rect 1894 568 1928 618
rect 1894 518 1928 534
rect 2002 568 2036 584
rect 2002 17 2036 534
rect 2110 568 2144 618
rect 2110 518 2144 534
rect 2214 568 2248 584
rect 2214 17 2248 534
rect 2318 109 2352 125
rect 2318 17 2352 75
rect 0 -17 2420 17
<< labels >>
rlabel locali s 81 1315 81 1315 4 A
port 1 nsew
rlabel locali s 1172 1315 1172 1315 4 Z
port 2 nsew
rlabel locali s 1210 0 1210 0 4 gnd
port 3 nsew
rlabel locali s 1210 2629 1210 2629 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2420 1994
<< end >>
