magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1296 -1277 3848 3436
<< nwell >>
rect -36 1017 2588 2176
<< locali >>
rect 0 2101 2552 2135
rect 64 988 98 1054
rect 179 1016 449 1050
rect 551 1006 925 1040
rect 1135 992 1617 1026
rect 2041 992 2075 1026
rect 0 -17 2552 17
use sky130_rom_krom_pinv  sky130_rom_krom_pinv_0
timestamp 1581321264
transform 1 0 0 0 1 0
box -36 -17 404 2176
use sky130_rom_krom_pinv_0  sky130_rom_krom_pinv_0_0
timestamp 1581321264
transform 1 0 368 0 1 0
box -36 -17 512 2176
use sky130_rom_krom_pinv_1  sky130_rom_krom_pinv_1_0
timestamp 1581321264
transform 1 0 844 0 1 0
box -36 -17 728 2176
use sky130_rom_krom_pinv_2  sky130_rom_krom_pinv_2_0
timestamp 1581321264
transform 1 0 1536 0 1 0
box -36 -17 1052 2176
<< labels >>
rlabel locali s 2058 1009 2058 1009 4 Z
port 1 nsew
rlabel locali s 81 1021 81 1021 4 A
port 2 nsew
rlabel locali s 1276 0 1276 0 4 gnd
port 3 nsew
rlabel locali s 1276 2118 1276 2118 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2552 2118
<< end >>
