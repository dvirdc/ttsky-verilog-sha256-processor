magic
tech sky130A
magscale 1 2
timestamp 1581398725
<< checkpaint >>
rect -1296 -1277 2312 3946
<< nwell >>
rect -36 1262 1052 2686
<< pwell >>
rect 28 159 878 677
rect 28 25 982 159
<< scnmos >>
rect 114 51 144 651
rect 222 51 252 651
rect 330 51 360 651
rect 438 51 468 651
rect 546 51 576 651
rect 654 51 684 651
rect 762 51 792 651
<< scpmos >>
rect 114 1578 144 2578
rect 222 1578 252 2578
rect 330 1578 360 2578
rect 438 1578 468 2578
rect 546 1578 576 2578
rect 654 1578 684 2578
rect 762 1578 792 2578
<< ndiff >>
rect 54 368 114 651
rect 54 334 62 368
rect 96 334 114 368
rect 54 51 114 334
rect 144 368 222 651
rect 144 334 166 368
rect 200 334 222 368
rect 144 51 222 334
rect 252 368 330 651
rect 252 334 274 368
rect 308 334 330 368
rect 252 51 330 334
rect 360 368 438 651
rect 360 334 382 368
rect 416 334 438 368
rect 360 51 438 334
rect 468 368 546 651
rect 468 334 490 368
rect 524 334 546 368
rect 468 51 546 334
rect 576 368 654 651
rect 576 334 598 368
rect 632 334 654 368
rect 576 51 654 334
rect 684 368 762 651
rect 684 334 706 368
rect 740 334 762 368
rect 684 51 762 334
rect 792 368 852 651
rect 792 334 810 368
rect 844 334 852 368
rect 792 51 852 334
<< pdiff >>
rect 54 2095 114 2578
rect 54 2061 62 2095
rect 96 2061 114 2095
rect 54 1578 114 2061
rect 144 2095 222 2578
rect 144 2061 166 2095
rect 200 2061 222 2095
rect 144 1578 222 2061
rect 252 2095 330 2578
rect 252 2061 274 2095
rect 308 2061 330 2095
rect 252 1578 330 2061
rect 360 2095 438 2578
rect 360 2061 382 2095
rect 416 2061 438 2095
rect 360 1578 438 2061
rect 468 2095 546 2578
rect 468 2061 490 2095
rect 524 2061 546 2095
rect 468 1578 546 2061
rect 576 2095 654 2578
rect 576 2061 598 2095
rect 632 2061 654 2095
rect 576 1578 654 2061
rect 684 2095 762 2578
rect 684 2061 706 2095
rect 740 2061 762 2095
rect 684 1578 762 2061
rect 792 2095 852 2578
rect 792 2061 810 2095
rect 844 2061 852 2095
rect 792 1578 852 2061
<< ndiffc >>
rect 62 334 96 368
rect 166 334 200 368
rect 274 334 308 368
rect 382 334 416 368
rect 490 334 524 368
rect 598 334 632 368
rect 706 334 740 368
rect 810 334 844 368
<< pdiffc >>
rect 62 2061 96 2095
rect 166 2061 200 2095
rect 274 2061 308 2095
rect 382 2061 416 2095
rect 490 2061 524 2095
rect 598 2061 632 2095
rect 706 2061 740 2095
rect 810 2061 844 2095
<< psubdiff >>
rect 906 109 956 133
rect 906 75 914 109
rect 948 75 956 109
rect 906 51 956 75
<< nsubdiff >>
rect 906 2541 956 2565
rect 906 2507 914 2541
rect 948 2507 956 2541
rect 906 2483 956 2507
<< psubdiffcont >>
rect 914 75 948 109
<< nsubdiffcont >>
rect 914 2507 948 2541
<< poly >>
rect 114 2578 144 2604
rect 222 2578 252 2604
rect 330 2578 360 2604
rect 438 2578 468 2604
rect 546 2578 576 2604
rect 654 2578 684 2604
rect 762 2578 792 2604
rect 114 1552 144 1578
rect 222 1552 252 1578
rect 330 1552 360 1578
rect 438 1552 468 1578
rect 546 1552 576 1578
rect 654 1552 684 1578
rect 762 1552 792 1578
rect 114 1522 792 1552
rect 114 1248 144 1522
rect 48 1232 144 1248
rect 48 1198 64 1232
rect 98 1198 144 1232
rect 48 1182 144 1198
rect 114 707 144 1182
rect 114 677 792 707
rect 114 651 144 677
rect 222 651 252 677
rect 330 651 360 677
rect 438 651 468 677
rect 546 651 576 677
rect 654 651 684 677
rect 762 651 792 677
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
rect 438 25 468 51
rect 546 25 576 51
rect 654 25 684 51
rect 762 25 792 51
<< polycont >>
rect 64 1198 98 1232
<< locali >>
rect 0 2612 1016 2646
rect 62 2095 96 2612
rect 62 2045 96 2061
rect 166 2095 200 2111
rect 166 2011 200 2061
rect 274 2095 308 2612
rect 274 2045 308 2061
rect 382 2095 416 2111
rect 382 2011 416 2061
rect 490 2095 524 2612
rect 490 2045 524 2061
rect 598 2095 632 2111
rect 598 2011 632 2061
rect 706 2095 740 2612
rect 914 2541 948 2612
rect 914 2491 948 2507
rect 706 2045 740 2061
rect 810 2095 844 2111
rect 810 2011 844 2061
rect 166 1977 844 2011
rect 64 1232 98 1248
rect 64 1182 98 1198
rect 488 1232 522 1977
rect 488 1198 539 1232
rect 488 452 522 1198
rect 166 418 844 452
rect 62 368 96 384
rect 62 17 96 334
rect 166 368 200 418
rect 166 318 200 334
rect 274 368 308 384
rect 274 17 308 334
rect 382 368 416 418
rect 382 318 416 334
rect 490 368 524 384
rect 490 17 524 334
rect 598 368 632 418
rect 598 318 632 334
rect 706 368 740 384
rect 706 17 740 334
rect 810 368 844 418
rect 810 318 844 334
rect 914 109 948 125
rect 914 17 948 75
rect 0 -17 1016 17
<< labels >>
rlabel locali s 81 1215 81 1215 4 A
port 1 nsew
rlabel locali s 522 1215 522 1215 4 Z
port 2 nsew
rlabel locali s 508 0 508 0 4 gnd
port 3 nsew
rlabel locali s 508 2629 508 2629 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1016 1994
<< end >>
