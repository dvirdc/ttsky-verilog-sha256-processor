magic
tech sky130A
magscale 1 2
timestamp 1581449089
<< checkpaint >>
rect -1260 -878 53535 4321
<< poly >>
rect 87 641 117 2272
rect 291 845 321 2272
rect 495 1049 525 2272
rect 699 1253 729 2272
rect 903 1457 933 2272
rect 1107 1661 1137 2272
rect 1311 1865 1341 2272
rect 1515 2069 1545 2272
rect 1606 2071 1672 2087
rect 1606 2069 1622 2071
rect 1515 2039 1622 2069
rect 1606 2037 1622 2039
rect 1656 2037 1672 2071
rect 1606 2021 1672 2037
rect 1402 1867 1468 1883
rect 1402 1865 1418 1867
rect 1311 1835 1418 1865
rect 1402 1833 1418 1835
rect 1452 1833 1468 1867
rect 1402 1817 1468 1833
rect 1198 1663 1264 1679
rect 1198 1661 1214 1663
rect 1107 1631 1214 1661
rect 1198 1629 1214 1631
rect 1248 1629 1264 1663
rect 1198 1613 1264 1629
rect 994 1459 1060 1475
rect 994 1457 1010 1459
rect 903 1427 1010 1457
rect 994 1425 1010 1427
rect 1044 1425 1060 1459
rect 994 1409 1060 1425
rect 790 1255 856 1271
rect 790 1253 806 1255
rect 699 1223 806 1253
rect 790 1221 806 1223
rect 840 1221 856 1255
rect 790 1205 856 1221
rect 586 1051 652 1067
rect 586 1049 602 1051
rect 495 1019 602 1049
rect 586 1017 602 1019
rect 636 1017 652 1051
rect 586 1001 652 1017
rect 382 847 448 863
rect 382 845 398 847
rect 291 815 398 845
rect 382 813 398 815
rect 432 813 448 847
rect 382 797 448 813
rect 178 643 244 659
rect 178 641 194 643
rect 87 611 194 641
rect 178 609 194 611
rect 228 609 244 643
rect 1719 641 1749 2272
rect 1923 845 1953 2272
rect 2127 1049 2157 2272
rect 2331 1253 2361 2272
rect 2535 1457 2565 2272
rect 2739 1661 2769 2272
rect 2943 1865 2973 2272
rect 3147 2069 3177 2272
rect 3238 2071 3304 2087
rect 3238 2069 3254 2071
rect 3147 2039 3254 2069
rect 3238 2037 3254 2039
rect 3288 2037 3304 2071
rect 3238 2021 3304 2037
rect 3034 1867 3100 1883
rect 3034 1865 3050 1867
rect 2943 1835 3050 1865
rect 3034 1833 3050 1835
rect 3084 1833 3100 1867
rect 3034 1817 3100 1833
rect 2830 1663 2896 1679
rect 2830 1661 2846 1663
rect 2739 1631 2846 1661
rect 2830 1629 2846 1631
rect 2880 1629 2896 1663
rect 2830 1613 2896 1629
rect 2626 1459 2692 1475
rect 2626 1457 2642 1459
rect 2535 1427 2642 1457
rect 2626 1425 2642 1427
rect 2676 1425 2692 1459
rect 2626 1409 2692 1425
rect 2422 1255 2488 1271
rect 2422 1253 2438 1255
rect 2331 1223 2438 1253
rect 2422 1221 2438 1223
rect 2472 1221 2488 1255
rect 2422 1205 2488 1221
rect 2218 1051 2284 1067
rect 2218 1049 2234 1051
rect 2127 1019 2234 1049
rect 2218 1017 2234 1019
rect 2268 1017 2284 1051
rect 2218 1001 2284 1017
rect 2014 847 2080 863
rect 2014 845 2030 847
rect 1923 815 2030 845
rect 2014 813 2030 815
rect 2064 813 2080 847
rect 2014 797 2080 813
rect 1810 643 1876 659
rect 1810 641 1826 643
rect 1719 611 1826 641
rect 178 593 244 609
rect 1810 609 1826 611
rect 1860 609 1876 643
rect 3351 641 3381 2272
rect 3555 845 3585 2272
rect 3759 1049 3789 2272
rect 3963 1253 3993 2272
rect 4167 1457 4197 2272
rect 4371 1661 4401 2272
rect 4575 1865 4605 2272
rect 4779 2069 4809 2272
rect 4870 2071 4936 2087
rect 4870 2069 4886 2071
rect 4779 2039 4886 2069
rect 4870 2037 4886 2039
rect 4920 2037 4936 2071
rect 4870 2021 4936 2037
rect 4666 1867 4732 1883
rect 4666 1865 4682 1867
rect 4575 1835 4682 1865
rect 4666 1833 4682 1835
rect 4716 1833 4732 1867
rect 4666 1817 4732 1833
rect 4462 1663 4528 1679
rect 4462 1661 4478 1663
rect 4371 1631 4478 1661
rect 4462 1629 4478 1631
rect 4512 1629 4528 1663
rect 4462 1613 4528 1629
rect 4258 1459 4324 1475
rect 4258 1457 4274 1459
rect 4167 1427 4274 1457
rect 4258 1425 4274 1427
rect 4308 1425 4324 1459
rect 4258 1409 4324 1425
rect 4054 1255 4120 1271
rect 4054 1253 4070 1255
rect 3963 1223 4070 1253
rect 4054 1221 4070 1223
rect 4104 1221 4120 1255
rect 4054 1205 4120 1221
rect 3850 1051 3916 1067
rect 3850 1049 3866 1051
rect 3759 1019 3866 1049
rect 3850 1017 3866 1019
rect 3900 1017 3916 1051
rect 3850 1001 3916 1017
rect 3646 847 3712 863
rect 3646 845 3662 847
rect 3555 815 3662 845
rect 3646 813 3662 815
rect 3696 813 3712 847
rect 3646 797 3712 813
rect 3442 643 3508 659
rect 3442 641 3458 643
rect 3351 611 3458 641
rect 1810 593 1876 609
rect 3442 609 3458 611
rect 3492 609 3508 643
rect 4983 641 5013 2272
rect 5187 845 5217 2272
rect 5391 1049 5421 2272
rect 5595 1253 5625 2272
rect 5799 1457 5829 2272
rect 6003 1661 6033 2272
rect 6207 1865 6237 2272
rect 6411 2069 6441 2272
rect 6502 2071 6568 2087
rect 6502 2069 6518 2071
rect 6411 2039 6518 2069
rect 6502 2037 6518 2039
rect 6552 2037 6568 2071
rect 6502 2021 6568 2037
rect 6298 1867 6364 1883
rect 6298 1865 6314 1867
rect 6207 1835 6314 1865
rect 6298 1833 6314 1835
rect 6348 1833 6364 1867
rect 6298 1817 6364 1833
rect 6094 1663 6160 1679
rect 6094 1661 6110 1663
rect 6003 1631 6110 1661
rect 6094 1629 6110 1631
rect 6144 1629 6160 1663
rect 6094 1613 6160 1629
rect 5890 1459 5956 1475
rect 5890 1457 5906 1459
rect 5799 1427 5906 1457
rect 5890 1425 5906 1427
rect 5940 1425 5956 1459
rect 5890 1409 5956 1425
rect 5686 1255 5752 1271
rect 5686 1253 5702 1255
rect 5595 1223 5702 1253
rect 5686 1221 5702 1223
rect 5736 1221 5752 1255
rect 5686 1205 5752 1221
rect 5482 1051 5548 1067
rect 5482 1049 5498 1051
rect 5391 1019 5498 1049
rect 5482 1017 5498 1019
rect 5532 1017 5548 1051
rect 5482 1001 5548 1017
rect 5278 847 5344 863
rect 5278 845 5294 847
rect 5187 815 5294 845
rect 5278 813 5294 815
rect 5328 813 5344 847
rect 5278 797 5344 813
rect 5074 643 5140 659
rect 5074 641 5090 643
rect 4983 611 5090 641
rect 3442 593 3508 609
rect 5074 609 5090 611
rect 5124 609 5140 643
rect 6615 641 6645 2272
rect 6819 845 6849 2272
rect 7023 1049 7053 2272
rect 7227 1253 7257 2272
rect 7431 1457 7461 2272
rect 7635 1661 7665 2272
rect 7839 1865 7869 2272
rect 8043 2069 8073 2272
rect 8134 2071 8200 2087
rect 8134 2069 8150 2071
rect 8043 2039 8150 2069
rect 8134 2037 8150 2039
rect 8184 2037 8200 2071
rect 8134 2021 8200 2037
rect 7930 1867 7996 1883
rect 7930 1865 7946 1867
rect 7839 1835 7946 1865
rect 7930 1833 7946 1835
rect 7980 1833 7996 1867
rect 7930 1817 7996 1833
rect 7726 1663 7792 1679
rect 7726 1661 7742 1663
rect 7635 1631 7742 1661
rect 7726 1629 7742 1631
rect 7776 1629 7792 1663
rect 7726 1613 7792 1629
rect 7522 1459 7588 1475
rect 7522 1457 7538 1459
rect 7431 1427 7538 1457
rect 7522 1425 7538 1427
rect 7572 1425 7588 1459
rect 7522 1409 7588 1425
rect 7318 1255 7384 1271
rect 7318 1253 7334 1255
rect 7227 1223 7334 1253
rect 7318 1221 7334 1223
rect 7368 1221 7384 1255
rect 7318 1205 7384 1221
rect 7114 1051 7180 1067
rect 7114 1049 7130 1051
rect 7023 1019 7130 1049
rect 7114 1017 7130 1019
rect 7164 1017 7180 1051
rect 7114 1001 7180 1017
rect 6910 847 6976 863
rect 6910 845 6926 847
rect 6819 815 6926 845
rect 6910 813 6926 815
rect 6960 813 6976 847
rect 6910 797 6976 813
rect 6706 643 6772 659
rect 6706 641 6722 643
rect 6615 611 6722 641
rect 5074 593 5140 609
rect 6706 609 6722 611
rect 6756 609 6772 643
rect 8247 641 8277 2272
rect 8451 845 8481 2272
rect 8655 1049 8685 2272
rect 8859 1253 8889 2272
rect 9063 1457 9093 2272
rect 9267 1661 9297 2272
rect 9471 1865 9501 2272
rect 9675 2069 9705 2272
rect 9766 2071 9832 2087
rect 9766 2069 9782 2071
rect 9675 2039 9782 2069
rect 9766 2037 9782 2039
rect 9816 2037 9832 2071
rect 9766 2021 9832 2037
rect 9562 1867 9628 1883
rect 9562 1865 9578 1867
rect 9471 1835 9578 1865
rect 9562 1833 9578 1835
rect 9612 1833 9628 1867
rect 9562 1817 9628 1833
rect 9358 1663 9424 1679
rect 9358 1661 9374 1663
rect 9267 1631 9374 1661
rect 9358 1629 9374 1631
rect 9408 1629 9424 1663
rect 9358 1613 9424 1629
rect 9154 1459 9220 1475
rect 9154 1457 9170 1459
rect 9063 1427 9170 1457
rect 9154 1425 9170 1427
rect 9204 1425 9220 1459
rect 9154 1409 9220 1425
rect 8950 1255 9016 1271
rect 8950 1253 8966 1255
rect 8859 1223 8966 1253
rect 8950 1221 8966 1223
rect 9000 1221 9016 1255
rect 8950 1205 9016 1221
rect 8746 1051 8812 1067
rect 8746 1049 8762 1051
rect 8655 1019 8762 1049
rect 8746 1017 8762 1019
rect 8796 1017 8812 1051
rect 8746 1001 8812 1017
rect 8542 847 8608 863
rect 8542 845 8558 847
rect 8451 815 8558 845
rect 8542 813 8558 815
rect 8592 813 8608 847
rect 8542 797 8608 813
rect 8338 643 8404 659
rect 8338 641 8354 643
rect 8247 611 8354 641
rect 6706 593 6772 609
rect 8338 609 8354 611
rect 8388 609 8404 643
rect 9879 641 9909 2272
rect 10083 845 10113 2272
rect 10287 1049 10317 2272
rect 10491 1253 10521 2272
rect 10695 1457 10725 2272
rect 10899 1661 10929 2272
rect 11103 1865 11133 2272
rect 11307 2069 11337 2272
rect 11398 2071 11464 2087
rect 11398 2069 11414 2071
rect 11307 2039 11414 2069
rect 11398 2037 11414 2039
rect 11448 2037 11464 2071
rect 11398 2021 11464 2037
rect 11194 1867 11260 1883
rect 11194 1865 11210 1867
rect 11103 1835 11210 1865
rect 11194 1833 11210 1835
rect 11244 1833 11260 1867
rect 11194 1817 11260 1833
rect 10990 1663 11056 1679
rect 10990 1661 11006 1663
rect 10899 1631 11006 1661
rect 10990 1629 11006 1631
rect 11040 1629 11056 1663
rect 10990 1613 11056 1629
rect 10786 1459 10852 1475
rect 10786 1457 10802 1459
rect 10695 1427 10802 1457
rect 10786 1425 10802 1427
rect 10836 1425 10852 1459
rect 10786 1409 10852 1425
rect 10582 1255 10648 1271
rect 10582 1253 10598 1255
rect 10491 1223 10598 1253
rect 10582 1221 10598 1223
rect 10632 1221 10648 1255
rect 10582 1205 10648 1221
rect 10378 1051 10444 1067
rect 10378 1049 10394 1051
rect 10287 1019 10394 1049
rect 10378 1017 10394 1019
rect 10428 1017 10444 1051
rect 10378 1001 10444 1017
rect 10174 847 10240 863
rect 10174 845 10190 847
rect 10083 815 10190 845
rect 10174 813 10190 815
rect 10224 813 10240 847
rect 10174 797 10240 813
rect 9970 643 10036 659
rect 9970 641 9986 643
rect 9879 611 9986 641
rect 8338 593 8404 609
rect 9970 609 9986 611
rect 10020 609 10036 643
rect 11511 641 11541 2272
rect 11715 845 11745 2272
rect 11919 1049 11949 2272
rect 12123 1253 12153 2272
rect 12327 1457 12357 2272
rect 12531 1661 12561 2272
rect 12735 1865 12765 2272
rect 12939 2069 12969 2272
rect 13030 2071 13096 2087
rect 13030 2069 13046 2071
rect 12939 2039 13046 2069
rect 13030 2037 13046 2039
rect 13080 2037 13096 2071
rect 13030 2021 13096 2037
rect 12826 1867 12892 1883
rect 12826 1865 12842 1867
rect 12735 1835 12842 1865
rect 12826 1833 12842 1835
rect 12876 1833 12892 1867
rect 12826 1817 12892 1833
rect 12622 1663 12688 1679
rect 12622 1661 12638 1663
rect 12531 1631 12638 1661
rect 12622 1629 12638 1631
rect 12672 1629 12688 1663
rect 12622 1613 12688 1629
rect 12418 1459 12484 1475
rect 12418 1457 12434 1459
rect 12327 1427 12434 1457
rect 12418 1425 12434 1427
rect 12468 1425 12484 1459
rect 12418 1409 12484 1425
rect 12214 1255 12280 1271
rect 12214 1253 12230 1255
rect 12123 1223 12230 1253
rect 12214 1221 12230 1223
rect 12264 1221 12280 1255
rect 12214 1205 12280 1221
rect 12010 1051 12076 1067
rect 12010 1049 12026 1051
rect 11919 1019 12026 1049
rect 12010 1017 12026 1019
rect 12060 1017 12076 1051
rect 12010 1001 12076 1017
rect 11806 847 11872 863
rect 11806 845 11822 847
rect 11715 815 11822 845
rect 11806 813 11822 815
rect 11856 813 11872 847
rect 11806 797 11872 813
rect 11602 643 11668 659
rect 11602 641 11618 643
rect 11511 611 11618 641
rect 9970 593 10036 609
rect 11602 609 11618 611
rect 11652 609 11668 643
rect 13143 641 13173 2272
rect 13347 845 13377 2272
rect 13551 1049 13581 2272
rect 13755 1253 13785 2272
rect 13959 1457 13989 2272
rect 14163 1661 14193 2272
rect 14367 1865 14397 2272
rect 14571 2069 14601 2272
rect 14662 2071 14728 2087
rect 14662 2069 14678 2071
rect 14571 2039 14678 2069
rect 14662 2037 14678 2039
rect 14712 2037 14728 2071
rect 14662 2021 14728 2037
rect 14458 1867 14524 1883
rect 14458 1865 14474 1867
rect 14367 1835 14474 1865
rect 14458 1833 14474 1835
rect 14508 1833 14524 1867
rect 14458 1817 14524 1833
rect 14254 1663 14320 1679
rect 14254 1661 14270 1663
rect 14163 1631 14270 1661
rect 14254 1629 14270 1631
rect 14304 1629 14320 1663
rect 14254 1613 14320 1629
rect 14050 1459 14116 1475
rect 14050 1457 14066 1459
rect 13959 1427 14066 1457
rect 14050 1425 14066 1427
rect 14100 1425 14116 1459
rect 14050 1409 14116 1425
rect 13846 1255 13912 1271
rect 13846 1253 13862 1255
rect 13755 1223 13862 1253
rect 13846 1221 13862 1223
rect 13896 1221 13912 1255
rect 13846 1205 13912 1221
rect 13642 1051 13708 1067
rect 13642 1049 13658 1051
rect 13551 1019 13658 1049
rect 13642 1017 13658 1019
rect 13692 1017 13708 1051
rect 13642 1001 13708 1017
rect 13438 847 13504 863
rect 13438 845 13454 847
rect 13347 815 13454 845
rect 13438 813 13454 815
rect 13488 813 13504 847
rect 13438 797 13504 813
rect 13234 643 13300 659
rect 13234 641 13250 643
rect 13143 611 13250 641
rect 11602 593 11668 609
rect 13234 609 13250 611
rect 13284 609 13300 643
rect 14775 641 14805 2272
rect 14979 845 15009 2272
rect 15183 1049 15213 2272
rect 15387 1253 15417 2272
rect 15591 1457 15621 2272
rect 15795 1661 15825 2272
rect 15999 1865 16029 2272
rect 16203 2069 16233 2272
rect 16294 2071 16360 2087
rect 16294 2069 16310 2071
rect 16203 2039 16310 2069
rect 16294 2037 16310 2039
rect 16344 2037 16360 2071
rect 16294 2021 16360 2037
rect 16090 1867 16156 1883
rect 16090 1865 16106 1867
rect 15999 1835 16106 1865
rect 16090 1833 16106 1835
rect 16140 1833 16156 1867
rect 16090 1817 16156 1833
rect 15886 1663 15952 1679
rect 15886 1661 15902 1663
rect 15795 1631 15902 1661
rect 15886 1629 15902 1631
rect 15936 1629 15952 1663
rect 15886 1613 15952 1629
rect 15682 1459 15748 1475
rect 15682 1457 15698 1459
rect 15591 1427 15698 1457
rect 15682 1425 15698 1427
rect 15732 1425 15748 1459
rect 15682 1409 15748 1425
rect 15478 1255 15544 1271
rect 15478 1253 15494 1255
rect 15387 1223 15494 1253
rect 15478 1221 15494 1223
rect 15528 1221 15544 1255
rect 15478 1205 15544 1221
rect 15274 1051 15340 1067
rect 15274 1049 15290 1051
rect 15183 1019 15290 1049
rect 15274 1017 15290 1019
rect 15324 1017 15340 1051
rect 15274 1001 15340 1017
rect 15070 847 15136 863
rect 15070 845 15086 847
rect 14979 815 15086 845
rect 15070 813 15086 815
rect 15120 813 15136 847
rect 15070 797 15136 813
rect 14866 643 14932 659
rect 14866 641 14882 643
rect 14775 611 14882 641
rect 13234 593 13300 609
rect 14866 609 14882 611
rect 14916 609 14932 643
rect 16407 641 16437 2272
rect 16611 845 16641 2272
rect 16815 1049 16845 2272
rect 17019 1253 17049 2272
rect 17223 1457 17253 2272
rect 17427 1661 17457 2272
rect 17631 1865 17661 2272
rect 17835 2069 17865 2272
rect 17926 2071 17992 2087
rect 17926 2069 17942 2071
rect 17835 2039 17942 2069
rect 17926 2037 17942 2039
rect 17976 2037 17992 2071
rect 17926 2021 17992 2037
rect 17722 1867 17788 1883
rect 17722 1865 17738 1867
rect 17631 1835 17738 1865
rect 17722 1833 17738 1835
rect 17772 1833 17788 1867
rect 17722 1817 17788 1833
rect 17518 1663 17584 1679
rect 17518 1661 17534 1663
rect 17427 1631 17534 1661
rect 17518 1629 17534 1631
rect 17568 1629 17584 1663
rect 17518 1613 17584 1629
rect 17314 1459 17380 1475
rect 17314 1457 17330 1459
rect 17223 1427 17330 1457
rect 17314 1425 17330 1427
rect 17364 1425 17380 1459
rect 17314 1409 17380 1425
rect 17110 1255 17176 1271
rect 17110 1253 17126 1255
rect 17019 1223 17126 1253
rect 17110 1221 17126 1223
rect 17160 1221 17176 1255
rect 17110 1205 17176 1221
rect 16906 1051 16972 1067
rect 16906 1049 16922 1051
rect 16815 1019 16922 1049
rect 16906 1017 16922 1019
rect 16956 1017 16972 1051
rect 16906 1001 16972 1017
rect 16702 847 16768 863
rect 16702 845 16718 847
rect 16611 815 16718 845
rect 16702 813 16718 815
rect 16752 813 16768 847
rect 16702 797 16768 813
rect 16498 643 16564 659
rect 16498 641 16514 643
rect 16407 611 16514 641
rect 14866 593 14932 609
rect 16498 609 16514 611
rect 16548 609 16564 643
rect 18039 641 18069 2272
rect 18243 845 18273 2272
rect 18447 1049 18477 2272
rect 18651 1253 18681 2272
rect 18855 1457 18885 2272
rect 19059 1661 19089 2272
rect 19263 1865 19293 2272
rect 19467 2069 19497 2272
rect 19558 2071 19624 2087
rect 19558 2069 19574 2071
rect 19467 2039 19574 2069
rect 19558 2037 19574 2039
rect 19608 2037 19624 2071
rect 19558 2021 19624 2037
rect 19354 1867 19420 1883
rect 19354 1865 19370 1867
rect 19263 1835 19370 1865
rect 19354 1833 19370 1835
rect 19404 1833 19420 1867
rect 19354 1817 19420 1833
rect 19150 1663 19216 1679
rect 19150 1661 19166 1663
rect 19059 1631 19166 1661
rect 19150 1629 19166 1631
rect 19200 1629 19216 1663
rect 19150 1613 19216 1629
rect 18946 1459 19012 1475
rect 18946 1457 18962 1459
rect 18855 1427 18962 1457
rect 18946 1425 18962 1427
rect 18996 1425 19012 1459
rect 18946 1409 19012 1425
rect 18742 1255 18808 1271
rect 18742 1253 18758 1255
rect 18651 1223 18758 1253
rect 18742 1221 18758 1223
rect 18792 1221 18808 1255
rect 18742 1205 18808 1221
rect 18538 1051 18604 1067
rect 18538 1049 18554 1051
rect 18447 1019 18554 1049
rect 18538 1017 18554 1019
rect 18588 1017 18604 1051
rect 18538 1001 18604 1017
rect 18334 847 18400 863
rect 18334 845 18350 847
rect 18243 815 18350 845
rect 18334 813 18350 815
rect 18384 813 18400 847
rect 18334 797 18400 813
rect 18130 643 18196 659
rect 18130 641 18146 643
rect 18039 611 18146 641
rect 16498 593 16564 609
rect 18130 609 18146 611
rect 18180 609 18196 643
rect 19671 641 19701 2272
rect 19875 845 19905 2272
rect 20079 1049 20109 2272
rect 20283 1253 20313 2272
rect 20487 1457 20517 2272
rect 20691 1661 20721 2272
rect 20895 1865 20925 2272
rect 21099 2069 21129 2272
rect 21190 2071 21256 2087
rect 21190 2069 21206 2071
rect 21099 2039 21206 2069
rect 21190 2037 21206 2039
rect 21240 2037 21256 2071
rect 21190 2021 21256 2037
rect 20986 1867 21052 1883
rect 20986 1865 21002 1867
rect 20895 1835 21002 1865
rect 20986 1833 21002 1835
rect 21036 1833 21052 1867
rect 20986 1817 21052 1833
rect 20782 1663 20848 1679
rect 20782 1661 20798 1663
rect 20691 1631 20798 1661
rect 20782 1629 20798 1631
rect 20832 1629 20848 1663
rect 20782 1613 20848 1629
rect 20578 1459 20644 1475
rect 20578 1457 20594 1459
rect 20487 1427 20594 1457
rect 20578 1425 20594 1427
rect 20628 1425 20644 1459
rect 20578 1409 20644 1425
rect 20374 1255 20440 1271
rect 20374 1253 20390 1255
rect 20283 1223 20390 1253
rect 20374 1221 20390 1223
rect 20424 1221 20440 1255
rect 20374 1205 20440 1221
rect 20170 1051 20236 1067
rect 20170 1049 20186 1051
rect 20079 1019 20186 1049
rect 20170 1017 20186 1019
rect 20220 1017 20236 1051
rect 20170 1001 20236 1017
rect 19966 847 20032 863
rect 19966 845 19982 847
rect 19875 815 19982 845
rect 19966 813 19982 815
rect 20016 813 20032 847
rect 19966 797 20032 813
rect 19762 643 19828 659
rect 19762 641 19778 643
rect 19671 611 19778 641
rect 18130 593 18196 609
rect 19762 609 19778 611
rect 19812 609 19828 643
rect 21303 641 21333 2272
rect 21507 845 21537 2272
rect 21711 1049 21741 2272
rect 21915 1253 21945 2272
rect 22119 1457 22149 2272
rect 22323 1661 22353 2272
rect 22527 1865 22557 2272
rect 22731 2069 22761 2272
rect 22822 2071 22888 2087
rect 22822 2069 22838 2071
rect 22731 2039 22838 2069
rect 22822 2037 22838 2039
rect 22872 2037 22888 2071
rect 22822 2021 22888 2037
rect 22618 1867 22684 1883
rect 22618 1865 22634 1867
rect 22527 1835 22634 1865
rect 22618 1833 22634 1835
rect 22668 1833 22684 1867
rect 22618 1817 22684 1833
rect 22414 1663 22480 1679
rect 22414 1661 22430 1663
rect 22323 1631 22430 1661
rect 22414 1629 22430 1631
rect 22464 1629 22480 1663
rect 22414 1613 22480 1629
rect 22210 1459 22276 1475
rect 22210 1457 22226 1459
rect 22119 1427 22226 1457
rect 22210 1425 22226 1427
rect 22260 1425 22276 1459
rect 22210 1409 22276 1425
rect 22006 1255 22072 1271
rect 22006 1253 22022 1255
rect 21915 1223 22022 1253
rect 22006 1221 22022 1223
rect 22056 1221 22072 1255
rect 22006 1205 22072 1221
rect 21802 1051 21868 1067
rect 21802 1049 21818 1051
rect 21711 1019 21818 1049
rect 21802 1017 21818 1019
rect 21852 1017 21868 1051
rect 21802 1001 21868 1017
rect 21598 847 21664 863
rect 21598 845 21614 847
rect 21507 815 21614 845
rect 21598 813 21614 815
rect 21648 813 21664 847
rect 21598 797 21664 813
rect 21394 643 21460 659
rect 21394 641 21410 643
rect 21303 611 21410 641
rect 19762 593 19828 609
rect 21394 609 21410 611
rect 21444 609 21460 643
rect 22935 641 22965 2272
rect 23139 845 23169 2272
rect 23343 1049 23373 2272
rect 23547 1253 23577 2272
rect 23751 1457 23781 2272
rect 23955 1661 23985 2272
rect 24159 1865 24189 2272
rect 24363 2069 24393 2272
rect 24454 2071 24520 2087
rect 24454 2069 24470 2071
rect 24363 2039 24470 2069
rect 24454 2037 24470 2039
rect 24504 2037 24520 2071
rect 24454 2021 24520 2037
rect 24250 1867 24316 1883
rect 24250 1865 24266 1867
rect 24159 1835 24266 1865
rect 24250 1833 24266 1835
rect 24300 1833 24316 1867
rect 24250 1817 24316 1833
rect 24046 1663 24112 1679
rect 24046 1661 24062 1663
rect 23955 1631 24062 1661
rect 24046 1629 24062 1631
rect 24096 1629 24112 1663
rect 24046 1613 24112 1629
rect 23842 1459 23908 1475
rect 23842 1457 23858 1459
rect 23751 1427 23858 1457
rect 23842 1425 23858 1427
rect 23892 1425 23908 1459
rect 23842 1409 23908 1425
rect 23638 1255 23704 1271
rect 23638 1253 23654 1255
rect 23547 1223 23654 1253
rect 23638 1221 23654 1223
rect 23688 1221 23704 1255
rect 23638 1205 23704 1221
rect 23434 1051 23500 1067
rect 23434 1049 23450 1051
rect 23343 1019 23450 1049
rect 23434 1017 23450 1019
rect 23484 1017 23500 1051
rect 23434 1001 23500 1017
rect 23230 847 23296 863
rect 23230 845 23246 847
rect 23139 815 23246 845
rect 23230 813 23246 815
rect 23280 813 23296 847
rect 23230 797 23296 813
rect 23026 643 23092 659
rect 23026 641 23042 643
rect 22935 611 23042 641
rect 21394 593 21460 609
rect 23026 609 23042 611
rect 23076 609 23092 643
rect 24567 641 24597 2272
rect 24771 845 24801 2272
rect 24975 1049 25005 2272
rect 25179 1253 25209 2272
rect 25383 1457 25413 2272
rect 25587 1661 25617 2272
rect 25791 1865 25821 2272
rect 25995 2069 26025 2272
rect 26086 2071 26152 2087
rect 26086 2069 26102 2071
rect 25995 2039 26102 2069
rect 26086 2037 26102 2039
rect 26136 2037 26152 2071
rect 26086 2021 26152 2037
rect 25882 1867 25948 1883
rect 25882 1865 25898 1867
rect 25791 1835 25898 1865
rect 25882 1833 25898 1835
rect 25932 1833 25948 1867
rect 25882 1817 25948 1833
rect 25678 1663 25744 1679
rect 25678 1661 25694 1663
rect 25587 1631 25694 1661
rect 25678 1629 25694 1631
rect 25728 1629 25744 1663
rect 25678 1613 25744 1629
rect 25474 1459 25540 1475
rect 25474 1457 25490 1459
rect 25383 1427 25490 1457
rect 25474 1425 25490 1427
rect 25524 1425 25540 1459
rect 25474 1409 25540 1425
rect 25270 1255 25336 1271
rect 25270 1253 25286 1255
rect 25179 1223 25286 1253
rect 25270 1221 25286 1223
rect 25320 1221 25336 1255
rect 25270 1205 25336 1221
rect 25066 1051 25132 1067
rect 25066 1049 25082 1051
rect 24975 1019 25082 1049
rect 25066 1017 25082 1019
rect 25116 1017 25132 1051
rect 25066 1001 25132 1017
rect 24862 847 24928 863
rect 24862 845 24878 847
rect 24771 815 24878 845
rect 24862 813 24878 815
rect 24912 813 24928 847
rect 24862 797 24928 813
rect 24658 643 24724 659
rect 24658 641 24674 643
rect 24567 611 24674 641
rect 23026 593 23092 609
rect 24658 609 24674 611
rect 24708 609 24724 643
rect 26199 641 26229 2272
rect 26403 845 26433 2272
rect 26607 1049 26637 2272
rect 26811 1253 26841 2272
rect 27015 1457 27045 2272
rect 27219 1661 27249 2272
rect 27423 1865 27453 2272
rect 27627 2069 27657 2272
rect 27718 2071 27784 2087
rect 27718 2069 27734 2071
rect 27627 2039 27734 2069
rect 27718 2037 27734 2039
rect 27768 2037 27784 2071
rect 27718 2021 27784 2037
rect 27514 1867 27580 1883
rect 27514 1865 27530 1867
rect 27423 1835 27530 1865
rect 27514 1833 27530 1835
rect 27564 1833 27580 1867
rect 27514 1817 27580 1833
rect 27310 1663 27376 1679
rect 27310 1661 27326 1663
rect 27219 1631 27326 1661
rect 27310 1629 27326 1631
rect 27360 1629 27376 1663
rect 27310 1613 27376 1629
rect 27106 1459 27172 1475
rect 27106 1457 27122 1459
rect 27015 1427 27122 1457
rect 27106 1425 27122 1427
rect 27156 1425 27172 1459
rect 27106 1409 27172 1425
rect 26902 1255 26968 1271
rect 26902 1253 26918 1255
rect 26811 1223 26918 1253
rect 26902 1221 26918 1223
rect 26952 1221 26968 1255
rect 26902 1205 26968 1221
rect 26698 1051 26764 1067
rect 26698 1049 26714 1051
rect 26607 1019 26714 1049
rect 26698 1017 26714 1019
rect 26748 1017 26764 1051
rect 26698 1001 26764 1017
rect 26494 847 26560 863
rect 26494 845 26510 847
rect 26403 815 26510 845
rect 26494 813 26510 815
rect 26544 813 26560 847
rect 26494 797 26560 813
rect 26290 643 26356 659
rect 26290 641 26306 643
rect 26199 611 26306 641
rect 24658 593 24724 609
rect 26290 609 26306 611
rect 26340 609 26356 643
rect 27831 641 27861 2272
rect 28035 845 28065 2272
rect 28239 1049 28269 2272
rect 28443 1253 28473 2272
rect 28647 1457 28677 2272
rect 28851 1661 28881 2272
rect 29055 1865 29085 2272
rect 29259 2069 29289 2272
rect 29350 2071 29416 2087
rect 29350 2069 29366 2071
rect 29259 2039 29366 2069
rect 29350 2037 29366 2039
rect 29400 2037 29416 2071
rect 29350 2021 29416 2037
rect 29146 1867 29212 1883
rect 29146 1865 29162 1867
rect 29055 1835 29162 1865
rect 29146 1833 29162 1835
rect 29196 1833 29212 1867
rect 29146 1817 29212 1833
rect 28942 1663 29008 1679
rect 28942 1661 28958 1663
rect 28851 1631 28958 1661
rect 28942 1629 28958 1631
rect 28992 1629 29008 1663
rect 28942 1613 29008 1629
rect 28738 1459 28804 1475
rect 28738 1457 28754 1459
rect 28647 1427 28754 1457
rect 28738 1425 28754 1427
rect 28788 1425 28804 1459
rect 28738 1409 28804 1425
rect 28534 1255 28600 1271
rect 28534 1253 28550 1255
rect 28443 1223 28550 1253
rect 28534 1221 28550 1223
rect 28584 1221 28600 1255
rect 28534 1205 28600 1221
rect 28330 1051 28396 1067
rect 28330 1049 28346 1051
rect 28239 1019 28346 1049
rect 28330 1017 28346 1019
rect 28380 1017 28396 1051
rect 28330 1001 28396 1017
rect 28126 847 28192 863
rect 28126 845 28142 847
rect 28035 815 28142 845
rect 28126 813 28142 815
rect 28176 813 28192 847
rect 28126 797 28192 813
rect 27922 643 27988 659
rect 27922 641 27938 643
rect 27831 611 27938 641
rect 26290 593 26356 609
rect 27922 609 27938 611
rect 27972 609 27988 643
rect 29463 641 29493 2272
rect 29667 845 29697 2272
rect 29871 1049 29901 2272
rect 30075 1253 30105 2272
rect 30279 1457 30309 2272
rect 30483 1661 30513 2272
rect 30687 1865 30717 2272
rect 30891 2069 30921 2272
rect 30982 2071 31048 2087
rect 30982 2069 30998 2071
rect 30891 2039 30998 2069
rect 30982 2037 30998 2039
rect 31032 2037 31048 2071
rect 30982 2021 31048 2037
rect 30778 1867 30844 1883
rect 30778 1865 30794 1867
rect 30687 1835 30794 1865
rect 30778 1833 30794 1835
rect 30828 1833 30844 1867
rect 30778 1817 30844 1833
rect 30574 1663 30640 1679
rect 30574 1661 30590 1663
rect 30483 1631 30590 1661
rect 30574 1629 30590 1631
rect 30624 1629 30640 1663
rect 30574 1613 30640 1629
rect 30370 1459 30436 1475
rect 30370 1457 30386 1459
rect 30279 1427 30386 1457
rect 30370 1425 30386 1427
rect 30420 1425 30436 1459
rect 30370 1409 30436 1425
rect 30166 1255 30232 1271
rect 30166 1253 30182 1255
rect 30075 1223 30182 1253
rect 30166 1221 30182 1223
rect 30216 1221 30232 1255
rect 30166 1205 30232 1221
rect 29962 1051 30028 1067
rect 29962 1049 29978 1051
rect 29871 1019 29978 1049
rect 29962 1017 29978 1019
rect 30012 1017 30028 1051
rect 29962 1001 30028 1017
rect 29758 847 29824 863
rect 29758 845 29774 847
rect 29667 815 29774 845
rect 29758 813 29774 815
rect 29808 813 29824 847
rect 29758 797 29824 813
rect 29554 643 29620 659
rect 29554 641 29570 643
rect 29463 611 29570 641
rect 27922 593 27988 609
rect 29554 609 29570 611
rect 29604 609 29620 643
rect 31095 641 31125 2272
rect 31299 845 31329 2272
rect 31503 1049 31533 2272
rect 31707 1253 31737 2272
rect 31911 1457 31941 2272
rect 32115 1661 32145 2272
rect 32319 1865 32349 2272
rect 32523 2069 32553 2272
rect 32614 2071 32680 2087
rect 32614 2069 32630 2071
rect 32523 2039 32630 2069
rect 32614 2037 32630 2039
rect 32664 2037 32680 2071
rect 32614 2021 32680 2037
rect 32410 1867 32476 1883
rect 32410 1865 32426 1867
rect 32319 1835 32426 1865
rect 32410 1833 32426 1835
rect 32460 1833 32476 1867
rect 32410 1817 32476 1833
rect 32206 1663 32272 1679
rect 32206 1661 32222 1663
rect 32115 1631 32222 1661
rect 32206 1629 32222 1631
rect 32256 1629 32272 1663
rect 32206 1613 32272 1629
rect 32002 1459 32068 1475
rect 32002 1457 32018 1459
rect 31911 1427 32018 1457
rect 32002 1425 32018 1427
rect 32052 1425 32068 1459
rect 32002 1409 32068 1425
rect 31798 1255 31864 1271
rect 31798 1253 31814 1255
rect 31707 1223 31814 1253
rect 31798 1221 31814 1223
rect 31848 1221 31864 1255
rect 31798 1205 31864 1221
rect 31594 1051 31660 1067
rect 31594 1049 31610 1051
rect 31503 1019 31610 1049
rect 31594 1017 31610 1019
rect 31644 1017 31660 1051
rect 31594 1001 31660 1017
rect 31390 847 31456 863
rect 31390 845 31406 847
rect 31299 815 31406 845
rect 31390 813 31406 815
rect 31440 813 31456 847
rect 31390 797 31456 813
rect 31186 643 31252 659
rect 31186 641 31202 643
rect 31095 611 31202 641
rect 29554 593 29620 609
rect 31186 609 31202 611
rect 31236 609 31252 643
rect 32727 641 32757 2272
rect 32931 845 32961 2272
rect 33135 1049 33165 2272
rect 33339 1253 33369 2272
rect 33543 1457 33573 2272
rect 33747 1661 33777 2272
rect 33951 1865 33981 2272
rect 34155 2069 34185 2272
rect 34246 2071 34312 2087
rect 34246 2069 34262 2071
rect 34155 2039 34262 2069
rect 34246 2037 34262 2039
rect 34296 2037 34312 2071
rect 34246 2021 34312 2037
rect 34042 1867 34108 1883
rect 34042 1865 34058 1867
rect 33951 1835 34058 1865
rect 34042 1833 34058 1835
rect 34092 1833 34108 1867
rect 34042 1817 34108 1833
rect 33838 1663 33904 1679
rect 33838 1661 33854 1663
rect 33747 1631 33854 1661
rect 33838 1629 33854 1631
rect 33888 1629 33904 1663
rect 33838 1613 33904 1629
rect 33634 1459 33700 1475
rect 33634 1457 33650 1459
rect 33543 1427 33650 1457
rect 33634 1425 33650 1427
rect 33684 1425 33700 1459
rect 33634 1409 33700 1425
rect 33430 1255 33496 1271
rect 33430 1253 33446 1255
rect 33339 1223 33446 1253
rect 33430 1221 33446 1223
rect 33480 1221 33496 1255
rect 33430 1205 33496 1221
rect 33226 1051 33292 1067
rect 33226 1049 33242 1051
rect 33135 1019 33242 1049
rect 33226 1017 33242 1019
rect 33276 1017 33292 1051
rect 33226 1001 33292 1017
rect 33022 847 33088 863
rect 33022 845 33038 847
rect 32931 815 33038 845
rect 33022 813 33038 815
rect 33072 813 33088 847
rect 33022 797 33088 813
rect 32818 643 32884 659
rect 32818 641 32834 643
rect 32727 611 32834 641
rect 31186 593 31252 609
rect 32818 609 32834 611
rect 32868 609 32884 643
rect 34359 641 34389 2272
rect 34563 845 34593 2272
rect 34767 1049 34797 2272
rect 34971 1253 35001 2272
rect 35175 1457 35205 2272
rect 35379 1661 35409 2272
rect 35583 1865 35613 2272
rect 35787 2069 35817 2272
rect 35878 2071 35944 2087
rect 35878 2069 35894 2071
rect 35787 2039 35894 2069
rect 35878 2037 35894 2039
rect 35928 2037 35944 2071
rect 35878 2021 35944 2037
rect 35674 1867 35740 1883
rect 35674 1865 35690 1867
rect 35583 1835 35690 1865
rect 35674 1833 35690 1835
rect 35724 1833 35740 1867
rect 35674 1817 35740 1833
rect 35470 1663 35536 1679
rect 35470 1661 35486 1663
rect 35379 1631 35486 1661
rect 35470 1629 35486 1631
rect 35520 1629 35536 1663
rect 35470 1613 35536 1629
rect 35266 1459 35332 1475
rect 35266 1457 35282 1459
rect 35175 1427 35282 1457
rect 35266 1425 35282 1427
rect 35316 1425 35332 1459
rect 35266 1409 35332 1425
rect 35062 1255 35128 1271
rect 35062 1253 35078 1255
rect 34971 1223 35078 1253
rect 35062 1221 35078 1223
rect 35112 1221 35128 1255
rect 35062 1205 35128 1221
rect 34858 1051 34924 1067
rect 34858 1049 34874 1051
rect 34767 1019 34874 1049
rect 34858 1017 34874 1019
rect 34908 1017 34924 1051
rect 34858 1001 34924 1017
rect 34654 847 34720 863
rect 34654 845 34670 847
rect 34563 815 34670 845
rect 34654 813 34670 815
rect 34704 813 34720 847
rect 34654 797 34720 813
rect 34450 643 34516 659
rect 34450 641 34466 643
rect 34359 611 34466 641
rect 32818 593 32884 609
rect 34450 609 34466 611
rect 34500 609 34516 643
rect 35991 641 36021 2272
rect 36195 845 36225 2272
rect 36399 1049 36429 2272
rect 36603 1253 36633 2272
rect 36807 1457 36837 2272
rect 37011 1661 37041 2272
rect 37215 1865 37245 2272
rect 37419 2069 37449 2272
rect 37510 2071 37576 2087
rect 37510 2069 37526 2071
rect 37419 2039 37526 2069
rect 37510 2037 37526 2039
rect 37560 2037 37576 2071
rect 37510 2021 37576 2037
rect 37306 1867 37372 1883
rect 37306 1865 37322 1867
rect 37215 1835 37322 1865
rect 37306 1833 37322 1835
rect 37356 1833 37372 1867
rect 37306 1817 37372 1833
rect 37102 1663 37168 1679
rect 37102 1661 37118 1663
rect 37011 1631 37118 1661
rect 37102 1629 37118 1631
rect 37152 1629 37168 1663
rect 37102 1613 37168 1629
rect 36898 1459 36964 1475
rect 36898 1457 36914 1459
rect 36807 1427 36914 1457
rect 36898 1425 36914 1427
rect 36948 1425 36964 1459
rect 36898 1409 36964 1425
rect 36694 1255 36760 1271
rect 36694 1253 36710 1255
rect 36603 1223 36710 1253
rect 36694 1221 36710 1223
rect 36744 1221 36760 1255
rect 36694 1205 36760 1221
rect 36490 1051 36556 1067
rect 36490 1049 36506 1051
rect 36399 1019 36506 1049
rect 36490 1017 36506 1019
rect 36540 1017 36556 1051
rect 36490 1001 36556 1017
rect 36286 847 36352 863
rect 36286 845 36302 847
rect 36195 815 36302 845
rect 36286 813 36302 815
rect 36336 813 36352 847
rect 36286 797 36352 813
rect 36082 643 36148 659
rect 36082 641 36098 643
rect 35991 611 36098 641
rect 34450 593 34516 609
rect 36082 609 36098 611
rect 36132 609 36148 643
rect 37623 641 37653 2272
rect 37827 845 37857 2272
rect 38031 1049 38061 2272
rect 38235 1253 38265 2272
rect 38439 1457 38469 2272
rect 38643 1661 38673 2272
rect 38847 1865 38877 2272
rect 39051 2069 39081 2272
rect 39142 2071 39208 2087
rect 39142 2069 39158 2071
rect 39051 2039 39158 2069
rect 39142 2037 39158 2039
rect 39192 2037 39208 2071
rect 39142 2021 39208 2037
rect 38938 1867 39004 1883
rect 38938 1865 38954 1867
rect 38847 1835 38954 1865
rect 38938 1833 38954 1835
rect 38988 1833 39004 1867
rect 38938 1817 39004 1833
rect 38734 1663 38800 1679
rect 38734 1661 38750 1663
rect 38643 1631 38750 1661
rect 38734 1629 38750 1631
rect 38784 1629 38800 1663
rect 38734 1613 38800 1629
rect 38530 1459 38596 1475
rect 38530 1457 38546 1459
rect 38439 1427 38546 1457
rect 38530 1425 38546 1427
rect 38580 1425 38596 1459
rect 38530 1409 38596 1425
rect 38326 1255 38392 1271
rect 38326 1253 38342 1255
rect 38235 1223 38342 1253
rect 38326 1221 38342 1223
rect 38376 1221 38392 1255
rect 38326 1205 38392 1221
rect 38122 1051 38188 1067
rect 38122 1049 38138 1051
rect 38031 1019 38138 1049
rect 38122 1017 38138 1019
rect 38172 1017 38188 1051
rect 38122 1001 38188 1017
rect 37918 847 37984 863
rect 37918 845 37934 847
rect 37827 815 37934 845
rect 37918 813 37934 815
rect 37968 813 37984 847
rect 37918 797 37984 813
rect 37714 643 37780 659
rect 37714 641 37730 643
rect 37623 611 37730 641
rect 36082 593 36148 609
rect 37714 609 37730 611
rect 37764 609 37780 643
rect 39255 641 39285 2272
rect 39459 845 39489 2272
rect 39663 1049 39693 2272
rect 39867 1253 39897 2272
rect 40071 1457 40101 2272
rect 40275 1661 40305 2272
rect 40479 1865 40509 2272
rect 40683 2069 40713 2272
rect 40774 2071 40840 2087
rect 40774 2069 40790 2071
rect 40683 2039 40790 2069
rect 40774 2037 40790 2039
rect 40824 2037 40840 2071
rect 40774 2021 40840 2037
rect 40570 1867 40636 1883
rect 40570 1865 40586 1867
rect 40479 1835 40586 1865
rect 40570 1833 40586 1835
rect 40620 1833 40636 1867
rect 40570 1817 40636 1833
rect 40366 1663 40432 1679
rect 40366 1661 40382 1663
rect 40275 1631 40382 1661
rect 40366 1629 40382 1631
rect 40416 1629 40432 1663
rect 40366 1613 40432 1629
rect 40162 1459 40228 1475
rect 40162 1457 40178 1459
rect 40071 1427 40178 1457
rect 40162 1425 40178 1427
rect 40212 1425 40228 1459
rect 40162 1409 40228 1425
rect 39958 1255 40024 1271
rect 39958 1253 39974 1255
rect 39867 1223 39974 1253
rect 39958 1221 39974 1223
rect 40008 1221 40024 1255
rect 39958 1205 40024 1221
rect 39754 1051 39820 1067
rect 39754 1049 39770 1051
rect 39663 1019 39770 1049
rect 39754 1017 39770 1019
rect 39804 1017 39820 1051
rect 39754 1001 39820 1017
rect 39550 847 39616 863
rect 39550 845 39566 847
rect 39459 815 39566 845
rect 39550 813 39566 815
rect 39600 813 39616 847
rect 39550 797 39616 813
rect 39346 643 39412 659
rect 39346 641 39362 643
rect 39255 611 39362 641
rect 37714 593 37780 609
rect 39346 609 39362 611
rect 39396 609 39412 643
rect 40887 641 40917 2272
rect 41091 845 41121 2272
rect 41295 1049 41325 2272
rect 41499 1253 41529 2272
rect 41703 1457 41733 2272
rect 41907 1661 41937 2272
rect 42111 1865 42141 2272
rect 42315 2069 42345 2272
rect 42406 2071 42472 2087
rect 42406 2069 42422 2071
rect 42315 2039 42422 2069
rect 42406 2037 42422 2039
rect 42456 2037 42472 2071
rect 42406 2021 42472 2037
rect 42202 1867 42268 1883
rect 42202 1865 42218 1867
rect 42111 1835 42218 1865
rect 42202 1833 42218 1835
rect 42252 1833 42268 1867
rect 42202 1817 42268 1833
rect 41998 1663 42064 1679
rect 41998 1661 42014 1663
rect 41907 1631 42014 1661
rect 41998 1629 42014 1631
rect 42048 1629 42064 1663
rect 41998 1613 42064 1629
rect 41794 1459 41860 1475
rect 41794 1457 41810 1459
rect 41703 1427 41810 1457
rect 41794 1425 41810 1427
rect 41844 1425 41860 1459
rect 41794 1409 41860 1425
rect 41590 1255 41656 1271
rect 41590 1253 41606 1255
rect 41499 1223 41606 1253
rect 41590 1221 41606 1223
rect 41640 1221 41656 1255
rect 41590 1205 41656 1221
rect 41386 1051 41452 1067
rect 41386 1049 41402 1051
rect 41295 1019 41402 1049
rect 41386 1017 41402 1019
rect 41436 1017 41452 1051
rect 41386 1001 41452 1017
rect 41182 847 41248 863
rect 41182 845 41198 847
rect 41091 815 41198 845
rect 41182 813 41198 815
rect 41232 813 41248 847
rect 41182 797 41248 813
rect 40978 643 41044 659
rect 40978 641 40994 643
rect 40887 611 40994 641
rect 39346 593 39412 609
rect 40978 609 40994 611
rect 41028 609 41044 643
rect 42519 641 42549 2272
rect 42723 845 42753 2272
rect 42927 1049 42957 2272
rect 43131 1253 43161 2272
rect 43335 1457 43365 2272
rect 43539 1661 43569 2272
rect 43743 1865 43773 2272
rect 43947 2069 43977 2272
rect 44038 2071 44104 2087
rect 44038 2069 44054 2071
rect 43947 2039 44054 2069
rect 44038 2037 44054 2039
rect 44088 2037 44104 2071
rect 44038 2021 44104 2037
rect 43834 1867 43900 1883
rect 43834 1865 43850 1867
rect 43743 1835 43850 1865
rect 43834 1833 43850 1835
rect 43884 1833 43900 1867
rect 43834 1817 43900 1833
rect 43630 1663 43696 1679
rect 43630 1661 43646 1663
rect 43539 1631 43646 1661
rect 43630 1629 43646 1631
rect 43680 1629 43696 1663
rect 43630 1613 43696 1629
rect 43426 1459 43492 1475
rect 43426 1457 43442 1459
rect 43335 1427 43442 1457
rect 43426 1425 43442 1427
rect 43476 1425 43492 1459
rect 43426 1409 43492 1425
rect 43222 1255 43288 1271
rect 43222 1253 43238 1255
rect 43131 1223 43238 1253
rect 43222 1221 43238 1223
rect 43272 1221 43288 1255
rect 43222 1205 43288 1221
rect 43018 1051 43084 1067
rect 43018 1049 43034 1051
rect 42927 1019 43034 1049
rect 43018 1017 43034 1019
rect 43068 1017 43084 1051
rect 43018 1001 43084 1017
rect 42814 847 42880 863
rect 42814 845 42830 847
rect 42723 815 42830 845
rect 42814 813 42830 815
rect 42864 813 42880 847
rect 42814 797 42880 813
rect 42610 643 42676 659
rect 42610 641 42626 643
rect 42519 611 42626 641
rect 40978 593 41044 609
rect 42610 609 42626 611
rect 42660 609 42676 643
rect 44151 641 44181 2272
rect 44355 845 44385 2272
rect 44559 1049 44589 2272
rect 44763 1253 44793 2272
rect 44967 1457 44997 2272
rect 45171 1661 45201 2272
rect 45375 1865 45405 2272
rect 45579 2069 45609 2272
rect 45670 2071 45736 2087
rect 45670 2069 45686 2071
rect 45579 2039 45686 2069
rect 45670 2037 45686 2039
rect 45720 2037 45736 2071
rect 45670 2021 45736 2037
rect 45466 1867 45532 1883
rect 45466 1865 45482 1867
rect 45375 1835 45482 1865
rect 45466 1833 45482 1835
rect 45516 1833 45532 1867
rect 45466 1817 45532 1833
rect 45262 1663 45328 1679
rect 45262 1661 45278 1663
rect 45171 1631 45278 1661
rect 45262 1629 45278 1631
rect 45312 1629 45328 1663
rect 45262 1613 45328 1629
rect 45058 1459 45124 1475
rect 45058 1457 45074 1459
rect 44967 1427 45074 1457
rect 45058 1425 45074 1427
rect 45108 1425 45124 1459
rect 45058 1409 45124 1425
rect 44854 1255 44920 1271
rect 44854 1253 44870 1255
rect 44763 1223 44870 1253
rect 44854 1221 44870 1223
rect 44904 1221 44920 1255
rect 44854 1205 44920 1221
rect 44650 1051 44716 1067
rect 44650 1049 44666 1051
rect 44559 1019 44666 1049
rect 44650 1017 44666 1019
rect 44700 1017 44716 1051
rect 44650 1001 44716 1017
rect 44446 847 44512 863
rect 44446 845 44462 847
rect 44355 815 44462 845
rect 44446 813 44462 815
rect 44496 813 44512 847
rect 44446 797 44512 813
rect 44242 643 44308 659
rect 44242 641 44258 643
rect 44151 611 44258 641
rect 42610 593 42676 609
rect 44242 609 44258 611
rect 44292 609 44308 643
rect 45783 641 45813 2272
rect 45987 845 46017 2272
rect 46191 1049 46221 2272
rect 46395 1253 46425 2272
rect 46599 1457 46629 2272
rect 46803 1661 46833 2272
rect 47007 1865 47037 2272
rect 47211 2069 47241 2272
rect 47302 2071 47368 2087
rect 47302 2069 47318 2071
rect 47211 2039 47318 2069
rect 47302 2037 47318 2039
rect 47352 2037 47368 2071
rect 47302 2021 47368 2037
rect 47098 1867 47164 1883
rect 47098 1865 47114 1867
rect 47007 1835 47114 1865
rect 47098 1833 47114 1835
rect 47148 1833 47164 1867
rect 47098 1817 47164 1833
rect 46894 1663 46960 1679
rect 46894 1661 46910 1663
rect 46803 1631 46910 1661
rect 46894 1629 46910 1631
rect 46944 1629 46960 1663
rect 46894 1613 46960 1629
rect 46690 1459 46756 1475
rect 46690 1457 46706 1459
rect 46599 1427 46706 1457
rect 46690 1425 46706 1427
rect 46740 1425 46756 1459
rect 46690 1409 46756 1425
rect 46486 1255 46552 1271
rect 46486 1253 46502 1255
rect 46395 1223 46502 1253
rect 46486 1221 46502 1223
rect 46536 1221 46552 1255
rect 46486 1205 46552 1221
rect 46282 1051 46348 1067
rect 46282 1049 46298 1051
rect 46191 1019 46298 1049
rect 46282 1017 46298 1019
rect 46332 1017 46348 1051
rect 46282 1001 46348 1017
rect 46078 847 46144 863
rect 46078 845 46094 847
rect 45987 815 46094 845
rect 46078 813 46094 815
rect 46128 813 46144 847
rect 46078 797 46144 813
rect 45874 643 45940 659
rect 45874 641 45890 643
rect 45783 611 45890 641
rect 44242 593 44308 609
rect 45874 609 45890 611
rect 45924 609 45940 643
rect 47415 641 47445 2272
rect 47619 845 47649 2272
rect 47823 1049 47853 2272
rect 48027 1253 48057 2272
rect 48231 1457 48261 2272
rect 48435 1661 48465 2272
rect 48639 1865 48669 2272
rect 48843 2069 48873 2272
rect 48934 2071 49000 2087
rect 48934 2069 48950 2071
rect 48843 2039 48950 2069
rect 48934 2037 48950 2039
rect 48984 2037 49000 2071
rect 48934 2021 49000 2037
rect 48730 1867 48796 1883
rect 48730 1865 48746 1867
rect 48639 1835 48746 1865
rect 48730 1833 48746 1835
rect 48780 1833 48796 1867
rect 48730 1817 48796 1833
rect 48526 1663 48592 1679
rect 48526 1661 48542 1663
rect 48435 1631 48542 1661
rect 48526 1629 48542 1631
rect 48576 1629 48592 1663
rect 48526 1613 48592 1629
rect 48322 1459 48388 1475
rect 48322 1457 48338 1459
rect 48231 1427 48338 1457
rect 48322 1425 48338 1427
rect 48372 1425 48388 1459
rect 48322 1409 48388 1425
rect 48118 1255 48184 1271
rect 48118 1253 48134 1255
rect 48027 1223 48134 1253
rect 48118 1221 48134 1223
rect 48168 1221 48184 1255
rect 48118 1205 48184 1221
rect 47914 1051 47980 1067
rect 47914 1049 47930 1051
rect 47823 1019 47930 1049
rect 47914 1017 47930 1019
rect 47964 1017 47980 1051
rect 47914 1001 47980 1017
rect 47710 847 47776 863
rect 47710 845 47726 847
rect 47619 815 47726 845
rect 47710 813 47726 815
rect 47760 813 47776 847
rect 47710 797 47776 813
rect 47506 643 47572 659
rect 47506 641 47522 643
rect 47415 611 47522 641
rect 45874 593 45940 609
rect 47506 609 47522 611
rect 47556 609 47572 643
rect 49047 641 49077 2272
rect 49251 845 49281 2272
rect 49455 1049 49485 2272
rect 49659 1253 49689 2272
rect 49863 1457 49893 2272
rect 50067 1661 50097 2272
rect 50271 1865 50301 2272
rect 50475 2069 50505 2272
rect 50566 2071 50632 2087
rect 50566 2069 50582 2071
rect 50475 2039 50582 2069
rect 50566 2037 50582 2039
rect 50616 2037 50632 2071
rect 50566 2021 50632 2037
rect 50362 1867 50428 1883
rect 50362 1865 50378 1867
rect 50271 1835 50378 1865
rect 50362 1833 50378 1835
rect 50412 1833 50428 1867
rect 50362 1817 50428 1833
rect 50158 1663 50224 1679
rect 50158 1661 50174 1663
rect 50067 1631 50174 1661
rect 50158 1629 50174 1631
rect 50208 1629 50224 1663
rect 50158 1613 50224 1629
rect 49954 1459 50020 1475
rect 49954 1457 49970 1459
rect 49863 1427 49970 1457
rect 49954 1425 49970 1427
rect 50004 1425 50020 1459
rect 49954 1409 50020 1425
rect 49750 1255 49816 1271
rect 49750 1253 49766 1255
rect 49659 1223 49766 1253
rect 49750 1221 49766 1223
rect 49800 1221 49816 1255
rect 49750 1205 49816 1221
rect 49546 1051 49612 1067
rect 49546 1049 49562 1051
rect 49455 1019 49562 1049
rect 49546 1017 49562 1019
rect 49596 1017 49612 1051
rect 49546 1001 49612 1017
rect 49342 847 49408 863
rect 49342 845 49358 847
rect 49251 815 49358 845
rect 49342 813 49358 815
rect 49392 813 49408 847
rect 49342 797 49408 813
rect 49138 643 49204 659
rect 49138 641 49154 643
rect 49047 611 49154 641
rect 47506 593 47572 609
rect 49138 609 49154 611
rect 49188 609 49204 643
rect 50679 641 50709 2272
rect 50883 845 50913 2272
rect 51087 1049 51117 2272
rect 51291 1253 51321 2272
rect 51495 1457 51525 2272
rect 51699 1661 51729 2272
rect 51903 1865 51933 2272
rect 52107 2069 52137 2272
rect 52198 2071 52264 2087
rect 52198 2069 52214 2071
rect 52107 2039 52214 2069
rect 52198 2037 52214 2039
rect 52248 2037 52264 2071
rect 52198 2021 52264 2037
rect 51994 1867 52060 1883
rect 51994 1865 52010 1867
rect 51903 1835 52010 1865
rect 51994 1833 52010 1835
rect 52044 1833 52060 1867
rect 51994 1817 52060 1833
rect 51790 1663 51856 1679
rect 51790 1661 51806 1663
rect 51699 1631 51806 1661
rect 51790 1629 51806 1631
rect 51840 1629 51856 1663
rect 51790 1613 51856 1629
rect 51586 1459 51652 1475
rect 51586 1457 51602 1459
rect 51495 1427 51602 1457
rect 51586 1425 51602 1427
rect 51636 1425 51652 1459
rect 51586 1409 51652 1425
rect 51382 1255 51448 1271
rect 51382 1253 51398 1255
rect 51291 1223 51398 1253
rect 51382 1221 51398 1223
rect 51432 1221 51448 1255
rect 51382 1205 51448 1221
rect 51178 1051 51244 1067
rect 51178 1049 51194 1051
rect 51087 1019 51194 1049
rect 51178 1017 51194 1019
rect 51228 1017 51244 1051
rect 51178 1001 51244 1017
rect 50974 847 51040 863
rect 50974 845 50990 847
rect 50883 815 50990 845
rect 50974 813 50990 815
rect 51024 813 51040 847
rect 50974 797 51040 813
rect 50770 643 50836 659
rect 50770 641 50786 643
rect 50679 611 50786 641
rect 49138 593 49204 609
rect 50770 609 50786 611
rect 50820 609 50836 643
rect 50770 593 50836 609
<< polycont >>
rect 1622 2037 1656 2071
rect 1418 1833 1452 1867
rect 1214 1629 1248 1663
rect 1010 1425 1044 1459
rect 806 1221 840 1255
rect 602 1017 636 1051
rect 398 813 432 847
rect 194 609 228 643
rect 3254 2037 3288 2071
rect 3050 1833 3084 1867
rect 2846 1629 2880 1663
rect 2642 1425 2676 1459
rect 2438 1221 2472 1255
rect 2234 1017 2268 1051
rect 2030 813 2064 847
rect 1826 609 1860 643
rect 4886 2037 4920 2071
rect 4682 1833 4716 1867
rect 4478 1629 4512 1663
rect 4274 1425 4308 1459
rect 4070 1221 4104 1255
rect 3866 1017 3900 1051
rect 3662 813 3696 847
rect 3458 609 3492 643
rect 6518 2037 6552 2071
rect 6314 1833 6348 1867
rect 6110 1629 6144 1663
rect 5906 1425 5940 1459
rect 5702 1221 5736 1255
rect 5498 1017 5532 1051
rect 5294 813 5328 847
rect 5090 609 5124 643
rect 8150 2037 8184 2071
rect 7946 1833 7980 1867
rect 7742 1629 7776 1663
rect 7538 1425 7572 1459
rect 7334 1221 7368 1255
rect 7130 1017 7164 1051
rect 6926 813 6960 847
rect 6722 609 6756 643
rect 9782 2037 9816 2071
rect 9578 1833 9612 1867
rect 9374 1629 9408 1663
rect 9170 1425 9204 1459
rect 8966 1221 9000 1255
rect 8762 1017 8796 1051
rect 8558 813 8592 847
rect 8354 609 8388 643
rect 11414 2037 11448 2071
rect 11210 1833 11244 1867
rect 11006 1629 11040 1663
rect 10802 1425 10836 1459
rect 10598 1221 10632 1255
rect 10394 1017 10428 1051
rect 10190 813 10224 847
rect 9986 609 10020 643
rect 13046 2037 13080 2071
rect 12842 1833 12876 1867
rect 12638 1629 12672 1663
rect 12434 1425 12468 1459
rect 12230 1221 12264 1255
rect 12026 1017 12060 1051
rect 11822 813 11856 847
rect 11618 609 11652 643
rect 14678 2037 14712 2071
rect 14474 1833 14508 1867
rect 14270 1629 14304 1663
rect 14066 1425 14100 1459
rect 13862 1221 13896 1255
rect 13658 1017 13692 1051
rect 13454 813 13488 847
rect 13250 609 13284 643
rect 16310 2037 16344 2071
rect 16106 1833 16140 1867
rect 15902 1629 15936 1663
rect 15698 1425 15732 1459
rect 15494 1221 15528 1255
rect 15290 1017 15324 1051
rect 15086 813 15120 847
rect 14882 609 14916 643
rect 17942 2037 17976 2071
rect 17738 1833 17772 1867
rect 17534 1629 17568 1663
rect 17330 1425 17364 1459
rect 17126 1221 17160 1255
rect 16922 1017 16956 1051
rect 16718 813 16752 847
rect 16514 609 16548 643
rect 19574 2037 19608 2071
rect 19370 1833 19404 1867
rect 19166 1629 19200 1663
rect 18962 1425 18996 1459
rect 18758 1221 18792 1255
rect 18554 1017 18588 1051
rect 18350 813 18384 847
rect 18146 609 18180 643
rect 21206 2037 21240 2071
rect 21002 1833 21036 1867
rect 20798 1629 20832 1663
rect 20594 1425 20628 1459
rect 20390 1221 20424 1255
rect 20186 1017 20220 1051
rect 19982 813 20016 847
rect 19778 609 19812 643
rect 22838 2037 22872 2071
rect 22634 1833 22668 1867
rect 22430 1629 22464 1663
rect 22226 1425 22260 1459
rect 22022 1221 22056 1255
rect 21818 1017 21852 1051
rect 21614 813 21648 847
rect 21410 609 21444 643
rect 24470 2037 24504 2071
rect 24266 1833 24300 1867
rect 24062 1629 24096 1663
rect 23858 1425 23892 1459
rect 23654 1221 23688 1255
rect 23450 1017 23484 1051
rect 23246 813 23280 847
rect 23042 609 23076 643
rect 26102 2037 26136 2071
rect 25898 1833 25932 1867
rect 25694 1629 25728 1663
rect 25490 1425 25524 1459
rect 25286 1221 25320 1255
rect 25082 1017 25116 1051
rect 24878 813 24912 847
rect 24674 609 24708 643
rect 27734 2037 27768 2071
rect 27530 1833 27564 1867
rect 27326 1629 27360 1663
rect 27122 1425 27156 1459
rect 26918 1221 26952 1255
rect 26714 1017 26748 1051
rect 26510 813 26544 847
rect 26306 609 26340 643
rect 29366 2037 29400 2071
rect 29162 1833 29196 1867
rect 28958 1629 28992 1663
rect 28754 1425 28788 1459
rect 28550 1221 28584 1255
rect 28346 1017 28380 1051
rect 28142 813 28176 847
rect 27938 609 27972 643
rect 30998 2037 31032 2071
rect 30794 1833 30828 1867
rect 30590 1629 30624 1663
rect 30386 1425 30420 1459
rect 30182 1221 30216 1255
rect 29978 1017 30012 1051
rect 29774 813 29808 847
rect 29570 609 29604 643
rect 32630 2037 32664 2071
rect 32426 1833 32460 1867
rect 32222 1629 32256 1663
rect 32018 1425 32052 1459
rect 31814 1221 31848 1255
rect 31610 1017 31644 1051
rect 31406 813 31440 847
rect 31202 609 31236 643
rect 34262 2037 34296 2071
rect 34058 1833 34092 1867
rect 33854 1629 33888 1663
rect 33650 1425 33684 1459
rect 33446 1221 33480 1255
rect 33242 1017 33276 1051
rect 33038 813 33072 847
rect 32834 609 32868 643
rect 35894 2037 35928 2071
rect 35690 1833 35724 1867
rect 35486 1629 35520 1663
rect 35282 1425 35316 1459
rect 35078 1221 35112 1255
rect 34874 1017 34908 1051
rect 34670 813 34704 847
rect 34466 609 34500 643
rect 37526 2037 37560 2071
rect 37322 1833 37356 1867
rect 37118 1629 37152 1663
rect 36914 1425 36948 1459
rect 36710 1221 36744 1255
rect 36506 1017 36540 1051
rect 36302 813 36336 847
rect 36098 609 36132 643
rect 39158 2037 39192 2071
rect 38954 1833 38988 1867
rect 38750 1629 38784 1663
rect 38546 1425 38580 1459
rect 38342 1221 38376 1255
rect 38138 1017 38172 1051
rect 37934 813 37968 847
rect 37730 609 37764 643
rect 40790 2037 40824 2071
rect 40586 1833 40620 1867
rect 40382 1629 40416 1663
rect 40178 1425 40212 1459
rect 39974 1221 40008 1255
rect 39770 1017 39804 1051
rect 39566 813 39600 847
rect 39362 609 39396 643
rect 42422 2037 42456 2071
rect 42218 1833 42252 1867
rect 42014 1629 42048 1663
rect 41810 1425 41844 1459
rect 41606 1221 41640 1255
rect 41402 1017 41436 1051
rect 41198 813 41232 847
rect 40994 609 41028 643
rect 44054 2037 44088 2071
rect 43850 1833 43884 1867
rect 43646 1629 43680 1663
rect 43442 1425 43476 1459
rect 43238 1221 43272 1255
rect 43034 1017 43068 1051
rect 42830 813 42864 847
rect 42626 609 42660 643
rect 45686 2037 45720 2071
rect 45482 1833 45516 1867
rect 45278 1629 45312 1663
rect 45074 1425 45108 1459
rect 44870 1221 44904 1255
rect 44666 1017 44700 1051
rect 44462 813 44496 847
rect 44258 609 44292 643
rect 47318 2037 47352 2071
rect 47114 1833 47148 1867
rect 46910 1629 46944 1663
rect 46706 1425 46740 1459
rect 46502 1221 46536 1255
rect 46298 1017 46332 1051
rect 46094 813 46128 847
rect 45890 609 45924 643
rect 48950 2037 48984 2071
rect 48746 1833 48780 1867
rect 48542 1629 48576 1663
rect 48338 1425 48372 1459
rect 48134 1221 48168 1255
rect 47930 1017 47964 1051
rect 47726 813 47760 847
rect 47522 609 47556 643
rect 50582 2037 50616 2071
rect 50378 1833 50412 1867
rect 50174 1629 50208 1663
rect 49970 1425 50004 1459
rect 49766 1221 49800 1255
rect 49562 1017 49596 1051
rect 49358 813 49392 847
rect 49154 609 49188 643
rect 52214 2037 52248 2071
rect 52010 1833 52044 1867
rect 51806 1629 51840 1663
rect 51602 1425 51636 1459
rect 51398 1221 51432 1255
rect 51194 1017 51228 1051
rect 50990 813 51024 847
rect 50786 609 50820 643
<< locali >>
rect 1606 2037 1622 2071
rect 1656 2037 1672 2071
rect 3238 2037 3254 2071
rect 3288 2037 3304 2071
rect 4870 2037 4886 2071
rect 4920 2037 4936 2071
rect 6502 2037 6518 2071
rect 6552 2037 6568 2071
rect 8134 2037 8150 2071
rect 8184 2037 8200 2071
rect 9766 2037 9782 2071
rect 9816 2037 9832 2071
rect 11398 2037 11414 2071
rect 11448 2037 11464 2071
rect 13030 2037 13046 2071
rect 13080 2037 13096 2071
rect 14662 2037 14678 2071
rect 14712 2037 14728 2071
rect 16294 2037 16310 2071
rect 16344 2037 16360 2071
rect 17926 2037 17942 2071
rect 17976 2037 17992 2071
rect 19558 2037 19574 2071
rect 19608 2037 19624 2071
rect 21190 2037 21206 2071
rect 21240 2037 21256 2071
rect 22822 2037 22838 2071
rect 22872 2037 22888 2071
rect 24454 2037 24470 2071
rect 24504 2037 24520 2071
rect 26086 2037 26102 2071
rect 26136 2037 26152 2071
rect 27718 2037 27734 2071
rect 27768 2037 27784 2071
rect 29350 2037 29366 2071
rect 29400 2037 29416 2071
rect 30982 2037 30998 2071
rect 31032 2037 31048 2071
rect 32614 2037 32630 2071
rect 32664 2037 32680 2071
rect 34246 2037 34262 2071
rect 34296 2037 34312 2071
rect 35878 2037 35894 2071
rect 35928 2037 35944 2071
rect 37510 2037 37526 2071
rect 37560 2037 37576 2071
rect 39142 2037 39158 2071
rect 39192 2037 39208 2071
rect 40774 2037 40790 2071
rect 40824 2037 40840 2071
rect 42406 2037 42422 2071
rect 42456 2037 42472 2071
rect 44038 2037 44054 2071
rect 44088 2037 44104 2071
rect 45670 2037 45686 2071
rect 45720 2037 45736 2071
rect 47302 2037 47318 2071
rect 47352 2037 47368 2071
rect 48934 2037 48950 2071
rect 48984 2037 49000 2071
rect 50566 2037 50582 2071
rect 50616 2037 50632 2071
rect 52198 2037 52214 2071
rect 52248 2037 52264 2071
rect 1402 1833 1418 1867
rect 1452 1833 1468 1867
rect 3034 1833 3050 1867
rect 3084 1833 3100 1867
rect 4666 1833 4682 1867
rect 4716 1833 4732 1867
rect 6298 1833 6314 1867
rect 6348 1833 6364 1867
rect 7930 1833 7946 1867
rect 7980 1833 7996 1867
rect 9562 1833 9578 1867
rect 9612 1833 9628 1867
rect 11194 1833 11210 1867
rect 11244 1833 11260 1867
rect 12826 1833 12842 1867
rect 12876 1833 12892 1867
rect 14458 1833 14474 1867
rect 14508 1833 14524 1867
rect 16090 1833 16106 1867
rect 16140 1833 16156 1867
rect 17722 1833 17738 1867
rect 17772 1833 17788 1867
rect 19354 1833 19370 1867
rect 19404 1833 19420 1867
rect 20986 1833 21002 1867
rect 21036 1833 21052 1867
rect 22618 1833 22634 1867
rect 22668 1833 22684 1867
rect 24250 1833 24266 1867
rect 24300 1833 24316 1867
rect 25882 1833 25898 1867
rect 25932 1833 25948 1867
rect 27514 1833 27530 1867
rect 27564 1833 27580 1867
rect 29146 1833 29162 1867
rect 29196 1833 29212 1867
rect 30778 1833 30794 1867
rect 30828 1833 30844 1867
rect 32410 1833 32426 1867
rect 32460 1833 32476 1867
rect 34042 1833 34058 1867
rect 34092 1833 34108 1867
rect 35674 1833 35690 1867
rect 35724 1833 35740 1867
rect 37306 1833 37322 1867
rect 37356 1833 37372 1867
rect 38938 1833 38954 1867
rect 38988 1833 39004 1867
rect 40570 1833 40586 1867
rect 40620 1833 40636 1867
rect 42202 1833 42218 1867
rect 42252 1833 42268 1867
rect 43834 1833 43850 1867
rect 43884 1833 43900 1867
rect 45466 1833 45482 1867
rect 45516 1833 45532 1867
rect 47098 1833 47114 1867
rect 47148 1833 47164 1867
rect 48730 1833 48746 1867
rect 48780 1833 48796 1867
rect 50362 1833 50378 1867
rect 50412 1833 50428 1867
rect 51994 1833 52010 1867
rect 52044 1833 52060 1867
rect 1198 1629 1214 1663
rect 1248 1629 1264 1663
rect 2830 1629 2846 1663
rect 2880 1629 2896 1663
rect 4462 1629 4478 1663
rect 4512 1629 4528 1663
rect 6094 1629 6110 1663
rect 6144 1629 6160 1663
rect 7726 1629 7742 1663
rect 7776 1629 7792 1663
rect 9358 1629 9374 1663
rect 9408 1629 9424 1663
rect 10990 1629 11006 1663
rect 11040 1629 11056 1663
rect 12622 1629 12638 1663
rect 12672 1629 12688 1663
rect 14254 1629 14270 1663
rect 14304 1629 14320 1663
rect 15886 1629 15902 1663
rect 15936 1629 15952 1663
rect 17518 1629 17534 1663
rect 17568 1629 17584 1663
rect 19150 1629 19166 1663
rect 19200 1629 19216 1663
rect 20782 1629 20798 1663
rect 20832 1629 20848 1663
rect 22414 1629 22430 1663
rect 22464 1629 22480 1663
rect 24046 1629 24062 1663
rect 24096 1629 24112 1663
rect 25678 1629 25694 1663
rect 25728 1629 25744 1663
rect 27310 1629 27326 1663
rect 27360 1629 27376 1663
rect 28942 1629 28958 1663
rect 28992 1629 29008 1663
rect 30574 1629 30590 1663
rect 30624 1629 30640 1663
rect 32206 1629 32222 1663
rect 32256 1629 32272 1663
rect 33838 1629 33854 1663
rect 33888 1629 33904 1663
rect 35470 1629 35486 1663
rect 35520 1629 35536 1663
rect 37102 1629 37118 1663
rect 37152 1629 37168 1663
rect 38734 1629 38750 1663
rect 38784 1629 38800 1663
rect 40366 1629 40382 1663
rect 40416 1629 40432 1663
rect 41998 1629 42014 1663
rect 42048 1629 42064 1663
rect 43630 1629 43646 1663
rect 43680 1629 43696 1663
rect 45262 1629 45278 1663
rect 45312 1629 45328 1663
rect 46894 1629 46910 1663
rect 46944 1629 46960 1663
rect 48526 1629 48542 1663
rect 48576 1629 48592 1663
rect 50158 1629 50174 1663
rect 50208 1629 50224 1663
rect 51790 1629 51806 1663
rect 51840 1629 51856 1663
rect 994 1425 1010 1459
rect 1044 1425 1060 1459
rect 2626 1425 2642 1459
rect 2676 1425 2692 1459
rect 4258 1425 4274 1459
rect 4308 1425 4324 1459
rect 5890 1425 5906 1459
rect 5940 1425 5956 1459
rect 7522 1425 7538 1459
rect 7572 1425 7588 1459
rect 9154 1425 9170 1459
rect 9204 1425 9220 1459
rect 10786 1425 10802 1459
rect 10836 1425 10852 1459
rect 12418 1425 12434 1459
rect 12468 1425 12484 1459
rect 14050 1425 14066 1459
rect 14100 1425 14116 1459
rect 15682 1425 15698 1459
rect 15732 1425 15748 1459
rect 17314 1425 17330 1459
rect 17364 1425 17380 1459
rect 18946 1425 18962 1459
rect 18996 1425 19012 1459
rect 20578 1425 20594 1459
rect 20628 1425 20644 1459
rect 22210 1425 22226 1459
rect 22260 1425 22276 1459
rect 23842 1425 23858 1459
rect 23892 1425 23908 1459
rect 25474 1425 25490 1459
rect 25524 1425 25540 1459
rect 27106 1425 27122 1459
rect 27156 1425 27172 1459
rect 28738 1425 28754 1459
rect 28788 1425 28804 1459
rect 30370 1425 30386 1459
rect 30420 1425 30436 1459
rect 32002 1425 32018 1459
rect 32052 1425 32068 1459
rect 33634 1425 33650 1459
rect 33684 1425 33700 1459
rect 35266 1425 35282 1459
rect 35316 1425 35332 1459
rect 36898 1425 36914 1459
rect 36948 1425 36964 1459
rect 38530 1425 38546 1459
rect 38580 1425 38596 1459
rect 40162 1425 40178 1459
rect 40212 1425 40228 1459
rect 41794 1425 41810 1459
rect 41844 1425 41860 1459
rect 43426 1425 43442 1459
rect 43476 1425 43492 1459
rect 45058 1425 45074 1459
rect 45108 1425 45124 1459
rect 46690 1425 46706 1459
rect 46740 1425 46756 1459
rect 48322 1425 48338 1459
rect 48372 1425 48388 1459
rect 49954 1425 49970 1459
rect 50004 1425 50020 1459
rect 51586 1425 51602 1459
rect 51636 1425 51652 1459
rect 790 1221 806 1255
rect 840 1221 856 1255
rect 2422 1221 2438 1255
rect 2472 1221 2488 1255
rect 4054 1221 4070 1255
rect 4104 1221 4120 1255
rect 5686 1221 5702 1255
rect 5736 1221 5752 1255
rect 7318 1221 7334 1255
rect 7368 1221 7384 1255
rect 8950 1221 8966 1255
rect 9000 1221 9016 1255
rect 10582 1221 10598 1255
rect 10632 1221 10648 1255
rect 12214 1221 12230 1255
rect 12264 1221 12280 1255
rect 13846 1221 13862 1255
rect 13896 1221 13912 1255
rect 15478 1221 15494 1255
rect 15528 1221 15544 1255
rect 17110 1221 17126 1255
rect 17160 1221 17176 1255
rect 18742 1221 18758 1255
rect 18792 1221 18808 1255
rect 20374 1221 20390 1255
rect 20424 1221 20440 1255
rect 22006 1221 22022 1255
rect 22056 1221 22072 1255
rect 23638 1221 23654 1255
rect 23688 1221 23704 1255
rect 25270 1221 25286 1255
rect 25320 1221 25336 1255
rect 26902 1221 26918 1255
rect 26952 1221 26968 1255
rect 28534 1221 28550 1255
rect 28584 1221 28600 1255
rect 30166 1221 30182 1255
rect 30216 1221 30232 1255
rect 31798 1221 31814 1255
rect 31848 1221 31864 1255
rect 33430 1221 33446 1255
rect 33480 1221 33496 1255
rect 35062 1221 35078 1255
rect 35112 1221 35128 1255
rect 36694 1221 36710 1255
rect 36744 1221 36760 1255
rect 38326 1221 38342 1255
rect 38376 1221 38392 1255
rect 39958 1221 39974 1255
rect 40008 1221 40024 1255
rect 41590 1221 41606 1255
rect 41640 1221 41656 1255
rect 43222 1221 43238 1255
rect 43272 1221 43288 1255
rect 44854 1221 44870 1255
rect 44904 1221 44920 1255
rect 46486 1221 46502 1255
rect 46536 1221 46552 1255
rect 48118 1221 48134 1255
rect 48168 1221 48184 1255
rect 49750 1221 49766 1255
rect 49800 1221 49816 1255
rect 51382 1221 51398 1255
rect 51432 1221 51448 1255
rect 586 1017 602 1051
rect 636 1017 652 1051
rect 2218 1017 2234 1051
rect 2268 1017 2284 1051
rect 3850 1017 3866 1051
rect 3900 1017 3916 1051
rect 5482 1017 5498 1051
rect 5532 1017 5548 1051
rect 7114 1017 7130 1051
rect 7164 1017 7180 1051
rect 8746 1017 8762 1051
rect 8796 1017 8812 1051
rect 10378 1017 10394 1051
rect 10428 1017 10444 1051
rect 12010 1017 12026 1051
rect 12060 1017 12076 1051
rect 13642 1017 13658 1051
rect 13692 1017 13708 1051
rect 15274 1017 15290 1051
rect 15324 1017 15340 1051
rect 16906 1017 16922 1051
rect 16956 1017 16972 1051
rect 18538 1017 18554 1051
rect 18588 1017 18604 1051
rect 20170 1017 20186 1051
rect 20220 1017 20236 1051
rect 21802 1017 21818 1051
rect 21852 1017 21868 1051
rect 23434 1017 23450 1051
rect 23484 1017 23500 1051
rect 25066 1017 25082 1051
rect 25116 1017 25132 1051
rect 26698 1017 26714 1051
rect 26748 1017 26764 1051
rect 28330 1017 28346 1051
rect 28380 1017 28396 1051
rect 29962 1017 29978 1051
rect 30012 1017 30028 1051
rect 31594 1017 31610 1051
rect 31644 1017 31660 1051
rect 33226 1017 33242 1051
rect 33276 1017 33292 1051
rect 34858 1017 34874 1051
rect 34908 1017 34924 1051
rect 36490 1017 36506 1051
rect 36540 1017 36556 1051
rect 38122 1017 38138 1051
rect 38172 1017 38188 1051
rect 39754 1017 39770 1051
rect 39804 1017 39820 1051
rect 41386 1017 41402 1051
rect 41436 1017 41452 1051
rect 43018 1017 43034 1051
rect 43068 1017 43084 1051
rect 44650 1017 44666 1051
rect 44700 1017 44716 1051
rect 46282 1017 46298 1051
rect 46332 1017 46348 1051
rect 47914 1017 47930 1051
rect 47964 1017 47980 1051
rect 49546 1017 49562 1051
rect 49596 1017 49612 1051
rect 51178 1017 51194 1051
rect 51228 1017 51244 1051
rect 382 813 398 847
rect 432 813 448 847
rect 2014 813 2030 847
rect 2064 813 2080 847
rect 3646 813 3662 847
rect 3696 813 3712 847
rect 5278 813 5294 847
rect 5328 813 5344 847
rect 6910 813 6926 847
rect 6960 813 6976 847
rect 8542 813 8558 847
rect 8592 813 8608 847
rect 10174 813 10190 847
rect 10224 813 10240 847
rect 11806 813 11822 847
rect 11856 813 11872 847
rect 13438 813 13454 847
rect 13488 813 13504 847
rect 15070 813 15086 847
rect 15120 813 15136 847
rect 16702 813 16718 847
rect 16752 813 16768 847
rect 18334 813 18350 847
rect 18384 813 18400 847
rect 19966 813 19982 847
rect 20016 813 20032 847
rect 21598 813 21614 847
rect 21648 813 21664 847
rect 23230 813 23246 847
rect 23280 813 23296 847
rect 24862 813 24878 847
rect 24912 813 24928 847
rect 26494 813 26510 847
rect 26544 813 26560 847
rect 28126 813 28142 847
rect 28176 813 28192 847
rect 29758 813 29774 847
rect 29808 813 29824 847
rect 31390 813 31406 847
rect 31440 813 31456 847
rect 33022 813 33038 847
rect 33072 813 33088 847
rect 34654 813 34670 847
rect 34704 813 34720 847
rect 36286 813 36302 847
rect 36336 813 36352 847
rect 37918 813 37934 847
rect 37968 813 37984 847
rect 39550 813 39566 847
rect 39600 813 39616 847
rect 41182 813 41198 847
rect 41232 813 41248 847
rect 42814 813 42830 847
rect 42864 813 42880 847
rect 44446 813 44462 847
rect 44496 813 44512 847
rect 46078 813 46094 847
rect 46128 813 46144 847
rect 47710 813 47726 847
rect 47760 813 47776 847
rect 49342 813 49358 847
rect 49392 813 49408 847
rect 50974 813 50990 847
rect 51024 813 51040 847
rect 178 609 194 643
rect 228 609 244 643
rect 1810 609 1826 643
rect 1860 609 1876 643
rect 3442 609 3458 643
rect 3492 609 3508 643
rect 5074 609 5090 643
rect 5124 609 5140 643
rect 6706 609 6722 643
rect 6756 609 6772 643
rect 8338 609 8354 643
rect 8388 609 8404 643
rect 9970 609 9986 643
rect 10020 609 10036 643
rect 11602 609 11618 643
rect 11652 609 11668 643
rect 13234 609 13250 643
rect 13284 609 13300 643
rect 14866 609 14882 643
rect 14916 609 14932 643
rect 16498 609 16514 643
rect 16548 609 16564 643
rect 18130 609 18146 643
rect 18180 609 18196 643
rect 19762 609 19778 643
rect 19812 609 19828 643
rect 21394 609 21410 643
rect 21444 609 21460 643
rect 23026 609 23042 643
rect 23076 609 23092 643
rect 24658 609 24674 643
rect 24708 609 24724 643
rect 26290 609 26306 643
rect 26340 609 26356 643
rect 27922 609 27938 643
rect 27972 609 27988 643
rect 29554 609 29570 643
rect 29604 609 29620 643
rect 31186 609 31202 643
rect 31236 609 31252 643
rect 32818 609 32834 643
rect 32868 609 32884 643
rect 34450 609 34466 643
rect 34500 609 34516 643
rect 36082 609 36098 643
rect 36132 609 36148 643
rect 37714 609 37730 643
rect 37764 609 37780 643
rect 39346 609 39362 643
rect 39396 609 39412 643
rect 40978 609 40994 643
rect 41028 609 41044 643
rect 42610 609 42626 643
rect 42660 609 42676 643
rect 44242 609 44258 643
rect 44292 609 44308 643
rect 45874 609 45890 643
rect 45924 609 45940 643
rect 47506 609 47522 643
rect 47556 609 47572 643
rect 49138 609 49154 643
rect 49188 609 49204 643
rect 50770 609 50786 643
rect 50820 609 50836 643
<< viali >>
rect 1622 2037 1656 2071
rect 3254 2037 3288 2071
rect 4886 2037 4920 2071
rect 6518 2037 6552 2071
rect 8150 2037 8184 2071
rect 9782 2037 9816 2071
rect 11414 2037 11448 2071
rect 13046 2037 13080 2071
rect 14678 2037 14712 2071
rect 16310 2037 16344 2071
rect 17942 2037 17976 2071
rect 19574 2037 19608 2071
rect 21206 2037 21240 2071
rect 22838 2037 22872 2071
rect 24470 2037 24504 2071
rect 26102 2037 26136 2071
rect 27734 2037 27768 2071
rect 29366 2037 29400 2071
rect 30998 2037 31032 2071
rect 32630 2037 32664 2071
rect 34262 2037 34296 2071
rect 35894 2037 35928 2071
rect 37526 2037 37560 2071
rect 39158 2037 39192 2071
rect 40790 2037 40824 2071
rect 42422 2037 42456 2071
rect 44054 2037 44088 2071
rect 45686 2037 45720 2071
rect 47318 2037 47352 2071
rect 48950 2037 48984 2071
rect 50582 2037 50616 2071
rect 52214 2037 52248 2071
rect 1418 1833 1452 1867
rect 3050 1833 3084 1867
rect 4682 1833 4716 1867
rect 6314 1833 6348 1867
rect 7946 1833 7980 1867
rect 9578 1833 9612 1867
rect 11210 1833 11244 1867
rect 12842 1833 12876 1867
rect 14474 1833 14508 1867
rect 16106 1833 16140 1867
rect 17738 1833 17772 1867
rect 19370 1833 19404 1867
rect 21002 1833 21036 1867
rect 22634 1833 22668 1867
rect 24266 1833 24300 1867
rect 25898 1833 25932 1867
rect 27530 1833 27564 1867
rect 29162 1833 29196 1867
rect 30794 1833 30828 1867
rect 32426 1833 32460 1867
rect 34058 1833 34092 1867
rect 35690 1833 35724 1867
rect 37322 1833 37356 1867
rect 38954 1833 38988 1867
rect 40586 1833 40620 1867
rect 42218 1833 42252 1867
rect 43850 1833 43884 1867
rect 45482 1833 45516 1867
rect 47114 1833 47148 1867
rect 48746 1833 48780 1867
rect 50378 1833 50412 1867
rect 52010 1833 52044 1867
rect 1214 1629 1248 1663
rect 2846 1629 2880 1663
rect 4478 1629 4512 1663
rect 6110 1629 6144 1663
rect 7742 1629 7776 1663
rect 9374 1629 9408 1663
rect 11006 1629 11040 1663
rect 12638 1629 12672 1663
rect 14270 1629 14304 1663
rect 15902 1629 15936 1663
rect 17534 1629 17568 1663
rect 19166 1629 19200 1663
rect 20798 1629 20832 1663
rect 22430 1629 22464 1663
rect 24062 1629 24096 1663
rect 25694 1629 25728 1663
rect 27326 1629 27360 1663
rect 28958 1629 28992 1663
rect 30590 1629 30624 1663
rect 32222 1629 32256 1663
rect 33854 1629 33888 1663
rect 35486 1629 35520 1663
rect 37118 1629 37152 1663
rect 38750 1629 38784 1663
rect 40382 1629 40416 1663
rect 42014 1629 42048 1663
rect 43646 1629 43680 1663
rect 45278 1629 45312 1663
rect 46910 1629 46944 1663
rect 48542 1629 48576 1663
rect 50174 1629 50208 1663
rect 51806 1629 51840 1663
rect 1010 1425 1044 1459
rect 2642 1425 2676 1459
rect 4274 1425 4308 1459
rect 5906 1425 5940 1459
rect 7538 1425 7572 1459
rect 9170 1425 9204 1459
rect 10802 1425 10836 1459
rect 12434 1425 12468 1459
rect 14066 1425 14100 1459
rect 15698 1425 15732 1459
rect 17330 1425 17364 1459
rect 18962 1425 18996 1459
rect 20594 1425 20628 1459
rect 22226 1425 22260 1459
rect 23858 1425 23892 1459
rect 25490 1425 25524 1459
rect 27122 1425 27156 1459
rect 28754 1425 28788 1459
rect 30386 1425 30420 1459
rect 32018 1425 32052 1459
rect 33650 1425 33684 1459
rect 35282 1425 35316 1459
rect 36914 1425 36948 1459
rect 38546 1425 38580 1459
rect 40178 1425 40212 1459
rect 41810 1425 41844 1459
rect 43442 1425 43476 1459
rect 45074 1425 45108 1459
rect 46706 1425 46740 1459
rect 48338 1425 48372 1459
rect 49970 1425 50004 1459
rect 51602 1425 51636 1459
rect 806 1221 840 1255
rect 2438 1221 2472 1255
rect 4070 1221 4104 1255
rect 5702 1221 5736 1255
rect 7334 1221 7368 1255
rect 8966 1221 9000 1255
rect 10598 1221 10632 1255
rect 12230 1221 12264 1255
rect 13862 1221 13896 1255
rect 15494 1221 15528 1255
rect 17126 1221 17160 1255
rect 18758 1221 18792 1255
rect 20390 1221 20424 1255
rect 22022 1221 22056 1255
rect 23654 1221 23688 1255
rect 25286 1221 25320 1255
rect 26918 1221 26952 1255
rect 28550 1221 28584 1255
rect 30182 1221 30216 1255
rect 31814 1221 31848 1255
rect 33446 1221 33480 1255
rect 35078 1221 35112 1255
rect 36710 1221 36744 1255
rect 38342 1221 38376 1255
rect 39974 1221 40008 1255
rect 41606 1221 41640 1255
rect 43238 1221 43272 1255
rect 44870 1221 44904 1255
rect 46502 1221 46536 1255
rect 48134 1221 48168 1255
rect 49766 1221 49800 1255
rect 51398 1221 51432 1255
rect 602 1017 636 1051
rect 2234 1017 2268 1051
rect 3866 1017 3900 1051
rect 5498 1017 5532 1051
rect 7130 1017 7164 1051
rect 8762 1017 8796 1051
rect 10394 1017 10428 1051
rect 12026 1017 12060 1051
rect 13658 1017 13692 1051
rect 15290 1017 15324 1051
rect 16922 1017 16956 1051
rect 18554 1017 18588 1051
rect 20186 1017 20220 1051
rect 21818 1017 21852 1051
rect 23450 1017 23484 1051
rect 25082 1017 25116 1051
rect 26714 1017 26748 1051
rect 28346 1017 28380 1051
rect 29978 1017 30012 1051
rect 31610 1017 31644 1051
rect 33242 1017 33276 1051
rect 34874 1017 34908 1051
rect 36506 1017 36540 1051
rect 38138 1017 38172 1051
rect 39770 1017 39804 1051
rect 41402 1017 41436 1051
rect 43034 1017 43068 1051
rect 44666 1017 44700 1051
rect 46298 1017 46332 1051
rect 47930 1017 47964 1051
rect 49562 1017 49596 1051
rect 51194 1017 51228 1051
rect 398 813 432 847
rect 2030 813 2064 847
rect 3662 813 3696 847
rect 5294 813 5328 847
rect 6926 813 6960 847
rect 8558 813 8592 847
rect 10190 813 10224 847
rect 11822 813 11856 847
rect 13454 813 13488 847
rect 15086 813 15120 847
rect 16718 813 16752 847
rect 18350 813 18384 847
rect 19982 813 20016 847
rect 21614 813 21648 847
rect 23246 813 23280 847
rect 24878 813 24912 847
rect 26510 813 26544 847
rect 28142 813 28176 847
rect 29774 813 29808 847
rect 31406 813 31440 847
rect 33038 813 33072 847
rect 34670 813 34704 847
rect 36302 813 36336 847
rect 37934 813 37968 847
rect 39566 813 39600 847
rect 41198 813 41232 847
rect 42830 813 42864 847
rect 44462 813 44496 847
rect 46094 813 46128 847
rect 47726 813 47760 847
rect 49358 813 49392 847
rect 50990 813 51024 847
rect 194 609 228 643
rect 1826 609 1860 643
rect 3458 609 3492 643
rect 5090 609 5124 643
rect 6722 609 6756 643
rect 8354 609 8388 643
rect 9986 609 10020 643
rect 11618 609 11652 643
rect 13250 609 13284 643
rect 14882 609 14916 643
rect 16514 609 16548 643
rect 18146 609 18180 643
rect 19778 609 19812 643
rect 21410 609 21444 643
rect 23042 609 23076 643
rect 24674 609 24708 643
rect 26306 609 26340 643
rect 27938 609 27972 643
rect 29570 609 29604 643
rect 31202 609 31236 643
rect 32834 609 32868 643
rect 34466 609 34500 643
rect 36098 609 36132 643
rect 37730 609 37764 643
rect 39362 609 39396 643
rect 40994 609 41028 643
rect 42626 609 42660 643
rect 44258 609 44292 643
rect 45890 609 45924 643
rect 47522 609 47556 643
rect 49154 609 49188 643
rect 50786 609 50820 643
<< metal1 >>
rect 80 2874 108 3026
rect 172 2968 178 3020
rect 230 2968 236 3020
rect 284 2874 312 3026
rect 376 2968 382 3020
rect 434 2968 440 3020
rect 488 2874 516 3026
rect 580 2968 586 3020
rect 638 2968 644 3020
rect 692 2874 720 3026
rect 784 2968 790 3020
rect 842 2968 848 3020
rect 896 2874 924 3026
rect 988 2968 994 3020
rect 1046 2968 1052 3020
rect 1100 2874 1128 3026
rect 1192 2968 1198 3020
rect 1250 2968 1256 3020
rect 1304 2874 1332 3026
rect 1396 2968 1402 3020
rect 1454 2968 1460 3020
rect 1508 2874 1536 3026
rect 1600 2968 1606 3020
rect 1658 2968 1664 3020
rect 1712 2874 1740 3026
rect 1804 2968 1810 3020
rect 1862 2968 1868 3020
rect 1916 2874 1944 3026
rect 2008 2968 2014 3020
rect 2066 2968 2072 3020
rect 2120 2874 2148 3026
rect 2212 2968 2218 3020
rect 2270 2968 2276 3020
rect 2324 2874 2352 3026
rect 2416 2968 2422 3020
rect 2474 2968 2480 3020
rect 2528 2874 2556 3026
rect 2620 2968 2626 3020
rect 2678 2968 2684 3020
rect 2732 2874 2760 3026
rect 2824 2968 2830 3020
rect 2882 2968 2888 3020
rect 2936 2874 2964 3026
rect 3028 2968 3034 3020
rect 3086 2968 3092 3020
rect 3140 2874 3168 3026
rect 3232 2968 3238 3020
rect 3290 2968 3296 3020
rect 3344 2874 3372 3026
rect 3436 2968 3442 3020
rect 3494 2968 3500 3020
rect 3548 2874 3576 3026
rect 3640 2968 3646 3020
rect 3698 2968 3704 3020
rect 3752 2874 3780 3026
rect 3844 2968 3850 3020
rect 3902 2968 3908 3020
rect 3956 2874 3984 3026
rect 4048 2968 4054 3020
rect 4106 2968 4112 3020
rect 4160 2874 4188 3026
rect 4252 2968 4258 3020
rect 4310 2968 4316 3020
rect 4364 2874 4392 3026
rect 4456 2968 4462 3020
rect 4514 2968 4520 3020
rect 4568 2874 4596 3026
rect 4660 2968 4666 3020
rect 4718 2968 4724 3020
rect 4772 2874 4800 3026
rect 4864 2968 4870 3020
rect 4922 2968 4928 3020
rect 4976 2874 5004 3026
rect 5068 2968 5074 3020
rect 5126 2968 5132 3020
rect 5180 2874 5208 3026
rect 5272 2968 5278 3020
rect 5330 2968 5336 3020
rect 5384 2874 5412 3026
rect 5476 2968 5482 3020
rect 5534 2968 5540 3020
rect 5588 2874 5616 3026
rect 5680 2968 5686 3020
rect 5738 2968 5744 3020
rect 5792 2874 5820 3026
rect 5884 2968 5890 3020
rect 5942 2968 5948 3020
rect 5996 2874 6024 3026
rect 6088 2968 6094 3020
rect 6146 2968 6152 3020
rect 6200 2874 6228 3026
rect 6292 2968 6298 3020
rect 6350 2968 6356 3020
rect 6404 2874 6432 3026
rect 6496 2968 6502 3020
rect 6554 2968 6560 3020
rect 6608 2874 6636 3026
rect 6700 2968 6706 3020
rect 6758 2968 6764 3020
rect 6812 2874 6840 3026
rect 6904 2968 6910 3020
rect 6962 2968 6968 3020
rect 7016 2874 7044 3026
rect 7108 2968 7114 3020
rect 7166 2968 7172 3020
rect 7220 2874 7248 3026
rect 7312 2968 7318 3020
rect 7370 2968 7376 3020
rect 7424 2874 7452 3026
rect 7516 2968 7522 3020
rect 7574 2968 7580 3020
rect 7628 2874 7656 3026
rect 7720 2968 7726 3020
rect 7778 2968 7784 3020
rect 7832 2874 7860 3026
rect 7924 2968 7930 3020
rect 7982 2968 7988 3020
rect 8036 2874 8064 3026
rect 8128 2968 8134 3020
rect 8186 2968 8192 3020
rect 8240 2874 8268 3026
rect 8332 2968 8338 3020
rect 8390 2968 8396 3020
rect 8444 2874 8472 3026
rect 8536 2968 8542 3020
rect 8594 2968 8600 3020
rect 8648 2874 8676 3026
rect 8740 2968 8746 3020
rect 8798 2968 8804 3020
rect 8852 2874 8880 3026
rect 8944 2968 8950 3020
rect 9002 2968 9008 3020
rect 9056 2874 9084 3026
rect 9148 2968 9154 3020
rect 9206 2968 9212 3020
rect 9260 2874 9288 3026
rect 9352 2968 9358 3020
rect 9410 2968 9416 3020
rect 9464 2874 9492 3026
rect 9556 2968 9562 3020
rect 9614 2968 9620 3020
rect 9668 2874 9696 3026
rect 9760 2968 9766 3020
rect 9818 2968 9824 3020
rect 9872 2874 9900 3026
rect 9964 2968 9970 3020
rect 10022 2968 10028 3020
rect 10076 2874 10104 3026
rect 10168 2968 10174 3020
rect 10226 2968 10232 3020
rect 10280 2874 10308 3026
rect 10372 2968 10378 3020
rect 10430 2968 10436 3020
rect 10484 2874 10512 3026
rect 10576 2968 10582 3020
rect 10634 2968 10640 3020
rect 10688 2874 10716 3026
rect 10780 2968 10786 3020
rect 10838 2968 10844 3020
rect 10892 2874 10920 3026
rect 10984 2968 10990 3020
rect 11042 2968 11048 3020
rect 11096 2874 11124 3026
rect 11188 2968 11194 3020
rect 11246 2968 11252 3020
rect 11300 2874 11328 3026
rect 11392 2968 11398 3020
rect 11450 2968 11456 3020
rect 11504 2874 11532 3026
rect 11596 2968 11602 3020
rect 11654 2968 11660 3020
rect 11708 2874 11736 3026
rect 11800 2968 11806 3020
rect 11858 2968 11864 3020
rect 11912 2874 11940 3026
rect 12004 2968 12010 3020
rect 12062 2968 12068 3020
rect 12116 2874 12144 3026
rect 12208 2968 12214 3020
rect 12266 2968 12272 3020
rect 12320 2874 12348 3026
rect 12412 2968 12418 3020
rect 12470 2968 12476 3020
rect 12524 2874 12552 3026
rect 12616 2968 12622 3020
rect 12674 2968 12680 3020
rect 12728 2874 12756 3026
rect 12820 2968 12826 3020
rect 12878 2968 12884 3020
rect 12932 2874 12960 3026
rect 13024 2968 13030 3020
rect 13082 2968 13088 3020
rect 13136 2874 13164 3026
rect 13228 2968 13234 3020
rect 13286 2968 13292 3020
rect 13340 2874 13368 3026
rect 13432 2968 13438 3020
rect 13490 2968 13496 3020
rect 13544 2874 13572 3026
rect 13636 2968 13642 3020
rect 13694 2968 13700 3020
rect 13748 2874 13776 3026
rect 13840 2968 13846 3020
rect 13898 2968 13904 3020
rect 13952 2874 13980 3026
rect 14044 2968 14050 3020
rect 14102 2968 14108 3020
rect 14156 2874 14184 3026
rect 14248 2968 14254 3020
rect 14306 2968 14312 3020
rect 14360 2874 14388 3026
rect 14452 2968 14458 3020
rect 14510 2968 14516 3020
rect 14564 2874 14592 3026
rect 14656 2968 14662 3020
rect 14714 2968 14720 3020
rect 14768 2874 14796 3026
rect 14860 2968 14866 3020
rect 14918 2968 14924 3020
rect 14972 2874 15000 3026
rect 15064 2968 15070 3020
rect 15122 2968 15128 3020
rect 15176 2874 15204 3026
rect 15268 2968 15274 3020
rect 15326 2968 15332 3020
rect 15380 2874 15408 3026
rect 15472 2968 15478 3020
rect 15530 2968 15536 3020
rect 15584 2874 15612 3026
rect 15676 2968 15682 3020
rect 15734 2968 15740 3020
rect 15788 2874 15816 3026
rect 15880 2968 15886 3020
rect 15938 2968 15944 3020
rect 15992 2874 16020 3026
rect 16084 2968 16090 3020
rect 16142 2968 16148 3020
rect 16196 2874 16224 3026
rect 16288 2968 16294 3020
rect 16346 2968 16352 3020
rect 16400 2874 16428 3026
rect 16492 2968 16498 3020
rect 16550 2968 16556 3020
rect 16604 2874 16632 3026
rect 16696 2968 16702 3020
rect 16754 2968 16760 3020
rect 16808 2874 16836 3026
rect 16900 2968 16906 3020
rect 16958 2968 16964 3020
rect 17012 2874 17040 3026
rect 17104 2968 17110 3020
rect 17162 2968 17168 3020
rect 17216 2874 17244 3026
rect 17308 2968 17314 3020
rect 17366 2968 17372 3020
rect 17420 2874 17448 3026
rect 17512 2968 17518 3020
rect 17570 2968 17576 3020
rect 17624 2874 17652 3026
rect 17716 2968 17722 3020
rect 17774 2968 17780 3020
rect 17828 2874 17856 3026
rect 17920 2968 17926 3020
rect 17978 2968 17984 3020
rect 18032 2874 18060 3026
rect 18124 2968 18130 3020
rect 18182 2968 18188 3020
rect 18236 2874 18264 3026
rect 18328 2968 18334 3020
rect 18386 2968 18392 3020
rect 18440 2874 18468 3026
rect 18532 2968 18538 3020
rect 18590 2968 18596 3020
rect 18644 2874 18672 3026
rect 18736 2968 18742 3020
rect 18794 2968 18800 3020
rect 18848 2874 18876 3026
rect 18940 2968 18946 3020
rect 18998 2968 19004 3020
rect 19052 2874 19080 3026
rect 19144 2968 19150 3020
rect 19202 2968 19208 3020
rect 19256 2874 19284 3026
rect 19348 2968 19354 3020
rect 19406 2968 19412 3020
rect 19460 2874 19488 3026
rect 19552 2968 19558 3020
rect 19610 2968 19616 3020
rect 19664 2874 19692 3026
rect 19756 2968 19762 3020
rect 19814 2968 19820 3020
rect 19868 2874 19896 3026
rect 19960 2968 19966 3020
rect 20018 2968 20024 3020
rect 20072 2874 20100 3026
rect 20164 2968 20170 3020
rect 20222 2968 20228 3020
rect 20276 2874 20304 3026
rect 20368 2968 20374 3020
rect 20426 2968 20432 3020
rect 20480 2874 20508 3026
rect 20572 2968 20578 3020
rect 20630 2968 20636 3020
rect 20684 2874 20712 3026
rect 20776 2968 20782 3020
rect 20834 2968 20840 3020
rect 20888 2874 20916 3026
rect 20980 2968 20986 3020
rect 21038 2968 21044 3020
rect 21092 2874 21120 3026
rect 21184 2968 21190 3020
rect 21242 2968 21248 3020
rect 21296 2874 21324 3026
rect 21388 2968 21394 3020
rect 21446 2968 21452 3020
rect 21500 2874 21528 3026
rect 21592 2968 21598 3020
rect 21650 2968 21656 3020
rect 21704 2874 21732 3026
rect 21796 2968 21802 3020
rect 21854 2968 21860 3020
rect 21908 2874 21936 3026
rect 22000 2968 22006 3020
rect 22058 2968 22064 3020
rect 22112 2874 22140 3026
rect 22204 2968 22210 3020
rect 22262 2968 22268 3020
rect 22316 2874 22344 3026
rect 22408 2968 22414 3020
rect 22466 2968 22472 3020
rect 22520 2874 22548 3026
rect 22612 2968 22618 3020
rect 22670 2968 22676 3020
rect 22724 2874 22752 3026
rect 22816 2968 22822 3020
rect 22874 2968 22880 3020
rect 22928 2874 22956 3026
rect 23020 2968 23026 3020
rect 23078 2968 23084 3020
rect 23132 2874 23160 3026
rect 23224 2968 23230 3020
rect 23282 2968 23288 3020
rect 23336 2874 23364 3026
rect 23428 2968 23434 3020
rect 23486 2968 23492 3020
rect 23540 2874 23568 3026
rect 23632 2968 23638 3020
rect 23690 2968 23696 3020
rect 23744 2874 23772 3026
rect 23836 2968 23842 3020
rect 23894 2968 23900 3020
rect 23948 2874 23976 3026
rect 24040 2968 24046 3020
rect 24098 2968 24104 3020
rect 24152 2874 24180 3026
rect 24244 2968 24250 3020
rect 24302 2968 24308 3020
rect 24356 2874 24384 3026
rect 24448 2968 24454 3020
rect 24506 2968 24512 3020
rect 24560 2874 24588 3026
rect 24652 2968 24658 3020
rect 24710 2968 24716 3020
rect 24764 2874 24792 3026
rect 24856 2968 24862 3020
rect 24914 2968 24920 3020
rect 24968 2874 24996 3026
rect 25060 2968 25066 3020
rect 25118 2968 25124 3020
rect 25172 2874 25200 3026
rect 25264 2968 25270 3020
rect 25322 2968 25328 3020
rect 25376 2874 25404 3026
rect 25468 2968 25474 3020
rect 25526 2968 25532 3020
rect 25580 2874 25608 3026
rect 25672 2968 25678 3020
rect 25730 2968 25736 3020
rect 25784 2874 25812 3026
rect 25876 2968 25882 3020
rect 25934 2968 25940 3020
rect 25988 2874 26016 3026
rect 26080 2968 26086 3020
rect 26138 2968 26144 3020
rect 26192 2874 26220 3026
rect 26284 2968 26290 3020
rect 26342 2968 26348 3020
rect 26396 2874 26424 3026
rect 26488 2968 26494 3020
rect 26546 2968 26552 3020
rect 26600 2874 26628 3026
rect 26692 2968 26698 3020
rect 26750 2968 26756 3020
rect 26804 2874 26832 3026
rect 26896 2968 26902 3020
rect 26954 2968 26960 3020
rect 27008 2874 27036 3026
rect 27100 2968 27106 3020
rect 27158 2968 27164 3020
rect 27212 2874 27240 3026
rect 27304 2968 27310 3020
rect 27362 2968 27368 3020
rect 27416 2874 27444 3026
rect 27508 2968 27514 3020
rect 27566 2968 27572 3020
rect 27620 2874 27648 3026
rect 27712 2968 27718 3020
rect 27770 2968 27776 3020
rect 27824 2874 27852 3026
rect 27916 2968 27922 3020
rect 27974 2968 27980 3020
rect 28028 2874 28056 3026
rect 28120 2968 28126 3020
rect 28178 2968 28184 3020
rect 28232 2874 28260 3026
rect 28324 2968 28330 3020
rect 28382 2968 28388 3020
rect 28436 2874 28464 3026
rect 28528 2968 28534 3020
rect 28586 2968 28592 3020
rect 28640 2874 28668 3026
rect 28732 2968 28738 3020
rect 28790 2968 28796 3020
rect 28844 2874 28872 3026
rect 28936 2968 28942 3020
rect 28994 2968 29000 3020
rect 29048 2874 29076 3026
rect 29140 2968 29146 3020
rect 29198 2968 29204 3020
rect 29252 2874 29280 3026
rect 29344 2968 29350 3020
rect 29402 2968 29408 3020
rect 29456 2874 29484 3026
rect 29548 2968 29554 3020
rect 29606 2968 29612 3020
rect 29660 2874 29688 3026
rect 29752 2968 29758 3020
rect 29810 2968 29816 3020
rect 29864 2874 29892 3026
rect 29956 2968 29962 3020
rect 30014 2968 30020 3020
rect 30068 2874 30096 3026
rect 30160 2968 30166 3020
rect 30218 2968 30224 3020
rect 30272 2874 30300 3026
rect 30364 2968 30370 3020
rect 30422 2968 30428 3020
rect 30476 2874 30504 3026
rect 30568 2968 30574 3020
rect 30626 2968 30632 3020
rect 30680 2874 30708 3026
rect 30772 2968 30778 3020
rect 30830 2968 30836 3020
rect 30884 2874 30912 3026
rect 30976 2968 30982 3020
rect 31034 2968 31040 3020
rect 31088 2874 31116 3026
rect 31180 2968 31186 3020
rect 31238 2968 31244 3020
rect 31292 2874 31320 3026
rect 31384 2968 31390 3020
rect 31442 2968 31448 3020
rect 31496 2874 31524 3026
rect 31588 2968 31594 3020
rect 31646 2968 31652 3020
rect 31700 2874 31728 3026
rect 31792 2968 31798 3020
rect 31850 2968 31856 3020
rect 31904 2874 31932 3026
rect 31996 2968 32002 3020
rect 32054 2968 32060 3020
rect 32108 2874 32136 3026
rect 32200 2968 32206 3020
rect 32258 2968 32264 3020
rect 32312 2874 32340 3026
rect 32404 2968 32410 3020
rect 32462 2968 32468 3020
rect 32516 2874 32544 3026
rect 32608 2968 32614 3020
rect 32666 2968 32672 3020
rect 32720 2874 32748 3026
rect 32812 2968 32818 3020
rect 32870 2968 32876 3020
rect 32924 2874 32952 3026
rect 33016 2968 33022 3020
rect 33074 2968 33080 3020
rect 33128 2874 33156 3026
rect 33220 2968 33226 3020
rect 33278 2968 33284 3020
rect 33332 2874 33360 3026
rect 33424 2968 33430 3020
rect 33482 2968 33488 3020
rect 33536 2874 33564 3026
rect 33628 2968 33634 3020
rect 33686 2968 33692 3020
rect 33740 2874 33768 3026
rect 33832 2968 33838 3020
rect 33890 2968 33896 3020
rect 33944 2874 33972 3026
rect 34036 2968 34042 3020
rect 34094 2968 34100 3020
rect 34148 2874 34176 3026
rect 34240 2968 34246 3020
rect 34298 2968 34304 3020
rect 34352 2874 34380 3026
rect 34444 2968 34450 3020
rect 34502 2968 34508 3020
rect 34556 2874 34584 3026
rect 34648 2968 34654 3020
rect 34706 2968 34712 3020
rect 34760 2874 34788 3026
rect 34852 2968 34858 3020
rect 34910 2968 34916 3020
rect 34964 2874 34992 3026
rect 35056 2968 35062 3020
rect 35114 2968 35120 3020
rect 35168 2874 35196 3026
rect 35260 2968 35266 3020
rect 35318 2968 35324 3020
rect 35372 2874 35400 3026
rect 35464 2968 35470 3020
rect 35522 2968 35528 3020
rect 35576 2874 35604 3026
rect 35668 2968 35674 3020
rect 35726 2968 35732 3020
rect 35780 2874 35808 3026
rect 35872 2968 35878 3020
rect 35930 2968 35936 3020
rect 35984 2874 36012 3026
rect 36076 2968 36082 3020
rect 36134 2968 36140 3020
rect 36188 2874 36216 3026
rect 36280 2968 36286 3020
rect 36338 2968 36344 3020
rect 36392 2874 36420 3026
rect 36484 2968 36490 3020
rect 36542 2968 36548 3020
rect 36596 2874 36624 3026
rect 36688 2968 36694 3020
rect 36746 2968 36752 3020
rect 36800 2874 36828 3026
rect 36892 2968 36898 3020
rect 36950 2968 36956 3020
rect 37004 2874 37032 3026
rect 37096 2968 37102 3020
rect 37154 2968 37160 3020
rect 37208 2874 37236 3026
rect 37300 2968 37306 3020
rect 37358 2968 37364 3020
rect 37412 2874 37440 3026
rect 37504 2968 37510 3020
rect 37562 2968 37568 3020
rect 37616 2874 37644 3026
rect 37708 2968 37714 3020
rect 37766 2968 37772 3020
rect 37820 2874 37848 3026
rect 37912 2968 37918 3020
rect 37970 2968 37976 3020
rect 38024 2874 38052 3026
rect 38116 2968 38122 3020
rect 38174 2968 38180 3020
rect 38228 2874 38256 3026
rect 38320 2968 38326 3020
rect 38378 2968 38384 3020
rect 38432 2874 38460 3026
rect 38524 2968 38530 3020
rect 38582 2968 38588 3020
rect 38636 2874 38664 3026
rect 38728 2968 38734 3020
rect 38786 2968 38792 3020
rect 38840 2874 38868 3026
rect 38932 2968 38938 3020
rect 38990 2968 38996 3020
rect 39044 2874 39072 3026
rect 39136 2968 39142 3020
rect 39194 2968 39200 3020
rect 39248 2874 39276 3026
rect 39340 2968 39346 3020
rect 39398 2968 39404 3020
rect 39452 2874 39480 3026
rect 39544 2968 39550 3020
rect 39602 2968 39608 3020
rect 39656 2874 39684 3026
rect 39748 2968 39754 3020
rect 39806 2968 39812 3020
rect 39860 2874 39888 3026
rect 39952 2968 39958 3020
rect 40010 2968 40016 3020
rect 40064 2874 40092 3026
rect 40156 2968 40162 3020
rect 40214 2968 40220 3020
rect 40268 2874 40296 3026
rect 40360 2968 40366 3020
rect 40418 2968 40424 3020
rect 40472 2874 40500 3026
rect 40564 2968 40570 3020
rect 40622 2968 40628 3020
rect 40676 2874 40704 3026
rect 40768 2968 40774 3020
rect 40826 2968 40832 3020
rect 40880 2874 40908 3026
rect 40972 2968 40978 3020
rect 41030 2968 41036 3020
rect 41084 2874 41112 3026
rect 41176 2968 41182 3020
rect 41234 2968 41240 3020
rect 41288 2874 41316 3026
rect 41380 2968 41386 3020
rect 41438 2968 41444 3020
rect 41492 2874 41520 3026
rect 41584 2968 41590 3020
rect 41642 2968 41648 3020
rect 41696 2874 41724 3026
rect 41788 2968 41794 3020
rect 41846 2968 41852 3020
rect 41900 2874 41928 3026
rect 41992 2968 41998 3020
rect 42050 2968 42056 3020
rect 42104 2874 42132 3026
rect 42196 2968 42202 3020
rect 42254 2968 42260 3020
rect 42308 2874 42336 3026
rect 42400 2968 42406 3020
rect 42458 2968 42464 3020
rect 42512 2874 42540 3026
rect 42604 2968 42610 3020
rect 42662 2968 42668 3020
rect 42716 2874 42744 3026
rect 42808 2968 42814 3020
rect 42866 2968 42872 3020
rect 42920 2874 42948 3026
rect 43012 2968 43018 3020
rect 43070 2968 43076 3020
rect 43124 2874 43152 3026
rect 43216 2968 43222 3020
rect 43274 2968 43280 3020
rect 43328 2874 43356 3026
rect 43420 2968 43426 3020
rect 43478 2968 43484 3020
rect 43532 2874 43560 3026
rect 43624 2968 43630 3020
rect 43682 2968 43688 3020
rect 43736 2874 43764 3026
rect 43828 2968 43834 3020
rect 43886 2968 43892 3020
rect 43940 2874 43968 3026
rect 44032 2968 44038 3020
rect 44090 2968 44096 3020
rect 44144 2874 44172 3026
rect 44236 2968 44242 3020
rect 44294 2968 44300 3020
rect 44348 2874 44376 3026
rect 44440 2968 44446 3020
rect 44498 2968 44504 3020
rect 44552 2874 44580 3026
rect 44644 2968 44650 3020
rect 44702 2968 44708 3020
rect 44756 2874 44784 3026
rect 44848 2968 44854 3020
rect 44906 2968 44912 3020
rect 44960 2874 44988 3026
rect 45052 2968 45058 3020
rect 45110 2968 45116 3020
rect 45164 2874 45192 3026
rect 45256 2968 45262 3020
rect 45314 2968 45320 3020
rect 45368 2874 45396 3026
rect 45460 2968 45466 3020
rect 45518 2968 45524 3020
rect 45572 2874 45600 3026
rect 45664 2968 45670 3020
rect 45722 2968 45728 3020
rect 45776 2874 45804 3026
rect 45868 2968 45874 3020
rect 45926 2968 45932 3020
rect 45980 2874 46008 3026
rect 46072 2968 46078 3020
rect 46130 2968 46136 3020
rect 46184 2874 46212 3026
rect 46276 2968 46282 3020
rect 46334 2968 46340 3020
rect 46388 2874 46416 3026
rect 46480 2968 46486 3020
rect 46538 2968 46544 3020
rect 46592 2874 46620 3026
rect 46684 2968 46690 3020
rect 46742 2968 46748 3020
rect 46796 2874 46824 3026
rect 46888 2968 46894 3020
rect 46946 2968 46952 3020
rect 47000 2874 47028 3026
rect 47092 2968 47098 3020
rect 47150 2968 47156 3020
rect 47204 2874 47232 3026
rect 47296 2968 47302 3020
rect 47354 2968 47360 3020
rect 47408 2874 47436 3026
rect 47500 2968 47506 3020
rect 47558 2968 47564 3020
rect 47612 2874 47640 3026
rect 47704 2968 47710 3020
rect 47762 2968 47768 3020
rect 47816 2874 47844 3026
rect 47908 2968 47914 3020
rect 47966 2968 47972 3020
rect 48020 2874 48048 3026
rect 48112 2968 48118 3020
rect 48170 2968 48176 3020
rect 48224 2874 48252 3026
rect 48316 2968 48322 3020
rect 48374 2968 48380 3020
rect 48428 2874 48456 3026
rect 48520 2968 48526 3020
rect 48578 2968 48584 3020
rect 48632 2874 48660 3026
rect 48724 2968 48730 3020
rect 48782 2968 48788 3020
rect 48836 2874 48864 3026
rect 48928 2968 48934 3020
rect 48986 2968 48992 3020
rect 49040 2874 49068 3026
rect 49132 2968 49138 3020
rect 49190 2968 49196 3020
rect 49244 2874 49272 3026
rect 49336 2968 49342 3020
rect 49394 2968 49400 3020
rect 49448 2874 49476 3026
rect 49540 2968 49546 3020
rect 49598 2968 49604 3020
rect 49652 2874 49680 3026
rect 49744 2968 49750 3020
rect 49802 2968 49808 3020
rect 49856 2874 49884 3026
rect 49948 2968 49954 3020
rect 50006 2968 50012 3020
rect 50060 2874 50088 3026
rect 50152 2968 50158 3020
rect 50210 2968 50216 3020
rect 50264 2874 50292 3026
rect 50356 2968 50362 3020
rect 50414 2968 50420 3020
rect 50468 2874 50496 3026
rect 50560 2968 50566 3020
rect 50618 2968 50624 3020
rect 50672 2874 50700 3026
rect 50764 2968 50770 3020
rect 50822 2968 50828 3020
rect 50876 2874 50904 3026
rect 50968 2968 50974 3020
rect 51026 2968 51032 3020
rect 51080 2874 51108 3026
rect 51172 2968 51178 3020
rect 51230 2968 51236 3020
rect 51284 2874 51312 3026
rect 51376 2968 51382 3020
rect 51434 2968 51440 3020
rect 51488 2874 51516 3026
rect 51580 2968 51586 3020
rect 51638 2968 51644 3020
rect 51692 2874 51720 3026
rect 51784 2968 51790 3020
rect 51842 2968 51848 3020
rect 51896 2874 51924 3026
rect 51988 2968 51994 3020
rect 52046 2968 52052 3020
rect 52100 2874 52128 3026
rect 52192 2968 52198 3020
rect 52250 2968 52256 3020
rect 80 434 108 2244
rect 179 600 185 652
rect 237 600 243 652
rect 284 434 312 2244
rect 383 804 389 856
rect 441 804 447 856
rect 488 434 516 2244
rect 587 1008 593 1060
rect 645 1008 651 1060
rect 692 434 720 2244
rect 791 1212 797 1264
rect 849 1212 855 1264
rect 896 434 924 2244
rect 995 1416 1001 1468
rect 1053 1416 1059 1468
rect 1100 434 1128 2244
rect 1199 1620 1205 1672
rect 1257 1620 1263 1672
rect 1304 434 1332 2244
rect 1403 1824 1409 1876
rect 1461 1824 1467 1876
rect 1508 434 1536 2244
rect 1607 2028 1613 2080
rect 1665 2028 1671 2080
rect 1712 434 1740 2244
rect 1811 600 1817 652
rect 1869 600 1875 652
rect 1916 434 1944 2244
rect 2015 804 2021 856
rect 2073 804 2079 856
rect 2120 434 2148 2244
rect 2219 1008 2225 1060
rect 2277 1008 2283 1060
rect 2324 434 2352 2244
rect 2423 1212 2429 1264
rect 2481 1212 2487 1264
rect 2528 434 2556 2244
rect 2627 1416 2633 1468
rect 2685 1416 2691 1468
rect 2732 434 2760 2244
rect 2831 1620 2837 1672
rect 2889 1620 2895 1672
rect 2936 434 2964 2244
rect 3035 1824 3041 1876
rect 3093 1824 3099 1876
rect 3140 434 3168 2244
rect 3239 2028 3245 2080
rect 3297 2028 3303 2080
rect 3344 434 3372 2244
rect 3443 600 3449 652
rect 3501 600 3507 652
rect 3548 434 3576 2244
rect 3647 804 3653 856
rect 3705 804 3711 856
rect 3752 434 3780 2244
rect 3851 1008 3857 1060
rect 3909 1008 3915 1060
rect 3956 434 3984 2244
rect 4055 1212 4061 1264
rect 4113 1212 4119 1264
rect 4160 434 4188 2244
rect 4259 1416 4265 1468
rect 4317 1416 4323 1468
rect 4364 434 4392 2244
rect 4463 1620 4469 1672
rect 4521 1620 4527 1672
rect 4568 434 4596 2244
rect 4667 1824 4673 1876
rect 4725 1824 4731 1876
rect 4772 434 4800 2244
rect 4871 2028 4877 2080
rect 4929 2028 4935 2080
rect 4976 434 5004 2244
rect 5075 600 5081 652
rect 5133 600 5139 652
rect 5180 434 5208 2244
rect 5279 804 5285 856
rect 5337 804 5343 856
rect 5384 434 5412 2244
rect 5483 1008 5489 1060
rect 5541 1008 5547 1060
rect 5588 434 5616 2244
rect 5687 1212 5693 1264
rect 5745 1212 5751 1264
rect 5792 434 5820 2244
rect 5891 1416 5897 1468
rect 5949 1416 5955 1468
rect 5996 434 6024 2244
rect 6095 1620 6101 1672
rect 6153 1620 6159 1672
rect 6200 434 6228 2244
rect 6299 1824 6305 1876
rect 6357 1824 6363 1876
rect 6404 434 6432 2244
rect 6503 2028 6509 2080
rect 6561 2028 6567 2080
rect 6608 434 6636 2244
rect 6707 600 6713 652
rect 6765 600 6771 652
rect 6812 434 6840 2244
rect 6911 804 6917 856
rect 6969 804 6975 856
rect 7016 434 7044 2244
rect 7115 1008 7121 1060
rect 7173 1008 7179 1060
rect 7220 434 7248 2244
rect 7319 1212 7325 1264
rect 7377 1212 7383 1264
rect 7424 434 7452 2244
rect 7523 1416 7529 1468
rect 7581 1416 7587 1468
rect 7628 434 7656 2244
rect 7727 1620 7733 1672
rect 7785 1620 7791 1672
rect 7832 434 7860 2244
rect 7931 1824 7937 1876
rect 7989 1824 7995 1876
rect 8036 434 8064 2244
rect 8135 2028 8141 2080
rect 8193 2028 8199 2080
rect 8240 434 8268 2244
rect 8339 600 8345 652
rect 8397 600 8403 652
rect 8444 434 8472 2244
rect 8543 804 8549 856
rect 8601 804 8607 856
rect 8648 434 8676 2244
rect 8747 1008 8753 1060
rect 8805 1008 8811 1060
rect 8852 434 8880 2244
rect 8951 1212 8957 1264
rect 9009 1212 9015 1264
rect 9056 434 9084 2244
rect 9155 1416 9161 1468
rect 9213 1416 9219 1468
rect 9260 434 9288 2244
rect 9359 1620 9365 1672
rect 9417 1620 9423 1672
rect 9464 434 9492 2244
rect 9563 1824 9569 1876
rect 9621 1824 9627 1876
rect 9668 434 9696 2244
rect 9767 2028 9773 2080
rect 9825 2028 9831 2080
rect 9872 434 9900 2244
rect 9971 600 9977 652
rect 10029 600 10035 652
rect 10076 434 10104 2244
rect 10175 804 10181 856
rect 10233 804 10239 856
rect 10280 434 10308 2244
rect 10379 1008 10385 1060
rect 10437 1008 10443 1060
rect 10484 434 10512 2244
rect 10583 1212 10589 1264
rect 10641 1212 10647 1264
rect 10688 434 10716 2244
rect 10787 1416 10793 1468
rect 10845 1416 10851 1468
rect 10892 434 10920 2244
rect 10991 1620 10997 1672
rect 11049 1620 11055 1672
rect 11096 434 11124 2244
rect 11195 1824 11201 1876
rect 11253 1824 11259 1876
rect 11300 434 11328 2244
rect 11399 2028 11405 2080
rect 11457 2028 11463 2080
rect 11504 434 11532 2244
rect 11603 600 11609 652
rect 11661 600 11667 652
rect 11708 434 11736 2244
rect 11807 804 11813 856
rect 11865 804 11871 856
rect 11912 434 11940 2244
rect 12011 1008 12017 1060
rect 12069 1008 12075 1060
rect 12116 434 12144 2244
rect 12215 1212 12221 1264
rect 12273 1212 12279 1264
rect 12320 434 12348 2244
rect 12419 1416 12425 1468
rect 12477 1416 12483 1468
rect 12524 434 12552 2244
rect 12623 1620 12629 1672
rect 12681 1620 12687 1672
rect 12728 434 12756 2244
rect 12827 1824 12833 1876
rect 12885 1824 12891 1876
rect 12932 434 12960 2244
rect 13031 2028 13037 2080
rect 13089 2028 13095 2080
rect 13136 434 13164 2244
rect 13235 600 13241 652
rect 13293 600 13299 652
rect 13340 434 13368 2244
rect 13439 804 13445 856
rect 13497 804 13503 856
rect 13544 434 13572 2244
rect 13643 1008 13649 1060
rect 13701 1008 13707 1060
rect 13748 434 13776 2244
rect 13847 1212 13853 1264
rect 13905 1212 13911 1264
rect 13952 434 13980 2244
rect 14051 1416 14057 1468
rect 14109 1416 14115 1468
rect 14156 434 14184 2244
rect 14255 1620 14261 1672
rect 14313 1620 14319 1672
rect 14360 434 14388 2244
rect 14459 1824 14465 1876
rect 14517 1824 14523 1876
rect 14564 434 14592 2244
rect 14663 2028 14669 2080
rect 14721 2028 14727 2080
rect 14768 434 14796 2244
rect 14867 600 14873 652
rect 14925 600 14931 652
rect 14972 434 15000 2244
rect 15071 804 15077 856
rect 15129 804 15135 856
rect 15176 434 15204 2244
rect 15275 1008 15281 1060
rect 15333 1008 15339 1060
rect 15380 434 15408 2244
rect 15479 1212 15485 1264
rect 15537 1212 15543 1264
rect 15584 434 15612 2244
rect 15683 1416 15689 1468
rect 15741 1416 15747 1468
rect 15788 434 15816 2244
rect 15887 1620 15893 1672
rect 15945 1620 15951 1672
rect 15992 434 16020 2244
rect 16091 1824 16097 1876
rect 16149 1824 16155 1876
rect 16196 434 16224 2244
rect 16295 2028 16301 2080
rect 16353 2028 16359 2080
rect 16400 434 16428 2244
rect 16499 600 16505 652
rect 16557 600 16563 652
rect 16604 434 16632 2244
rect 16703 804 16709 856
rect 16761 804 16767 856
rect 16808 434 16836 2244
rect 16907 1008 16913 1060
rect 16965 1008 16971 1060
rect 17012 434 17040 2244
rect 17111 1212 17117 1264
rect 17169 1212 17175 1264
rect 17216 434 17244 2244
rect 17315 1416 17321 1468
rect 17373 1416 17379 1468
rect 17420 434 17448 2244
rect 17519 1620 17525 1672
rect 17577 1620 17583 1672
rect 17624 434 17652 2244
rect 17723 1824 17729 1876
rect 17781 1824 17787 1876
rect 17828 434 17856 2244
rect 17927 2028 17933 2080
rect 17985 2028 17991 2080
rect 18032 434 18060 2244
rect 18131 600 18137 652
rect 18189 600 18195 652
rect 18236 434 18264 2244
rect 18335 804 18341 856
rect 18393 804 18399 856
rect 18440 434 18468 2244
rect 18539 1008 18545 1060
rect 18597 1008 18603 1060
rect 18644 434 18672 2244
rect 18743 1212 18749 1264
rect 18801 1212 18807 1264
rect 18848 434 18876 2244
rect 18947 1416 18953 1468
rect 19005 1416 19011 1468
rect 19052 434 19080 2244
rect 19151 1620 19157 1672
rect 19209 1620 19215 1672
rect 19256 434 19284 2244
rect 19355 1824 19361 1876
rect 19413 1824 19419 1876
rect 19460 434 19488 2244
rect 19559 2028 19565 2080
rect 19617 2028 19623 2080
rect 19664 434 19692 2244
rect 19763 600 19769 652
rect 19821 600 19827 652
rect 19868 434 19896 2244
rect 19967 804 19973 856
rect 20025 804 20031 856
rect 20072 434 20100 2244
rect 20171 1008 20177 1060
rect 20229 1008 20235 1060
rect 20276 434 20304 2244
rect 20375 1212 20381 1264
rect 20433 1212 20439 1264
rect 20480 434 20508 2244
rect 20579 1416 20585 1468
rect 20637 1416 20643 1468
rect 20684 434 20712 2244
rect 20783 1620 20789 1672
rect 20841 1620 20847 1672
rect 20888 434 20916 2244
rect 20987 1824 20993 1876
rect 21045 1824 21051 1876
rect 21092 434 21120 2244
rect 21191 2028 21197 2080
rect 21249 2028 21255 2080
rect 21296 434 21324 2244
rect 21395 600 21401 652
rect 21453 600 21459 652
rect 21500 434 21528 2244
rect 21599 804 21605 856
rect 21657 804 21663 856
rect 21704 434 21732 2244
rect 21803 1008 21809 1060
rect 21861 1008 21867 1060
rect 21908 434 21936 2244
rect 22007 1212 22013 1264
rect 22065 1212 22071 1264
rect 22112 434 22140 2244
rect 22211 1416 22217 1468
rect 22269 1416 22275 1468
rect 22316 434 22344 2244
rect 22415 1620 22421 1672
rect 22473 1620 22479 1672
rect 22520 434 22548 2244
rect 22619 1824 22625 1876
rect 22677 1824 22683 1876
rect 22724 434 22752 2244
rect 22823 2028 22829 2080
rect 22881 2028 22887 2080
rect 22928 434 22956 2244
rect 23027 600 23033 652
rect 23085 600 23091 652
rect 23132 434 23160 2244
rect 23231 804 23237 856
rect 23289 804 23295 856
rect 23336 434 23364 2244
rect 23435 1008 23441 1060
rect 23493 1008 23499 1060
rect 23540 434 23568 2244
rect 23639 1212 23645 1264
rect 23697 1212 23703 1264
rect 23744 434 23772 2244
rect 23843 1416 23849 1468
rect 23901 1416 23907 1468
rect 23948 434 23976 2244
rect 24047 1620 24053 1672
rect 24105 1620 24111 1672
rect 24152 434 24180 2244
rect 24251 1824 24257 1876
rect 24309 1824 24315 1876
rect 24356 434 24384 2244
rect 24455 2028 24461 2080
rect 24513 2028 24519 2080
rect 24560 434 24588 2244
rect 24659 600 24665 652
rect 24717 600 24723 652
rect 24764 434 24792 2244
rect 24863 804 24869 856
rect 24921 804 24927 856
rect 24968 434 24996 2244
rect 25067 1008 25073 1060
rect 25125 1008 25131 1060
rect 25172 434 25200 2244
rect 25271 1212 25277 1264
rect 25329 1212 25335 1264
rect 25376 434 25404 2244
rect 25475 1416 25481 1468
rect 25533 1416 25539 1468
rect 25580 434 25608 2244
rect 25679 1620 25685 1672
rect 25737 1620 25743 1672
rect 25784 434 25812 2244
rect 25883 1824 25889 1876
rect 25941 1824 25947 1876
rect 25988 434 26016 2244
rect 26087 2028 26093 2080
rect 26145 2028 26151 2080
rect 26192 434 26220 2244
rect 26291 600 26297 652
rect 26349 600 26355 652
rect 26396 434 26424 2244
rect 26495 804 26501 856
rect 26553 804 26559 856
rect 26600 434 26628 2244
rect 26699 1008 26705 1060
rect 26757 1008 26763 1060
rect 26804 434 26832 2244
rect 26903 1212 26909 1264
rect 26961 1212 26967 1264
rect 27008 434 27036 2244
rect 27107 1416 27113 1468
rect 27165 1416 27171 1468
rect 27212 434 27240 2244
rect 27311 1620 27317 1672
rect 27369 1620 27375 1672
rect 27416 434 27444 2244
rect 27515 1824 27521 1876
rect 27573 1824 27579 1876
rect 27620 434 27648 2244
rect 27719 2028 27725 2080
rect 27777 2028 27783 2080
rect 27824 434 27852 2244
rect 27923 600 27929 652
rect 27981 600 27987 652
rect 28028 434 28056 2244
rect 28127 804 28133 856
rect 28185 804 28191 856
rect 28232 434 28260 2244
rect 28331 1008 28337 1060
rect 28389 1008 28395 1060
rect 28436 434 28464 2244
rect 28535 1212 28541 1264
rect 28593 1212 28599 1264
rect 28640 434 28668 2244
rect 28739 1416 28745 1468
rect 28797 1416 28803 1468
rect 28844 434 28872 2244
rect 28943 1620 28949 1672
rect 29001 1620 29007 1672
rect 29048 434 29076 2244
rect 29147 1824 29153 1876
rect 29205 1824 29211 1876
rect 29252 434 29280 2244
rect 29351 2028 29357 2080
rect 29409 2028 29415 2080
rect 29456 434 29484 2244
rect 29555 600 29561 652
rect 29613 600 29619 652
rect 29660 434 29688 2244
rect 29759 804 29765 856
rect 29817 804 29823 856
rect 29864 434 29892 2244
rect 29963 1008 29969 1060
rect 30021 1008 30027 1060
rect 30068 434 30096 2244
rect 30167 1212 30173 1264
rect 30225 1212 30231 1264
rect 30272 434 30300 2244
rect 30371 1416 30377 1468
rect 30429 1416 30435 1468
rect 30476 434 30504 2244
rect 30575 1620 30581 1672
rect 30633 1620 30639 1672
rect 30680 434 30708 2244
rect 30779 1824 30785 1876
rect 30837 1824 30843 1876
rect 30884 434 30912 2244
rect 30983 2028 30989 2080
rect 31041 2028 31047 2080
rect 31088 434 31116 2244
rect 31187 600 31193 652
rect 31245 600 31251 652
rect 31292 434 31320 2244
rect 31391 804 31397 856
rect 31449 804 31455 856
rect 31496 434 31524 2244
rect 31595 1008 31601 1060
rect 31653 1008 31659 1060
rect 31700 434 31728 2244
rect 31799 1212 31805 1264
rect 31857 1212 31863 1264
rect 31904 434 31932 2244
rect 32003 1416 32009 1468
rect 32061 1416 32067 1468
rect 32108 434 32136 2244
rect 32207 1620 32213 1672
rect 32265 1620 32271 1672
rect 32312 434 32340 2244
rect 32411 1824 32417 1876
rect 32469 1824 32475 1876
rect 32516 434 32544 2244
rect 32615 2028 32621 2080
rect 32673 2028 32679 2080
rect 32720 434 32748 2244
rect 32819 600 32825 652
rect 32877 600 32883 652
rect 32924 434 32952 2244
rect 33023 804 33029 856
rect 33081 804 33087 856
rect 33128 434 33156 2244
rect 33227 1008 33233 1060
rect 33285 1008 33291 1060
rect 33332 434 33360 2244
rect 33431 1212 33437 1264
rect 33489 1212 33495 1264
rect 33536 434 33564 2244
rect 33635 1416 33641 1468
rect 33693 1416 33699 1468
rect 33740 434 33768 2244
rect 33839 1620 33845 1672
rect 33897 1620 33903 1672
rect 33944 434 33972 2244
rect 34043 1824 34049 1876
rect 34101 1824 34107 1876
rect 34148 434 34176 2244
rect 34247 2028 34253 2080
rect 34305 2028 34311 2080
rect 34352 434 34380 2244
rect 34451 600 34457 652
rect 34509 600 34515 652
rect 34556 434 34584 2244
rect 34655 804 34661 856
rect 34713 804 34719 856
rect 34760 434 34788 2244
rect 34859 1008 34865 1060
rect 34917 1008 34923 1060
rect 34964 434 34992 2244
rect 35063 1212 35069 1264
rect 35121 1212 35127 1264
rect 35168 434 35196 2244
rect 35267 1416 35273 1468
rect 35325 1416 35331 1468
rect 35372 434 35400 2244
rect 35471 1620 35477 1672
rect 35529 1620 35535 1672
rect 35576 434 35604 2244
rect 35675 1824 35681 1876
rect 35733 1824 35739 1876
rect 35780 434 35808 2244
rect 35879 2028 35885 2080
rect 35937 2028 35943 2080
rect 35984 434 36012 2244
rect 36083 600 36089 652
rect 36141 600 36147 652
rect 36188 434 36216 2244
rect 36287 804 36293 856
rect 36345 804 36351 856
rect 36392 434 36420 2244
rect 36491 1008 36497 1060
rect 36549 1008 36555 1060
rect 36596 434 36624 2244
rect 36695 1212 36701 1264
rect 36753 1212 36759 1264
rect 36800 434 36828 2244
rect 36899 1416 36905 1468
rect 36957 1416 36963 1468
rect 37004 434 37032 2244
rect 37103 1620 37109 1672
rect 37161 1620 37167 1672
rect 37208 434 37236 2244
rect 37307 1824 37313 1876
rect 37365 1824 37371 1876
rect 37412 434 37440 2244
rect 37511 2028 37517 2080
rect 37569 2028 37575 2080
rect 37616 434 37644 2244
rect 37715 600 37721 652
rect 37773 600 37779 652
rect 37820 434 37848 2244
rect 37919 804 37925 856
rect 37977 804 37983 856
rect 38024 434 38052 2244
rect 38123 1008 38129 1060
rect 38181 1008 38187 1060
rect 38228 434 38256 2244
rect 38327 1212 38333 1264
rect 38385 1212 38391 1264
rect 38432 434 38460 2244
rect 38531 1416 38537 1468
rect 38589 1416 38595 1468
rect 38636 434 38664 2244
rect 38735 1620 38741 1672
rect 38793 1620 38799 1672
rect 38840 434 38868 2244
rect 38939 1824 38945 1876
rect 38997 1824 39003 1876
rect 39044 434 39072 2244
rect 39143 2028 39149 2080
rect 39201 2028 39207 2080
rect 39248 434 39276 2244
rect 39347 600 39353 652
rect 39405 600 39411 652
rect 39452 434 39480 2244
rect 39551 804 39557 856
rect 39609 804 39615 856
rect 39656 434 39684 2244
rect 39755 1008 39761 1060
rect 39813 1008 39819 1060
rect 39860 434 39888 2244
rect 39959 1212 39965 1264
rect 40017 1212 40023 1264
rect 40064 434 40092 2244
rect 40163 1416 40169 1468
rect 40221 1416 40227 1468
rect 40268 434 40296 2244
rect 40367 1620 40373 1672
rect 40425 1620 40431 1672
rect 40472 434 40500 2244
rect 40571 1824 40577 1876
rect 40629 1824 40635 1876
rect 40676 434 40704 2244
rect 40775 2028 40781 2080
rect 40833 2028 40839 2080
rect 40880 434 40908 2244
rect 40979 600 40985 652
rect 41037 600 41043 652
rect 41084 434 41112 2244
rect 41183 804 41189 856
rect 41241 804 41247 856
rect 41288 434 41316 2244
rect 41387 1008 41393 1060
rect 41445 1008 41451 1060
rect 41492 434 41520 2244
rect 41591 1212 41597 1264
rect 41649 1212 41655 1264
rect 41696 434 41724 2244
rect 41795 1416 41801 1468
rect 41853 1416 41859 1468
rect 41900 434 41928 2244
rect 41999 1620 42005 1672
rect 42057 1620 42063 1672
rect 42104 434 42132 2244
rect 42203 1824 42209 1876
rect 42261 1824 42267 1876
rect 42308 434 42336 2244
rect 42407 2028 42413 2080
rect 42465 2028 42471 2080
rect 42512 434 42540 2244
rect 42611 600 42617 652
rect 42669 600 42675 652
rect 42716 434 42744 2244
rect 42815 804 42821 856
rect 42873 804 42879 856
rect 42920 434 42948 2244
rect 43019 1008 43025 1060
rect 43077 1008 43083 1060
rect 43124 434 43152 2244
rect 43223 1212 43229 1264
rect 43281 1212 43287 1264
rect 43328 434 43356 2244
rect 43427 1416 43433 1468
rect 43485 1416 43491 1468
rect 43532 434 43560 2244
rect 43631 1620 43637 1672
rect 43689 1620 43695 1672
rect 43736 434 43764 2244
rect 43835 1824 43841 1876
rect 43893 1824 43899 1876
rect 43940 434 43968 2244
rect 44039 2028 44045 2080
rect 44097 2028 44103 2080
rect 44144 434 44172 2244
rect 44243 600 44249 652
rect 44301 600 44307 652
rect 44348 434 44376 2244
rect 44447 804 44453 856
rect 44505 804 44511 856
rect 44552 434 44580 2244
rect 44651 1008 44657 1060
rect 44709 1008 44715 1060
rect 44756 434 44784 2244
rect 44855 1212 44861 1264
rect 44913 1212 44919 1264
rect 44960 434 44988 2244
rect 45059 1416 45065 1468
rect 45117 1416 45123 1468
rect 45164 434 45192 2244
rect 45263 1620 45269 1672
rect 45321 1620 45327 1672
rect 45368 434 45396 2244
rect 45467 1824 45473 1876
rect 45525 1824 45531 1876
rect 45572 434 45600 2244
rect 45671 2028 45677 2080
rect 45729 2028 45735 2080
rect 45776 434 45804 2244
rect 45875 600 45881 652
rect 45933 600 45939 652
rect 45980 434 46008 2244
rect 46079 804 46085 856
rect 46137 804 46143 856
rect 46184 434 46212 2244
rect 46283 1008 46289 1060
rect 46341 1008 46347 1060
rect 46388 434 46416 2244
rect 46487 1212 46493 1264
rect 46545 1212 46551 1264
rect 46592 434 46620 2244
rect 46691 1416 46697 1468
rect 46749 1416 46755 1468
rect 46796 434 46824 2244
rect 46895 1620 46901 1672
rect 46953 1620 46959 1672
rect 47000 434 47028 2244
rect 47099 1824 47105 1876
rect 47157 1824 47163 1876
rect 47204 434 47232 2244
rect 47303 2028 47309 2080
rect 47361 2028 47367 2080
rect 47408 434 47436 2244
rect 47507 600 47513 652
rect 47565 600 47571 652
rect 47612 434 47640 2244
rect 47711 804 47717 856
rect 47769 804 47775 856
rect 47816 434 47844 2244
rect 47915 1008 47921 1060
rect 47973 1008 47979 1060
rect 48020 434 48048 2244
rect 48119 1212 48125 1264
rect 48177 1212 48183 1264
rect 48224 434 48252 2244
rect 48323 1416 48329 1468
rect 48381 1416 48387 1468
rect 48428 434 48456 2244
rect 48527 1620 48533 1672
rect 48585 1620 48591 1672
rect 48632 434 48660 2244
rect 48731 1824 48737 1876
rect 48789 1824 48795 1876
rect 48836 434 48864 2244
rect 48935 2028 48941 2080
rect 48993 2028 48999 2080
rect 49040 434 49068 2244
rect 49139 600 49145 652
rect 49197 600 49203 652
rect 49244 434 49272 2244
rect 49343 804 49349 856
rect 49401 804 49407 856
rect 49448 434 49476 2244
rect 49547 1008 49553 1060
rect 49605 1008 49611 1060
rect 49652 434 49680 2244
rect 49751 1212 49757 1264
rect 49809 1212 49815 1264
rect 49856 434 49884 2244
rect 49955 1416 49961 1468
rect 50013 1416 50019 1468
rect 50060 434 50088 2244
rect 50159 1620 50165 1672
rect 50217 1620 50223 1672
rect 50264 434 50292 2244
rect 50363 1824 50369 1876
rect 50421 1824 50427 1876
rect 50468 434 50496 2244
rect 50567 2028 50573 2080
rect 50625 2028 50631 2080
rect 50672 434 50700 2244
rect 50771 600 50777 652
rect 50829 600 50835 652
rect 50876 434 50904 2244
rect 50975 804 50981 856
rect 51033 804 51039 856
rect 51080 434 51108 2244
rect 51179 1008 51185 1060
rect 51237 1008 51243 1060
rect 51284 434 51312 2244
rect 51383 1212 51389 1264
rect 51441 1212 51447 1264
rect 51488 434 51516 2244
rect 51587 1416 51593 1468
rect 51645 1416 51651 1468
rect 51692 434 51720 2244
rect 51791 1620 51797 1672
rect 51849 1620 51855 1672
rect 51896 434 51924 2244
rect 51995 1824 52001 1876
rect 52053 1824 52059 1876
rect 52100 434 52128 2244
rect 52199 2028 52205 2080
rect 52257 2028 52263 2080
rect 62 382 68 434
rect 120 382 126 434
rect 266 382 272 434
rect 324 382 330 434
rect 470 382 476 434
rect 528 382 534 434
rect 674 382 680 434
rect 732 382 738 434
rect 878 382 884 434
rect 936 382 942 434
rect 1082 382 1088 434
rect 1140 382 1146 434
rect 1286 382 1292 434
rect 1344 382 1350 434
rect 1490 382 1496 434
rect 1548 382 1554 434
rect 1694 382 1700 434
rect 1752 382 1758 434
rect 1898 382 1904 434
rect 1956 382 1962 434
rect 2102 382 2108 434
rect 2160 382 2166 434
rect 2306 382 2312 434
rect 2364 382 2370 434
rect 2510 382 2516 434
rect 2568 382 2574 434
rect 2714 382 2720 434
rect 2772 382 2778 434
rect 2918 382 2924 434
rect 2976 382 2982 434
rect 3122 382 3128 434
rect 3180 382 3186 434
rect 3326 382 3332 434
rect 3384 382 3390 434
rect 3530 382 3536 434
rect 3588 382 3594 434
rect 3734 382 3740 434
rect 3792 382 3798 434
rect 3938 382 3944 434
rect 3996 382 4002 434
rect 4142 382 4148 434
rect 4200 382 4206 434
rect 4346 382 4352 434
rect 4404 382 4410 434
rect 4550 382 4556 434
rect 4608 382 4614 434
rect 4754 382 4760 434
rect 4812 382 4818 434
rect 4958 382 4964 434
rect 5016 382 5022 434
rect 5162 382 5168 434
rect 5220 382 5226 434
rect 5366 382 5372 434
rect 5424 382 5430 434
rect 5570 382 5576 434
rect 5628 382 5634 434
rect 5774 382 5780 434
rect 5832 382 5838 434
rect 5978 382 5984 434
rect 6036 382 6042 434
rect 6182 382 6188 434
rect 6240 382 6246 434
rect 6386 382 6392 434
rect 6444 382 6450 434
rect 6590 382 6596 434
rect 6648 382 6654 434
rect 6794 382 6800 434
rect 6852 382 6858 434
rect 6998 382 7004 434
rect 7056 382 7062 434
rect 7202 382 7208 434
rect 7260 382 7266 434
rect 7406 382 7412 434
rect 7464 382 7470 434
rect 7610 382 7616 434
rect 7668 382 7674 434
rect 7814 382 7820 434
rect 7872 382 7878 434
rect 8018 382 8024 434
rect 8076 382 8082 434
rect 8222 382 8228 434
rect 8280 382 8286 434
rect 8426 382 8432 434
rect 8484 382 8490 434
rect 8630 382 8636 434
rect 8688 382 8694 434
rect 8834 382 8840 434
rect 8892 382 8898 434
rect 9038 382 9044 434
rect 9096 382 9102 434
rect 9242 382 9248 434
rect 9300 382 9306 434
rect 9446 382 9452 434
rect 9504 382 9510 434
rect 9650 382 9656 434
rect 9708 382 9714 434
rect 9854 382 9860 434
rect 9912 382 9918 434
rect 10058 382 10064 434
rect 10116 382 10122 434
rect 10262 382 10268 434
rect 10320 382 10326 434
rect 10466 382 10472 434
rect 10524 382 10530 434
rect 10670 382 10676 434
rect 10728 382 10734 434
rect 10874 382 10880 434
rect 10932 382 10938 434
rect 11078 382 11084 434
rect 11136 382 11142 434
rect 11282 382 11288 434
rect 11340 382 11346 434
rect 11486 382 11492 434
rect 11544 382 11550 434
rect 11690 382 11696 434
rect 11748 382 11754 434
rect 11894 382 11900 434
rect 11952 382 11958 434
rect 12098 382 12104 434
rect 12156 382 12162 434
rect 12302 382 12308 434
rect 12360 382 12366 434
rect 12506 382 12512 434
rect 12564 382 12570 434
rect 12710 382 12716 434
rect 12768 382 12774 434
rect 12914 382 12920 434
rect 12972 382 12978 434
rect 13118 382 13124 434
rect 13176 382 13182 434
rect 13322 382 13328 434
rect 13380 382 13386 434
rect 13526 382 13532 434
rect 13584 382 13590 434
rect 13730 382 13736 434
rect 13788 382 13794 434
rect 13934 382 13940 434
rect 13992 382 13998 434
rect 14138 382 14144 434
rect 14196 382 14202 434
rect 14342 382 14348 434
rect 14400 382 14406 434
rect 14546 382 14552 434
rect 14604 382 14610 434
rect 14750 382 14756 434
rect 14808 382 14814 434
rect 14954 382 14960 434
rect 15012 382 15018 434
rect 15158 382 15164 434
rect 15216 382 15222 434
rect 15362 382 15368 434
rect 15420 382 15426 434
rect 15566 382 15572 434
rect 15624 382 15630 434
rect 15770 382 15776 434
rect 15828 382 15834 434
rect 15974 382 15980 434
rect 16032 382 16038 434
rect 16178 382 16184 434
rect 16236 382 16242 434
rect 16382 382 16388 434
rect 16440 382 16446 434
rect 16586 382 16592 434
rect 16644 382 16650 434
rect 16790 382 16796 434
rect 16848 382 16854 434
rect 16994 382 17000 434
rect 17052 382 17058 434
rect 17198 382 17204 434
rect 17256 382 17262 434
rect 17402 382 17408 434
rect 17460 382 17466 434
rect 17606 382 17612 434
rect 17664 382 17670 434
rect 17810 382 17816 434
rect 17868 382 17874 434
rect 18014 382 18020 434
rect 18072 382 18078 434
rect 18218 382 18224 434
rect 18276 382 18282 434
rect 18422 382 18428 434
rect 18480 382 18486 434
rect 18626 382 18632 434
rect 18684 382 18690 434
rect 18830 382 18836 434
rect 18888 382 18894 434
rect 19034 382 19040 434
rect 19092 382 19098 434
rect 19238 382 19244 434
rect 19296 382 19302 434
rect 19442 382 19448 434
rect 19500 382 19506 434
rect 19646 382 19652 434
rect 19704 382 19710 434
rect 19850 382 19856 434
rect 19908 382 19914 434
rect 20054 382 20060 434
rect 20112 382 20118 434
rect 20258 382 20264 434
rect 20316 382 20322 434
rect 20462 382 20468 434
rect 20520 382 20526 434
rect 20666 382 20672 434
rect 20724 382 20730 434
rect 20870 382 20876 434
rect 20928 382 20934 434
rect 21074 382 21080 434
rect 21132 382 21138 434
rect 21278 382 21284 434
rect 21336 382 21342 434
rect 21482 382 21488 434
rect 21540 382 21546 434
rect 21686 382 21692 434
rect 21744 382 21750 434
rect 21890 382 21896 434
rect 21948 382 21954 434
rect 22094 382 22100 434
rect 22152 382 22158 434
rect 22298 382 22304 434
rect 22356 382 22362 434
rect 22502 382 22508 434
rect 22560 382 22566 434
rect 22706 382 22712 434
rect 22764 382 22770 434
rect 22910 382 22916 434
rect 22968 382 22974 434
rect 23114 382 23120 434
rect 23172 382 23178 434
rect 23318 382 23324 434
rect 23376 382 23382 434
rect 23522 382 23528 434
rect 23580 382 23586 434
rect 23726 382 23732 434
rect 23784 382 23790 434
rect 23930 382 23936 434
rect 23988 382 23994 434
rect 24134 382 24140 434
rect 24192 382 24198 434
rect 24338 382 24344 434
rect 24396 382 24402 434
rect 24542 382 24548 434
rect 24600 382 24606 434
rect 24746 382 24752 434
rect 24804 382 24810 434
rect 24950 382 24956 434
rect 25008 382 25014 434
rect 25154 382 25160 434
rect 25212 382 25218 434
rect 25358 382 25364 434
rect 25416 382 25422 434
rect 25562 382 25568 434
rect 25620 382 25626 434
rect 25766 382 25772 434
rect 25824 382 25830 434
rect 25970 382 25976 434
rect 26028 382 26034 434
rect 26174 382 26180 434
rect 26232 382 26238 434
rect 26378 382 26384 434
rect 26436 382 26442 434
rect 26582 382 26588 434
rect 26640 382 26646 434
rect 26786 382 26792 434
rect 26844 382 26850 434
rect 26990 382 26996 434
rect 27048 382 27054 434
rect 27194 382 27200 434
rect 27252 382 27258 434
rect 27398 382 27404 434
rect 27456 382 27462 434
rect 27602 382 27608 434
rect 27660 382 27666 434
rect 27806 382 27812 434
rect 27864 382 27870 434
rect 28010 382 28016 434
rect 28068 382 28074 434
rect 28214 382 28220 434
rect 28272 382 28278 434
rect 28418 382 28424 434
rect 28476 382 28482 434
rect 28622 382 28628 434
rect 28680 382 28686 434
rect 28826 382 28832 434
rect 28884 382 28890 434
rect 29030 382 29036 434
rect 29088 382 29094 434
rect 29234 382 29240 434
rect 29292 382 29298 434
rect 29438 382 29444 434
rect 29496 382 29502 434
rect 29642 382 29648 434
rect 29700 382 29706 434
rect 29846 382 29852 434
rect 29904 382 29910 434
rect 30050 382 30056 434
rect 30108 382 30114 434
rect 30254 382 30260 434
rect 30312 382 30318 434
rect 30458 382 30464 434
rect 30516 382 30522 434
rect 30662 382 30668 434
rect 30720 382 30726 434
rect 30866 382 30872 434
rect 30924 382 30930 434
rect 31070 382 31076 434
rect 31128 382 31134 434
rect 31274 382 31280 434
rect 31332 382 31338 434
rect 31478 382 31484 434
rect 31536 382 31542 434
rect 31682 382 31688 434
rect 31740 382 31746 434
rect 31886 382 31892 434
rect 31944 382 31950 434
rect 32090 382 32096 434
rect 32148 382 32154 434
rect 32294 382 32300 434
rect 32352 382 32358 434
rect 32498 382 32504 434
rect 32556 382 32562 434
rect 32702 382 32708 434
rect 32760 382 32766 434
rect 32906 382 32912 434
rect 32964 382 32970 434
rect 33110 382 33116 434
rect 33168 382 33174 434
rect 33314 382 33320 434
rect 33372 382 33378 434
rect 33518 382 33524 434
rect 33576 382 33582 434
rect 33722 382 33728 434
rect 33780 382 33786 434
rect 33926 382 33932 434
rect 33984 382 33990 434
rect 34130 382 34136 434
rect 34188 382 34194 434
rect 34334 382 34340 434
rect 34392 382 34398 434
rect 34538 382 34544 434
rect 34596 382 34602 434
rect 34742 382 34748 434
rect 34800 382 34806 434
rect 34946 382 34952 434
rect 35004 382 35010 434
rect 35150 382 35156 434
rect 35208 382 35214 434
rect 35354 382 35360 434
rect 35412 382 35418 434
rect 35558 382 35564 434
rect 35616 382 35622 434
rect 35762 382 35768 434
rect 35820 382 35826 434
rect 35966 382 35972 434
rect 36024 382 36030 434
rect 36170 382 36176 434
rect 36228 382 36234 434
rect 36374 382 36380 434
rect 36432 382 36438 434
rect 36578 382 36584 434
rect 36636 382 36642 434
rect 36782 382 36788 434
rect 36840 382 36846 434
rect 36986 382 36992 434
rect 37044 382 37050 434
rect 37190 382 37196 434
rect 37248 382 37254 434
rect 37394 382 37400 434
rect 37452 382 37458 434
rect 37598 382 37604 434
rect 37656 382 37662 434
rect 37802 382 37808 434
rect 37860 382 37866 434
rect 38006 382 38012 434
rect 38064 382 38070 434
rect 38210 382 38216 434
rect 38268 382 38274 434
rect 38414 382 38420 434
rect 38472 382 38478 434
rect 38618 382 38624 434
rect 38676 382 38682 434
rect 38822 382 38828 434
rect 38880 382 38886 434
rect 39026 382 39032 434
rect 39084 382 39090 434
rect 39230 382 39236 434
rect 39288 382 39294 434
rect 39434 382 39440 434
rect 39492 382 39498 434
rect 39638 382 39644 434
rect 39696 382 39702 434
rect 39842 382 39848 434
rect 39900 382 39906 434
rect 40046 382 40052 434
rect 40104 382 40110 434
rect 40250 382 40256 434
rect 40308 382 40314 434
rect 40454 382 40460 434
rect 40512 382 40518 434
rect 40658 382 40664 434
rect 40716 382 40722 434
rect 40862 382 40868 434
rect 40920 382 40926 434
rect 41066 382 41072 434
rect 41124 382 41130 434
rect 41270 382 41276 434
rect 41328 382 41334 434
rect 41474 382 41480 434
rect 41532 382 41538 434
rect 41678 382 41684 434
rect 41736 382 41742 434
rect 41882 382 41888 434
rect 41940 382 41946 434
rect 42086 382 42092 434
rect 42144 382 42150 434
rect 42290 382 42296 434
rect 42348 382 42354 434
rect 42494 382 42500 434
rect 42552 382 42558 434
rect 42698 382 42704 434
rect 42756 382 42762 434
rect 42902 382 42908 434
rect 42960 382 42966 434
rect 43106 382 43112 434
rect 43164 382 43170 434
rect 43310 382 43316 434
rect 43368 382 43374 434
rect 43514 382 43520 434
rect 43572 382 43578 434
rect 43718 382 43724 434
rect 43776 382 43782 434
rect 43922 382 43928 434
rect 43980 382 43986 434
rect 44126 382 44132 434
rect 44184 382 44190 434
rect 44330 382 44336 434
rect 44388 382 44394 434
rect 44534 382 44540 434
rect 44592 382 44598 434
rect 44738 382 44744 434
rect 44796 382 44802 434
rect 44942 382 44948 434
rect 45000 382 45006 434
rect 45146 382 45152 434
rect 45204 382 45210 434
rect 45350 382 45356 434
rect 45408 382 45414 434
rect 45554 382 45560 434
rect 45612 382 45618 434
rect 45758 382 45764 434
rect 45816 382 45822 434
rect 45962 382 45968 434
rect 46020 382 46026 434
rect 46166 382 46172 434
rect 46224 382 46230 434
rect 46370 382 46376 434
rect 46428 382 46434 434
rect 46574 382 46580 434
rect 46632 382 46638 434
rect 46778 382 46784 434
rect 46836 382 46842 434
rect 46982 382 46988 434
rect 47040 382 47046 434
rect 47186 382 47192 434
rect 47244 382 47250 434
rect 47390 382 47396 434
rect 47448 382 47454 434
rect 47594 382 47600 434
rect 47652 382 47658 434
rect 47798 382 47804 434
rect 47856 382 47862 434
rect 48002 382 48008 434
rect 48060 382 48066 434
rect 48206 382 48212 434
rect 48264 382 48270 434
rect 48410 382 48416 434
rect 48468 382 48474 434
rect 48614 382 48620 434
rect 48672 382 48678 434
rect 48818 382 48824 434
rect 48876 382 48882 434
rect 49022 382 49028 434
rect 49080 382 49086 434
rect 49226 382 49232 434
rect 49284 382 49290 434
rect 49430 382 49436 434
rect 49488 382 49494 434
rect 49634 382 49640 434
rect 49692 382 49698 434
rect 49838 382 49844 434
rect 49896 382 49902 434
rect 50042 382 50048 434
rect 50100 382 50106 434
rect 50246 382 50252 434
rect 50304 382 50310 434
rect 50450 382 50456 434
rect 50508 382 50514 434
rect 50654 382 50660 434
rect 50712 382 50718 434
rect 50858 382 50864 434
rect 50916 382 50922 434
rect 51062 382 51068 434
rect 51120 382 51126 434
rect 51266 382 51272 434
rect 51324 382 51330 434
rect 51470 382 51476 434
rect 51528 382 51534 434
rect 51674 382 51680 434
rect 51732 382 51738 434
rect 51878 382 51884 434
rect 51936 382 51942 434
rect 52082 382 52088 434
rect 52140 382 52146 434
<< via1 >>
rect 178 2968 230 3020
rect 382 2968 434 3020
rect 586 2968 638 3020
rect 790 2968 842 3020
rect 994 2968 1046 3020
rect 1198 2968 1250 3020
rect 1402 2968 1454 3020
rect 1606 2968 1658 3020
rect 1810 2968 1862 3020
rect 2014 2968 2066 3020
rect 2218 2968 2270 3020
rect 2422 2968 2474 3020
rect 2626 2968 2678 3020
rect 2830 2968 2882 3020
rect 3034 2968 3086 3020
rect 3238 2968 3290 3020
rect 3442 2968 3494 3020
rect 3646 2968 3698 3020
rect 3850 2968 3902 3020
rect 4054 2968 4106 3020
rect 4258 2968 4310 3020
rect 4462 2968 4514 3020
rect 4666 2968 4718 3020
rect 4870 2968 4922 3020
rect 5074 2968 5126 3020
rect 5278 2968 5330 3020
rect 5482 2968 5534 3020
rect 5686 2968 5738 3020
rect 5890 2968 5942 3020
rect 6094 2968 6146 3020
rect 6298 2968 6350 3020
rect 6502 2968 6554 3020
rect 6706 2968 6758 3020
rect 6910 2968 6962 3020
rect 7114 2968 7166 3020
rect 7318 2968 7370 3020
rect 7522 2968 7574 3020
rect 7726 2968 7778 3020
rect 7930 2968 7982 3020
rect 8134 2968 8186 3020
rect 8338 2968 8390 3020
rect 8542 2968 8594 3020
rect 8746 2968 8798 3020
rect 8950 2968 9002 3020
rect 9154 2968 9206 3020
rect 9358 2968 9410 3020
rect 9562 2968 9614 3020
rect 9766 2968 9818 3020
rect 9970 2968 10022 3020
rect 10174 2968 10226 3020
rect 10378 2968 10430 3020
rect 10582 2968 10634 3020
rect 10786 2968 10838 3020
rect 10990 2968 11042 3020
rect 11194 2968 11246 3020
rect 11398 2968 11450 3020
rect 11602 2968 11654 3020
rect 11806 2968 11858 3020
rect 12010 2968 12062 3020
rect 12214 2968 12266 3020
rect 12418 2968 12470 3020
rect 12622 2968 12674 3020
rect 12826 2968 12878 3020
rect 13030 2968 13082 3020
rect 13234 2968 13286 3020
rect 13438 2968 13490 3020
rect 13642 2968 13694 3020
rect 13846 2968 13898 3020
rect 14050 2968 14102 3020
rect 14254 2968 14306 3020
rect 14458 2968 14510 3020
rect 14662 2968 14714 3020
rect 14866 2968 14918 3020
rect 15070 2968 15122 3020
rect 15274 2968 15326 3020
rect 15478 2968 15530 3020
rect 15682 2968 15734 3020
rect 15886 2968 15938 3020
rect 16090 2968 16142 3020
rect 16294 2968 16346 3020
rect 16498 2968 16550 3020
rect 16702 2968 16754 3020
rect 16906 2968 16958 3020
rect 17110 2968 17162 3020
rect 17314 2968 17366 3020
rect 17518 2968 17570 3020
rect 17722 2968 17774 3020
rect 17926 2968 17978 3020
rect 18130 2968 18182 3020
rect 18334 2968 18386 3020
rect 18538 2968 18590 3020
rect 18742 2968 18794 3020
rect 18946 2968 18998 3020
rect 19150 2968 19202 3020
rect 19354 2968 19406 3020
rect 19558 2968 19610 3020
rect 19762 2968 19814 3020
rect 19966 2968 20018 3020
rect 20170 2968 20222 3020
rect 20374 2968 20426 3020
rect 20578 2968 20630 3020
rect 20782 2968 20834 3020
rect 20986 2968 21038 3020
rect 21190 2968 21242 3020
rect 21394 2968 21446 3020
rect 21598 2968 21650 3020
rect 21802 2968 21854 3020
rect 22006 2968 22058 3020
rect 22210 2968 22262 3020
rect 22414 2968 22466 3020
rect 22618 2968 22670 3020
rect 22822 2968 22874 3020
rect 23026 2968 23078 3020
rect 23230 2968 23282 3020
rect 23434 2968 23486 3020
rect 23638 2968 23690 3020
rect 23842 2968 23894 3020
rect 24046 2968 24098 3020
rect 24250 2968 24302 3020
rect 24454 2968 24506 3020
rect 24658 2968 24710 3020
rect 24862 2968 24914 3020
rect 25066 2968 25118 3020
rect 25270 2968 25322 3020
rect 25474 2968 25526 3020
rect 25678 2968 25730 3020
rect 25882 2968 25934 3020
rect 26086 2968 26138 3020
rect 26290 2968 26342 3020
rect 26494 2968 26546 3020
rect 26698 2968 26750 3020
rect 26902 2968 26954 3020
rect 27106 2968 27158 3020
rect 27310 2968 27362 3020
rect 27514 2968 27566 3020
rect 27718 2968 27770 3020
rect 27922 2968 27974 3020
rect 28126 2968 28178 3020
rect 28330 2968 28382 3020
rect 28534 2968 28586 3020
rect 28738 2968 28790 3020
rect 28942 2968 28994 3020
rect 29146 2968 29198 3020
rect 29350 2968 29402 3020
rect 29554 2968 29606 3020
rect 29758 2968 29810 3020
rect 29962 2968 30014 3020
rect 30166 2968 30218 3020
rect 30370 2968 30422 3020
rect 30574 2968 30626 3020
rect 30778 2968 30830 3020
rect 30982 2968 31034 3020
rect 31186 2968 31238 3020
rect 31390 2968 31442 3020
rect 31594 2968 31646 3020
rect 31798 2968 31850 3020
rect 32002 2968 32054 3020
rect 32206 2968 32258 3020
rect 32410 2968 32462 3020
rect 32614 2968 32666 3020
rect 32818 2968 32870 3020
rect 33022 2968 33074 3020
rect 33226 2968 33278 3020
rect 33430 2968 33482 3020
rect 33634 2968 33686 3020
rect 33838 2968 33890 3020
rect 34042 2968 34094 3020
rect 34246 2968 34298 3020
rect 34450 2968 34502 3020
rect 34654 2968 34706 3020
rect 34858 2968 34910 3020
rect 35062 2968 35114 3020
rect 35266 2968 35318 3020
rect 35470 2968 35522 3020
rect 35674 2968 35726 3020
rect 35878 2968 35930 3020
rect 36082 2968 36134 3020
rect 36286 2968 36338 3020
rect 36490 2968 36542 3020
rect 36694 2968 36746 3020
rect 36898 2968 36950 3020
rect 37102 2968 37154 3020
rect 37306 2968 37358 3020
rect 37510 2968 37562 3020
rect 37714 2968 37766 3020
rect 37918 2968 37970 3020
rect 38122 2968 38174 3020
rect 38326 2968 38378 3020
rect 38530 2968 38582 3020
rect 38734 2968 38786 3020
rect 38938 2968 38990 3020
rect 39142 2968 39194 3020
rect 39346 2968 39398 3020
rect 39550 2968 39602 3020
rect 39754 2968 39806 3020
rect 39958 2968 40010 3020
rect 40162 2968 40214 3020
rect 40366 2968 40418 3020
rect 40570 2968 40622 3020
rect 40774 2968 40826 3020
rect 40978 2968 41030 3020
rect 41182 2968 41234 3020
rect 41386 2968 41438 3020
rect 41590 2968 41642 3020
rect 41794 2968 41846 3020
rect 41998 2968 42050 3020
rect 42202 2968 42254 3020
rect 42406 2968 42458 3020
rect 42610 2968 42662 3020
rect 42814 2968 42866 3020
rect 43018 2968 43070 3020
rect 43222 2968 43274 3020
rect 43426 2968 43478 3020
rect 43630 2968 43682 3020
rect 43834 2968 43886 3020
rect 44038 2968 44090 3020
rect 44242 2968 44294 3020
rect 44446 2968 44498 3020
rect 44650 2968 44702 3020
rect 44854 2968 44906 3020
rect 45058 2968 45110 3020
rect 45262 2968 45314 3020
rect 45466 2968 45518 3020
rect 45670 2968 45722 3020
rect 45874 2968 45926 3020
rect 46078 2968 46130 3020
rect 46282 2968 46334 3020
rect 46486 2968 46538 3020
rect 46690 2968 46742 3020
rect 46894 2968 46946 3020
rect 47098 2968 47150 3020
rect 47302 2968 47354 3020
rect 47506 2968 47558 3020
rect 47710 2968 47762 3020
rect 47914 2968 47966 3020
rect 48118 2968 48170 3020
rect 48322 2968 48374 3020
rect 48526 2968 48578 3020
rect 48730 2968 48782 3020
rect 48934 2968 48986 3020
rect 49138 2968 49190 3020
rect 49342 2968 49394 3020
rect 49546 2968 49598 3020
rect 49750 2968 49802 3020
rect 49954 2968 50006 3020
rect 50158 2968 50210 3020
rect 50362 2968 50414 3020
rect 50566 2968 50618 3020
rect 50770 2968 50822 3020
rect 50974 2968 51026 3020
rect 51178 2968 51230 3020
rect 51382 2968 51434 3020
rect 51586 2968 51638 3020
rect 51790 2968 51842 3020
rect 51994 2968 52046 3020
rect 52198 2968 52250 3020
rect 185 643 237 652
rect 185 609 194 643
rect 194 609 228 643
rect 228 609 237 643
rect 185 600 237 609
rect 389 847 441 856
rect 389 813 398 847
rect 398 813 432 847
rect 432 813 441 847
rect 389 804 441 813
rect 593 1051 645 1060
rect 593 1017 602 1051
rect 602 1017 636 1051
rect 636 1017 645 1051
rect 593 1008 645 1017
rect 797 1255 849 1264
rect 797 1221 806 1255
rect 806 1221 840 1255
rect 840 1221 849 1255
rect 797 1212 849 1221
rect 1001 1459 1053 1468
rect 1001 1425 1010 1459
rect 1010 1425 1044 1459
rect 1044 1425 1053 1459
rect 1001 1416 1053 1425
rect 1205 1663 1257 1672
rect 1205 1629 1214 1663
rect 1214 1629 1248 1663
rect 1248 1629 1257 1663
rect 1205 1620 1257 1629
rect 1409 1867 1461 1876
rect 1409 1833 1418 1867
rect 1418 1833 1452 1867
rect 1452 1833 1461 1867
rect 1409 1824 1461 1833
rect 1613 2071 1665 2080
rect 1613 2037 1622 2071
rect 1622 2037 1656 2071
rect 1656 2037 1665 2071
rect 1613 2028 1665 2037
rect 1817 643 1869 652
rect 1817 609 1826 643
rect 1826 609 1860 643
rect 1860 609 1869 643
rect 1817 600 1869 609
rect 2021 847 2073 856
rect 2021 813 2030 847
rect 2030 813 2064 847
rect 2064 813 2073 847
rect 2021 804 2073 813
rect 2225 1051 2277 1060
rect 2225 1017 2234 1051
rect 2234 1017 2268 1051
rect 2268 1017 2277 1051
rect 2225 1008 2277 1017
rect 2429 1255 2481 1264
rect 2429 1221 2438 1255
rect 2438 1221 2472 1255
rect 2472 1221 2481 1255
rect 2429 1212 2481 1221
rect 2633 1459 2685 1468
rect 2633 1425 2642 1459
rect 2642 1425 2676 1459
rect 2676 1425 2685 1459
rect 2633 1416 2685 1425
rect 2837 1663 2889 1672
rect 2837 1629 2846 1663
rect 2846 1629 2880 1663
rect 2880 1629 2889 1663
rect 2837 1620 2889 1629
rect 3041 1867 3093 1876
rect 3041 1833 3050 1867
rect 3050 1833 3084 1867
rect 3084 1833 3093 1867
rect 3041 1824 3093 1833
rect 3245 2071 3297 2080
rect 3245 2037 3254 2071
rect 3254 2037 3288 2071
rect 3288 2037 3297 2071
rect 3245 2028 3297 2037
rect 3449 643 3501 652
rect 3449 609 3458 643
rect 3458 609 3492 643
rect 3492 609 3501 643
rect 3449 600 3501 609
rect 3653 847 3705 856
rect 3653 813 3662 847
rect 3662 813 3696 847
rect 3696 813 3705 847
rect 3653 804 3705 813
rect 3857 1051 3909 1060
rect 3857 1017 3866 1051
rect 3866 1017 3900 1051
rect 3900 1017 3909 1051
rect 3857 1008 3909 1017
rect 4061 1255 4113 1264
rect 4061 1221 4070 1255
rect 4070 1221 4104 1255
rect 4104 1221 4113 1255
rect 4061 1212 4113 1221
rect 4265 1459 4317 1468
rect 4265 1425 4274 1459
rect 4274 1425 4308 1459
rect 4308 1425 4317 1459
rect 4265 1416 4317 1425
rect 4469 1663 4521 1672
rect 4469 1629 4478 1663
rect 4478 1629 4512 1663
rect 4512 1629 4521 1663
rect 4469 1620 4521 1629
rect 4673 1867 4725 1876
rect 4673 1833 4682 1867
rect 4682 1833 4716 1867
rect 4716 1833 4725 1867
rect 4673 1824 4725 1833
rect 4877 2071 4929 2080
rect 4877 2037 4886 2071
rect 4886 2037 4920 2071
rect 4920 2037 4929 2071
rect 4877 2028 4929 2037
rect 5081 643 5133 652
rect 5081 609 5090 643
rect 5090 609 5124 643
rect 5124 609 5133 643
rect 5081 600 5133 609
rect 5285 847 5337 856
rect 5285 813 5294 847
rect 5294 813 5328 847
rect 5328 813 5337 847
rect 5285 804 5337 813
rect 5489 1051 5541 1060
rect 5489 1017 5498 1051
rect 5498 1017 5532 1051
rect 5532 1017 5541 1051
rect 5489 1008 5541 1017
rect 5693 1255 5745 1264
rect 5693 1221 5702 1255
rect 5702 1221 5736 1255
rect 5736 1221 5745 1255
rect 5693 1212 5745 1221
rect 5897 1459 5949 1468
rect 5897 1425 5906 1459
rect 5906 1425 5940 1459
rect 5940 1425 5949 1459
rect 5897 1416 5949 1425
rect 6101 1663 6153 1672
rect 6101 1629 6110 1663
rect 6110 1629 6144 1663
rect 6144 1629 6153 1663
rect 6101 1620 6153 1629
rect 6305 1867 6357 1876
rect 6305 1833 6314 1867
rect 6314 1833 6348 1867
rect 6348 1833 6357 1867
rect 6305 1824 6357 1833
rect 6509 2071 6561 2080
rect 6509 2037 6518 2071
rect 6518 2037 6552 2071
rect 6552 2037 6561 2071
rect 6509 2028 6561 2037
rect 6713 643 6765 652
rect 6713 609 6722 643
rect 6722 609 6756 643
rect 6756 609 6765 643
rect 6713 600 6765 609
rect 6917 847 6969 856
rect 6917 813 6926 847
rect 6926 813 6960 847
rect 6960 813 6969 847
rect 6917 804 6969 813
rect 7121 1051 7173 1060
rect 7121 1017 7130 1051
rect 7130 1017 7164 1051
rect 7164 1017 7173 1051
rect 7121 1008 7173 1017
rect 7325 1255 7377 1264
rect 7325 1221 7334 1255
rect 7334 1221 7368 1255
rect 7368 1221 7377 1255
rect 7325 1212 7377 1221
rect 7529 1459 7581 1468
rect 7529 1425 7538 1459
rect 7538 1425 7572 1459
rect 7572 1425 7581 1459
rect 7529 1416 7581 1425
rect 7733 1663 7785 1672
rect 7733 1629 7742 1663
rect 7742 1629 7776 1663
rect 7776 1629 7785 1663
rect 7733 1620 7785 1629
rect 7937 1867 7989 1876
rect 7937 1833 7946 1867
rect 7946 1833 7980 1867
rect 7980 1833 7989 1867
rect 7937 1824 7989 1833
rect 8141 2071 8193 2080
rect 8141 2037 8150 2071
rect 8150 2037 8184 2071
rect 8184 2037 8193 2071
rect 8141 2028 8193 2037
rect 8345 643 8397 652
rect 8345 609 8354 643
rect 8354 609 8388 643
rect 8388 609 8397 643
rect 8345 600 8397 609
rect 8549 847 8601 856
rect 8549 813 8558 847
rect 8558 813 8592 847
rect 8592 813 8601 847
rect 8549 804 8601 813
rect 8753 1051 8805 1060
rect 8753 1017 8762 1051
rect 8762 1017 8796 1051
rect 8796 1017 8805 1051
rect 8753 1008 8805 1017
rect 8957 1255 9009 1264
rect 8957 1221 8966 1255
rect 8966 1221 9000 1255
rect 9000 1221 9009 1255
rect 8957 1212 9009 1221
rect 9161 1459 9213 1468
rect 9161 1425 9170 1459
rect 9170 1425 9204 1459
rect 9204 1425 9213 1459
rect 9161 1416 9213 1425
rect 9365 1663 9417 1672
rect 9365 1629 9374 1663
rect 9374 1629 9408 1663
rect 9408 1629 9417 1663
rect 9365 1620 9417 1629
rect 9569 1867 9621 1876
rect 9569 1833 9578 1867
rect 9578 1833 9612 1867
rect 9612 1833 9621 1867
rect 9569 1824 9621 1833
rect 9773 2071 9825 2080
rect 9773 2037 9782 2071
rect 9782 2037 9816 2071
rect 9816 2037 9825 2071
rect 9773 2028 9825 2037
rect 9977 643 10029 652
rect 9977 609 9986 643
rect 9986 609 10020 643
rect 10020 609 10029 643
rect 9977 600 10029 609
rect 10181 847 10233 856
rect 10181 813 10190 847
rect 10190 813 10224 847
rect 10224 813 10233 847
rect 10181 804 10233 813
rect 10385 1051 10437 1060
rect 10385 1017 10394 1051
rect 10394 1017 10428 1051
rect 10428 1017 10437 1051
rect 10385 1008 10437 1017
rect 10589 1255 10641 1264
rect 10589 1221 10598 1255
rect 10598 1221 10632 1255
rect 10632 1221 10641 1255
rect 10589 1212 10641 1221
rect 10793 1459 10845 1468
rect 10793 1425 10802 1459
rect 10802 1425 10836 1459
rect 10836 1425 10845 1459
rect 10793 1416 10845 1425
rect 10997 1663 11049 1672
rect 10997 1629 11006 1663
rect 11006 1629 11040 1663
rect 11040 1629 11049 1663
rect 10997 1620 11049 1629
rect 11201 1867 11253 1876
rect 11201 1833 11210 1867
rect 11210 1833 11244 1867
rect 11244 1833 11253 1867
rect 11201 1824 11253 1833
rect 11405 2071 11457 2080
rect 11405 2037 11414 2071
rect 11414 2037 11448 2071
rect 11448 2037 11457 2071
rect 11405 2028 11457 2037
rect 11609 643 11661 652
rect 11609 609 11618 643
rect 11618 609 11652 643
rect 11652 609 11661 643
rect 11609 600 11661 609
rect 11813 847 11865 856
rect 11813 813 11822 847
rect 11822 813 11856 847
rect 11856 813 11865 847
rect 11813 804 11865 813
rect 12017 1051 12069 1060
rect 12017 1017 12026 1051
rect 12026 1017 12060 1051
rect 12060 1017 12069 1051
rect 12017 1008 12069 1017
rect 12221 1255 12273 1264
rect 12221 1221 12230 1255
rect 12230 1221 12264 1255
rect 12264 1221 12273 1255
rect 12221 1212 12273 1221
rect 12425 1459 12477 1468
rect 12425 1425 12434 1459
rect 12434 1425 12468 1459
rect 12468 1425 12477 1459
rect 12425 1416 12477 1425
rect 12629 1663 12681 1672
rect 12629 1629 12638 1663
rect 12638 1629 12672 1663
rect 12672 1629 12681 1663
rect 12629 1620 12681 1629
rect 12833 1867 12885 1876
rect 12833 1833 12842 1867
rect 12842 1833 12876 1867
rect 12876 1833 12885 1867
rect 12833 1824 12885 1833
rect 13037 2071 13089 2080
rect 13037 2037 13046 2071
rect 13046 2037 13080 2071
rect 13080 2037 13089 2071
rect 13037 2028 13089 2037
rect 13241 643 13293 652
rect 13241 609 13250 643
rect 13250 609 13284 643
rect 13284 609 13293 643
rect 13241 600 13293 609
rect 13445 847 13497 856
rect 13445 813 13454 847
rect 13454 813 13488 847
rect 13488 813 13497 847
rect 13445 804 13497 813
rect 13649 1051 13701 1060
rect 13649 1017 13658 1051
rect 13658 1017 13692 1051
rect 13692 1017 13701 1051
rect 13649 1008 13701 1017
rect 13853 1255 13905 1264
rect 13853 1221 13862 1255
rect 13862 1221 13896 1255
rect 13896 1221 13905 1255
rect 13853 1212 13905 1221
rect 14057 1459 14109 1468
rect 14057 1425 14066 1459
rect 14066 1425 14100 1459
rect 14100 1425 14109 1459
rect 14057 1416 14109 1425
rect 14261 1663 14313 1672
rect 14261 1629 14270 1663
rect 14270 1629 14304 1663
rect 14304 1629 14313 1663
rect 14261 1620 14313 1629
rect 14465 1867 14517 1876
rect 14465 1833 14474 1867
rect 14474 1833 14508 1867
rect 14508 1833 14517 1867
rect 14465 1824 14517 1833
rect 14669 2071 14721 2080
rect 14669 2037 14678 2071
rect 14678 2037 14712 2071
rect 14712 2037 14721 2071
rect 14669 2028 14721 2037
rect 14873 643 14925 652
rect 14873 609 14882 643
rect 14882 609 14916 643
rect 14916 609 14925 643
rect 14873 600 14925 609
rect 15077 847 15129 856
rect 15077 813 15086 847
rect 15086 813 15120 847
rect 15120 813 15129 847
rect 15077 804 15129 813
rect 15281 1051 15333 1060
rect 15281 1017 15290 1051
rect 15290 1017 15324 1051
rect 15324 1017 15333 1051
rect 15281 1008 15333 1017
rect 15485 1255 15537 1264
rect 15485 1221 15494 1255
rect 15494 1221 15528 1255
rect 15528 1221 15537 1255
rect 15485 1212 15537 1221
rect 15689 1459 15741 1468
rect 15689 1425 15698 1459
rect 15698 1425 15732 1459
rect 15732 1425 15741 1459
rect 15689 1416 15741 1425
rect 15893 1663 15945 1672
rect 15893 1629 15902 1663
rect 15902 1629 15936 1663
rect 15936 1629 15945 1663
rect 15893 1620 15945 1629
rect 16097 1867 16149 1876
rect 16097 1833 16106 1867
rect 16106 1833 16140 1867
rect 16140 1833 16149 1867
rect 16097 1824 16149 1833
rect 16301 2071 16353 2080
rect 16301 2037 16310 2071
rect 16310 2037 16344 2071
rect 16344 2037 16353 2071
rect 16301 2028 16353 2037
rect 16505 643 16557 652
rect 16505 609 16514 643
rect 16514 609 16548 643
rect 16548 609 16557 643
rect 16505 600 16557 609
rect 16709 847 16761 856
rect 16709 813 16718 847
rect 16718 813 16752 847
rect 16752 813 16761 847
rect 16709 804 16761 813
rect 16913 1051 16965 1060
rect 16913 1017 16922 1051
rect 16922 1017 16956 1051
rect 16956 1017 16965 1051
rect 16913 1008 16965 1017
rect 17117 1255 17169 1264
rect 17117 1221 17126 1255
rect 17126 1221 17160 1255
rect 17160 1221 17169 1255
rect 17117 1212 17169 1221
rect 17321 1459 17373 1468
rect 17321 1425 17330 1459
rect 17330 1425 17364 1459
rect 17364 1425 17373 1459
rect 17321 1416 17373 1425
rect 17525 1663 17577 1672
rect 17525 1629 17534 1663
rect 17534 1629 17568 1663
rect 17568 1629 17577 1663
rect 17525 1620 17577 1629
rect 17729 1867 17781 1876
rect 17729 1833 17738 1867
rect 17738 1833 17772 1867
rect 17772 1833 17781 1867
rect 17729 1824 17781 1833
rect 17933 2071 17985 2080
rect 17933 2037 17942 2071
rect 17942 2037 17976 2071
rect 17976 2037 17985 2071
rect 17933 2028 17985 2037
rect 18137 643 18189 652
rect 18137 609 18146 643
rect 18146 609 18180 643
rect 18180 609 18189 643
rect 18137 600 18189 609
rect 18341 847 18393 856
rect 18341 813 18350 847
rect 18350 813 18384 847
rect 18384 813 18393 847
rect 18341 804 18393 813
rect 18545 1051 18597 1060
rect 18545 1017 18554 1051
rect 18554 1017 18588 1051
rect 18588 1017 18597 1051
rect 18545 1008 18597 1017
rect 18749 1255 18801 1264
rect 18749 1221 18758 1255
rect 18758 1221 18792 1255
rect 18792 1221 18801 1255
rect 18749 1212 18801 1221
rect 18953 1459 19005 1468
rect 18953 1425 18962 1459
rect 18962 1425 18996 1459
rect 18996 1425 19005 1459
rect 18953 1416 19005 1425
rect 19157 1663 19209 1672
rect 19157 1629 19166 1663
rect 19166 1629 19200 1663
rect 19200 1629 19209 1663
rect 19157 1620 19209 1629
rect 19361 1867 19413 1876
rect 19361 1833 19370 1867
rect 19370 1833 19404 1867
rect 19404 1833 19413 1867
rect 19361 1824 19413 1833
rect 19565 2071 19617 2080
rect 19565 2037 19574 2071
rect 19574 2037 19608 2071
rect 19608 2037 19617 2071
rect 19565 2028 19617 2037
rect 19769 643 19821 652
rect 19769 609 19778 643
rect 19778 609 19812 643
rect 19812 609 19821 643
rect 19769 600 19821 609
rect 19973 847 20025 856
rect 19973 813 19982 847
rect 19982 813 20016 847
rect 20016 813 20025 847
rect 19973 804 20025 813
rect 20177 1051 20229 1060
rect 20177 1017 20186 1051
rect 20186 1017 20220 1051
rect 20220 1017 20229 1051
rect 20177 1008 20229 1017
rect 20381 1255 20433 1264
rect 20381 1221 20390 1255
rect 20390 1221 20424 1255
rect 20424 1221 20433 1255
rect 20381 1212 20433 1221
rect 20585 1459 20637 1468
rect 20585 1425 20594 1459
rect 20594 1425 20628 1459
rect 20628 1425 20637 1459
rect 20585 1416 20637 1425
rect 20789 1663 20841 1672
rect 20789 1629 20798 1663
rect 20798 1629 20832 1663
rect 20832 1629 20841 1663
rect 20789 1620 20841 1629
rect 20993 1867 21045 1876
rect 20993 1833 21002 1867
rect 21002 1833 21036 1867
rect 21036 1833 21045 1867
rect 20993 1824 21045 1833
rect 21197 2071 21249 2080
rect 21197 2037 21206 2071
rect 21206 2037 21240 2071
rect 21240 2037 21249 2071
rect 21197 2028 21249 2037
rect 21401 643 21453 652
rect 21401 609 21410 643
rect 21410 609 21444 643
rect 21444 609 21453 643
rect 21401 600 21453 609
rect 21605 847 21657 856
rect 21605 813 21614 847
rect 21614 813 21648 847
rect 21648 813 21657 847
rect 21605 804 21657 813
rect 21809 1051 21861 1060
rect 21809 1017 21818 1051
rect 21818 1017 21852 1051
rect 21852 1017 21861 1051
rect 21809 1008 21861 1017
rect 22013 1255 22065 1264
rect 22013 1221 22022 1255
rect 22022 1221 22056 1255
rect 22056 1221 22065 1255
rect 22013 1212 22065 1221
rect 22217 1459 22269 1468
rect 22217 1425 22226 1459
rect 22226 1425 22260 1459
rect 22260 1425 22269 1459
rect 22217 1416 22269 1425
rect 22421 1663 22473 1672
rect 22421 1629 22430 1663
rect 22430 1629 22464 1663
rect 22464 1629 22473 1663
rect 22421 1620 22473 1629
rect 22625 1867 22677 1876
rect 22625 1833 22634 1867
rect 22634 1833 22668 1867
rect 22668 1833 22677 1867
rect 22625 1824 22677 1833
rect 22829 2071 22881 2080
rect 22829 2037 22838 2071
rect 22838 2037 22872 2071
rect 22872 2037 22881 2071
rect 22829 2028 22881 2037
rect 23033 643 23085 652
rect 23033 609 23042 643
rect 23042 609 23076 643
rect 23076 609 23085 643
rect 23033 600 23085 609
rect 23237 847 23289 856
rect 23237 813 23246 847
rect 23246 813 23280 847
rect 23280 813 23289 847
rect 23237 804 23289 813
rect 23441 1051 23493 1060
rect 23441 1017 23450 1051
rect 23450 1017 23484 1051
rect 23484 1017 23493 1051
rect 23441 1008 23493 1017
rect 23645 1255 23697 1264
rect 23645 1221 23654 1255
rect 23654 1221 23688 1255
rect 23688 1221 23697 1255
rect 23645 1212 23697 1221
rect 23849 1459 23901 1468
rect 23849 1425 23858 1459
rect 23858 1425 23892 1459
rect 23892 1425 23901 1459
rect 23849 1416 23901 1425
rect 24053 1663 24105 1672
rect 24053 1629 24062 1663
rect 24062 1629 24096 1663
rect 24096 1629 24105 1663
rect 24053 1620 24105 1629
rect 24257 1867 24309 1876
rect 24257 1833 24266 1867
rect 24266 1833 24300 1867
rect 24300 1833 24309 1867
rect 24257 1824 24309 1833
rect 24461 2071 24513 2080
rect 24461 2037 24470 2071
rect 24470 2037 24504 2071
rect 24504 2037 24513 2071
rect 24461 2028 24513 2037
rect 24665 643 24717 652
rect 24665 609 24674 643
rect 24674 609 24708 643
rect 24708 609 24717 643
rect 24665 600 24717 609
rect 24869 847 24921 856
rect 24869 813 24878 847
rect 24878 813 24912 847
rect 24912 813 24921 847
rect 24869 804 24921 813
rect 25073 1051 25125 1060
rect 25073 1017 25082 1051
rect 25082 1017 25116 1051
rect 25116 1017 25125 1051
rect 25073 1008 25125 1017
rect 25277 1255 25329 1264
rect 25277 1221 25286 1255
rect 25286 1221 25320 1255
rect 25320 1221 25329 1255
rect 25277 1212 25329 1221
rect 25481 1459 25533 1468
rect 25481 1425 25490 1459
rect 25490 1425 25524 1459
rect 25524 1425 25533 1459
rect 25481 1416 25533 1425
rect 25685 1663 25737 1672
rect 25685 1629 25694 1663
rect 25694 1629 25728 1663
rect 25728 1629 25737 1663
rect 25685 1620 25737 1629
rect 25889 1867 25941 1876
rect 25889 1833 25898 1867
rect 25898 1833 25932 1867
rect 25932 1833 25941 1867
rect 25889 1824 25941 1833
rect 26093 2071 26145 2080
rect 26093 2037 26102 2071
rect 26102 2037 26136 2071
rect 26136 2037 26145 2071
rect 26093 2028 26145 2037
rect 26297 643 26349 652
rect 26297 609 26306 643
rect 26306 609 26340 643
rect 26340 609 26349 643
rect 26297 600 26349 609
rect 26501 847 26553 856
rect 26501 813 26510 847
rect 26510 813 26544 847
rect 26544 813 26553 847
rect 26501 804 26553 813
rect 26705 1051 26757 1060
rect 26705 1017 26714 1051
rect 26714 1017 26748 1051
rect 26748 1017 26757 1051
rect 26705 1008 26757 1017
rect 26909 1255 26961 1264
rect 26909 1221 26918 1255
rect 26918 1221 26952 1255
rect 26952 1221 26961 1255
rect 26909 1212 26961 1221
rect 27113 1459 27165 1468
rect 27113 1425 27122 1459
rect 27122 1425 27156 1459
rect 27156 1425 27165 1459
rect 27113 1416 27165 1425
rect 27317 1663 27369 1672
rect 27317 1629 27326 1663
rect 27326 1629 27360 1663
rect 27360 1629 27369 1663
rect 27317 1620 27369 1629
rect 27521 1867 27573 1876
rect 27521 1833 27530 1867
rect 27530 1833 27564 1867
rect 27564 1833 27573 1867
rect 27521 1824 27573 1833
rect 27725 2071 27777 2080
rect 27725 2037 27734 2071
rect 27734 2037 27768 2071
rect 27768 2037 27777 2071
rect 27725 2028 27777 2037
rect 27929 643 27981 652
rect 27929 609 27938 643
rect 27938 609 27972 643
rect 27972 609 27981 643
rect 27929 600 27981 609
rect 28133 847 28185 856
rect 28133 813 28142 847
rect 28142 813 28176 847
rect 28176 813 28185 847
rect 28133 804 28185 813
rect 28337 1051 28389 1060
rect 28337 1017 28346 1051
rect 28346 1017 28380 1051
rect 28380 1017 28389 1051
rect 28337 1008 28389 1017
rect 28541 1255 28593 1264
rect 28541 1221 28550 1255
rect 28550 1221 28584 1255
rect 28584 1221 28593 1255
rect 28541 1212 28593 1221
rect 28745 1459 28797 1468
rect 28745 1425 28754 1459
rect 28754 1425 28788 1459
rect 28788 1425 28797 1459
rect 28745 1416 28797 1425
rect 28949 1663 29001 1672
rect 28949 1629 28958 1663
rect 28958 1629 28992 1663
rect 28992 1629 29001 1663
rect 28949 1620 29001 1629
rect 29153 1867 29205 1876
rect 29153 1833 29162 1867
rect 29162 1833 29196 1867
rect 29196 1833 29205 1867
rect 29153 1824 29205 1833
rect 29357 2071 29409 2080
rect 29357 2037 29366 2071
rect 29366 2037 29400 2071
rect 29400 2037 29409 2071
rect 29357 2028 29409 2037
rect 29561 643 29613 652
rect 29561 609 29570 643
rect 29570 609 29604 643
rect 29604 609 29613 643
rect 29561 600 29613 609
rect 29765 847 29817 856
rect 29765 813 29774 847
rect 29774 813 29808 847
rect 29808 813 29817 847
rect 29765 804 29817 813
rect 29969 1051 30021 1060
rect 29969 1017 29978 1051
rect 29978 1017 30012 1051
rect 30012 1017 30021 1051
rect 29969 1008 30021 1017
rect 30173 1255 30225 1264
rect 30173 1221 30182 1255
rect 30182 1221 30216 1255
rect 30216 1221 30225 1255
rect 30173 1212 30225 1221
rect 30377 1459 30429 1468
rect 30377 1425 30386 1459
rect 30386 1425 30420 1459
rect 30420 1425 30429 1459
rect 30377 1416 30429 1425
rect 30581 1663 30633 1672
rect 30581 1629 30590 1663
rect 30590 1629 30624 1663
rect 30624 1629 30633 1663
rect 30581 1620 30633 1629
rect 30785 1867 30837 1876
rect 30785 1833 30794 1867
rect 30794 1833 30828 1867
rect 30828 1833 30837 1867
rect 30785 1824 30837 1833
rect 30989 2071 31041 2080
rect 30989 2037 30998 2071
rect 30998 2037 31032 2071
rect 31032 2037 31041 2071
rect 30989 2028 31041 2037
rect 31193 643 31245 652
rect 31193 609 31202 643
rect 31202 609 31236 643
rect 31236 609 31245 643
rect 31193 600 31245 609
rect 31397 847 31449 856
rect 31397 813 31406 847
rect 31406 813 31440 847
rect 31440 813 31449 847
rect 31397 804 31449 813
rect 31601 1051 31653 1060
rect 31601 1017 31610 1051
rect 31610 1017 31644 1051
rect 31644 1017 31653 1051
rect 31601 1008 31653 1017
rect 31805 1255 31857 1264
rect 31805 1221 31814 1255
rect 31814 1221 31848 1255
rect 31848 1221 31857 1255
rect 31805 1212 31857 1221
rect 32009 1459 32061 1468
rect 32009 1425 32018 1459
rect 32018 1425 32052 1459
rect 32052 1425 32061 1459
rect 32009 1416 32061 1425
rect 32213 1663 32265 1672
rect 32213 1629 32222 1663
rect 32222 1629 32256 1663
rect 32256 1629 32265 1663
rect 32213 1620 32265 1629
rect 32417 1867 32469 1876
rect 32417 1833 32426 1867
rect 32426 1833 32460 1867
rect 32460 1833 32469 1867
rect 32417 1824 32469 1833
rect 32621 2071 32673 2080
rect 32621 2037 32630 2071
rect 32630 2037 32664 2071
rect 32664 2037 32673 2071
rect 32621 2028 32673 2037
rect 32825 643 32877 652
rect 32825 609 32834 643
rect 32834 609 32868 643
rect 32868 609 32877 643
rect 32825 600 32877 609
rect 33029 847 33081 856
rect 33029 813 33038 847
rect 33038 813 33072 847
rect 33072 813 33081 847
rect 33029 804 33081 813
rect 33233 1051 33285 1060
rect 33233 1017 33242 1051
rect 33242 1017 33276 1051
rect 33276 1017 33285 1051
rect 33233 1008 33285 1017
rect 33437 1255 33489 1264
rect 33437 1221 33446 1255
rect 33446 1221 33480 1255
rect 33480 1221 33489 1255
rect 33437 1212 33489 1221
rect 33641 1459 33693 1468
rect 33641 1425 33650 1459
rect 33650 1425 33684 1459
rect 33684 1425 33693 1459
rect 33641 1416 33693 1425
rect 33845 1663 33897 1672
rect 33845 1629 33854 1663
rect 33854 1629 33888 1663
rect 33888 1629 33897 1663
rect 33845 1620 33897 1629
rect 34049 1867 34101 1876
rect 34049 1833 34058 1867
rect 34058 1833 34092 1867
rect 34092 1833 34101 1867
rect 34049 1824 34101 1833
rect 34253 2071 34305 2080
rect 34253 2037 34262 2071
rect 34262 2037 34296 2071
rect 34296 2037 34305 2071
rect 34253 2028 34305 2037
rect 34457 643 34509 652
rect 34457 609 34466 643
rect 34466 609 34500 643
rect 34500 609 34509 643
rect 34457 600 34509 609
rect 34661 847 34713 856
rect 34661 813 34670 847
rect 34670 813 34704 847
rect 34704 813 34713 847
rect 34661 804 34713 813
rect 34865 1051 34917 1060
rect 34865 1017 34874 1051
rect 34874 1017 34908 1051
rect 34908 1017 34917 1051
rect 34865 1008 34917 1017
rect 35069 1255 35121 1264
rect 35069 1221 35078 1255
rect 35078 1221 35112 1255
rect 35112 1221 35121 1255
rect 35069 1212 35121 1221
rect 35273 1459 35325 1468
rect 35273 1425 35282 1459
rect 35282 1425 35316 1459
rect 35316 1425 35325 1459
rect 35273 1416 35325 1425
rect 35477 1663 35529 1672
rect 35477 1629 35486 1663
rect 35486 1629 35520 1663
rect 35520 1629 35529 1663
rect 35477 1620 35529 1629
rect 35681 1867 35733 1876
rect 35681 1833 35690 1867
rect 35690 1833 35724 1867
rect 35724 1833 35733 1867
rect 35681 1824 35733 1833
rect 35885 2071 35937 2080
rect 35885 2037 35894 2071
rect 35894 2037 35928 2071
rect 35928 2037 35937 2071
rect 35885 2028 35937 2037
rect 36089 643 36141 652
rect 36089 609 36098 643
rect 36098 609 36132 643
rect 36132 609 36141 643
rect 36089 600 36141 609
rect 36293 847 36345 856
rect 36293 813 36302 847
rect 36302 813 36336 847
rect 36336 813 36345 847
rect 36293 804 36345 813
rect 36497 1051 36549 1060
rect 36497 1017 36506 1051
rect 36506 1017 36540 1051
rect 36540 1017 36549 1051
rect 36497 1008 36549 1017
rect 36701 1255 36753 1264
rect 36701 1221 36710 1255
rect 36710 1221 36744 1255
rect 36744 1221 36753 1255
rect 36701 1212 36753 1221
rect 36905 1459 36957 1468
rect 36905 1425 36914 1459
rect 36914 1425 36948 1459
rect 36948 1425 36957 1459
rect 36905 1416 36957 1425
rect 37109 1663 37161 1672
rect 37109 1629 37118 1663
rect 37118 1629 37152 1663
rect 37152 1629 37161 1663
rect 37109 1620 37161 1629
rect 37313 1867 37365 1876
rect 37313 1833 37322 1867
rect 37322 1833 37356 1867
rect 37356 1833 37365 1867
rect 37313 1824 37365 1833
rect 37517 2071 37569 2080
rect 37517 2037 37526 2071
rect 37526 2037 37560 2071
rect 37560 2037 37569 2071
rect 37517 2028 37569 2037
rect 37721 643 37773 652
rect 37721 609 37730 643
rect 37730 609 37764 643
rect 37764 609 37773 643
rect 37721 600 37773 609
rect 37925 847 37977 856
rect 37925 813 37934 847
rect 37934 813 37968 847
rect 37968 813 37977 847
rect 37925 804 37977 813
rect 38129 1051 38181 1060
rect 38129 1017 38138 1051
rect 38138 1017 38172 1051
rect 38172 1017 38181 1051
rect 38129 1008 38181 1017
rect 38333 1255 38385 1264
rect 38333 1221 38342 1255
rect 38342 1221 38376 1255
rect 38376 1221 38385 1255
rect 38333 1212 38385 1221
rect 38537 1459 38589 1468
rect 38537 1425 38546 1459
rect 38546 1425 38580 1459
rect 38580 1425 38589 1459
rect 38537 1416 38589 1425
rect 38741 1663 38793 1672
rect 38741 1629 38750 1663
rect 38750 1629 38784 1663
rect 38784 1629 38793 1663
rect 38741 1620 38793 1629
rect 38945 1867 38997 1876
rect 38945 1833 38954 1867
rect 38954 1833 38988 1867
rect 38988 1833 38997 1867
rect 38945 1824 38997 1833
rect 39149 2071 39201 2080
rect 39149 2037 39158 2071
rect 39158 2037 39192 2071
rect 39192 2037 39201 2071
rect 39149 2028 39201 2037
rect 39353 643 39405 652
rect 39353 609 39362 643
rect 39362 609 39396 643
rect 39396 609 39405 643
rect 39353 600 39405 609
rect 39557 847 39609 856
rect 39557 813 39566 847
rect 39566 813 39600 847
rect 39600 813 39609 847
rect 39557 804 39609 813
rect 39761 1051 39813 1060
rect 39761 1017 39770 1051
rect 39770 1017 39804 1051
rect 39804 1017 39813 1051
rect 39761 1008 39813 1017
rect 39965 1255 40017 1264
rect 39965 1221 39974 1255
rect 39974 1221 40008 1255
rect 40008 1221 40017 1255
rect 39965 1212 40017 1221
rect 40169 1459 40221 1468
rect 40169 1425 40178 1459
rect 40178 1425 40212 1459
rect 40212 1425 40221 1459
rect 40169 1416 40221 1425
rect 40373 1663 40425 1672
rect 40373 1629 40382 1663
rect 40382 1629 40416 1663
rect 40416 1629 40425 1663
rect 40373 1620 40425 1629
rect 40577 1867 40629 1876
rect 40577 1833 40586 1867
rect 40586 1833 40620 1867
rect 40620 1833 40629 1867
rect 40577 1824 40629 1833
rect 40781 2071 40833 2080
rect 40781 2037 40790 2071
rect 40790 2037 40824 2071
rect 40824 2037 40833 2071
rect 40781 2028 40833 2037
rect 40985 643 41037 652
rect 40985 609 40994 643
rect 40994 609 41028 643
rect 41028 609 41037 643
rect 40985 600 41037 609
rect 41189 847 41241 856
rect 41189 813 41198 847
rect 41198 813 41232 847
rect 41232 813 41241 847
rect 41189 804 41241 813
rect 41393 1051 41445 1060
rect 41393 1017 41402 1051
rect 41402 1017 41436 1051
rect 41436 1017 41445 1051
rect 41393 1008 41445 1017
rect 41597 1255 41649 1264
rect 41597 1221 41606 1255
rect 41606 1221 41640 1255
rect 41640 1221 41649 1255
rect 41597 1212 41649 1221
rect 41801 1459 41853 1468
rect 41801 1425 41810 1459
rect 41810 1425 41844 1459
rect 41844 1425 41853 1459
rect 41801 1416 41853 1425
rect 42005 1663 42057 1672
rect 42005 1629 42014 1663
rect 42014 1629 42048 1663
rect 42048 1629 42057 1663
rect 42005 1620 42057 1629
rect 42209 1867 42261 1876
rect 42209 1833 42218 1867
rect 42218 1833 42252 1867
rect 42252 1833 42261 1867
rect 42209 1824 42261 1833
rect 42413 2071 42465 2080
rect 42413 2037 42422 2071
rect 42422 2037 42456 2071
rect 42456 2037 42465 2071
rect 42413 2028 42465 2037
rect 42617 643 42669 652
rect 42617 609 42626 643
rect 42626 609 42660 643
rect 42660 609 42669 643
rect 42617 600 42669 609
rect 42821 847 42873 856
rect 42821 813 42830 847
rect 42830 813 42864 847
rect 42864 813 42873 847
rect 42821 804 42873 813
rect 43025 1051 43077 1060
rect 43025 1017 43034 1051
rect 43034 1017 43068 1051
rect 43068 1017 43077 1051
rect 43025 1008 43077 1017
rect 43229 1255 43281 1264
rect 43229 1221 43238 1255
rect 43238 1221 43272 1255
rect 43272 1221 43281 1255
rect 43229 1212 43281 1221
rect 43433 1459 43485 1468
rect 43433 1425 43442 1459
rect 43442 1425 43476 1459
rect 43476 1425 43485 1459
rect 43433 1416 43485 1425
rect 43637 1663 43689 1672
rect 43637 1629 43646 1663
rect 43646 1629 43680 1663
rect 43680 1629 43689 1663
rect 43637 1620 43689 1629
rect 43841 1867 43893 1876
rect 43841 1833 43850 1867
rect 43850 1833 43884 1867
rect 43884 1833 43893 1867
rect 43841 1824 43893 1833
rect 44045 2071 44097 2080
rect 44045 2037 44054 2071
rect 44054 2037 44088 2071
rect 44088 2037 44097 2071
rect 44045 2028 44097 2037
rect 44249 643 44301 652
rect 44249 609 44258 643
rect 44258 609 44292 643
rect 44292 609 44301 643
rect 44249 600 44301 609
rect 44453 847 44505 856
rect 44453 813 44462 847
rect 44462 813 44496 847
rect 44496 813 44505 847
rect 44453 804 44505 813
rect 44657 1051 44709 1060
rect 44657 1017 44666 1051
rect 44666 1017 44700 1051
rect 44700 1017 44709 1051
rect 44657 1008 44709 1017
rect 44861 1255 44913 1264
rect 44861 1221 44870 1255
rect 44870 1221 44904 1255
rect 44904 1221 44913 1255
rect 44861 1212 44913 1221
rect 45065 1459 45117 1468
rect 45065 1425 45074 1459
rect 45074 1425 45108 1459
rect 45108 1425 45117 1459
rect 45065 1416 45117 1425
rect 45269 1663 45321 1672
rect 45269 1629 45278 1663
rect 45278 1629 45312 1663
rect 45312 1629 45321 1663
rect 45269 1620 45321 1629
rect 45473 1867 45525 1876
rect 45473 1833 45482 1867
rect 45482 1833 45516 1867
rect 45516 1833 45525 1867
rect 45473 1824 45525 1833
rect 45677 2071 45729 2080
rect 45677 2037 45686 2071
rect 45686 2037 45720 2071
rect 45720 2037 45729 2071
rect 45677 2028 45729 2037
rect 45881 643 45933 652
rect 45881 609 45890 643
rect 45890 609 45924 643
rect 45924 609 45933 643
rect 45881 600 45933 609
rect 46085 847 46137 856
rect 46085 813 46094 847
rect 46094 813 46128 847
rect 46128 813 46137 847
rect 46085 804 46137 813
rect 46289 1051 46341 1060
rect 46289 1017 46298 1051
rect 46298 1017 46332 1051
rect 46332 1017 46341 1051
rect 46289 1008 46341 1017
rect 46493 1255 46545 1264
rect 46493 1221 46502 1255
rect 46502 1221 46536 1255
rect 46536 1221 46545 1255
rect 46493 1212 46545 1221
rect 46697 1459 46749 1468
rect 46697 1425 46706 1459
rect 46706 1425 46740 1459
rect 46740 1425 46749 1459
rect 46697 1416 46749 1425
rect 46901 1663 46953 1672
rect 46901 1629 46910 1663
rect 46910 1629 46944 1663
rect 46944 1629 46953 1663
rect 46901 1620 46953 1629
rect 47105 1867 47157 1876
rect 47105 1833 47114 1867
rect 47114 1833 47148 1867
rect 47148 1833 47157 1867
rect 47105 1824 47157 1833
rect 47309 2071 47361 2080
rect 47309 2037 47318 2071
rect 47318 2037 47352 2071
rect 47352 2037 47361 2071
rect 47309 2028 47361 2037
rect 47513 643 47565 652
rect 47513 609 47522 643
rect 47522 609 47556 643
rect 47556 609 47565 643
rect 47513 600 47565 609
rect 47717 847 47769 856
rect 47717 813 47726 847
rect 47726 813 47760 847
rect 47760 813 47769 847
rect 47717 804 47769 813
rect 47921 1051 47973 1060
rect 47921 1017 47930 1051
rect 47930 1017 47964 1051
rect 47964 1017 47973 1051
rect 47921 1008 47973 1017
rect 48125 1255 48177 1264
rect 48125 1221 48134 1255
rect 48134 1221 48168 1255
rect 48168 1221 48177 1255
rect 48125 1212 48177 1221
rect 48329 1459 48381 1468
rect 48329 1425 48338 1459
rect 48338 1425 48372 1459
rect 48372 1425 48381 1459
rect 48329 1416 48381 1425
rect 48533 1663 48585 1672
rect 48533 1629 48542 1663
rect 48542 1629 48576 1663
rect 48576 1629 48585 1663
rect 48533 1620 48585 1629
rect 48737 1867 48789 1876
rect 48737 1833 48746 1867
rect 48746 1833 48780 1867
rect 48780 1833 48789 1867
rect 48737 1824 48789 1833
rect 48941 2071 48993 2080
rect 48941 2037 48950 2071
rect 48950 2037 48984 2071
rect 48984 2037 48993 2071
rect 48941 2028 48993 2037
rect 49145 643 49197 652
rect 49145 609 49154 643
rect 49154 609 49188 643
rect 49188 609 49197 643
rect 49145 600 49197 609
rect 49349 847 49401 856
rect 49349 813 49358 847
rect 49358 813 49392 847
rect 49392 813 49401 847
rect 49349 804 49401 813
rect 49553 1051 49605 1060
rect 49553 1017 49562 1051
rect 49562 1017 49596 1051
rect 49596 1017 49605 1051
rect 49553 1008 49605 1017
rect 49757 1255 49809 1264
rect 49757 1221 49766 1255
rect 49766 1221 49800 1255
rect 49800 1221 49809 1255
rect 49757 1212 49809 1221
rect 49961 1459 50013 1468
rect 49961 1425 49970 1459
rect 49970 1425 50004 1459
rect 50004 1425 50013 1459
rect 49961 1416 50013 1425
rect 50165 1663 50217 1672
rect 50165 1629 50174 1663
rect 50174 1629 50208 1663
rect 50208 1629 50217 1663
rect 50165 1620 50217 1629
rect 50369 1867 50421 1876
rect 50369 1833 50378 1867
rect 50378 1833 50412 1867
rect 50412 1833 50421 1867
rect 50369 1824 50421 1833
rect 50573 2071 50625 2080
rect 50573 2037 50582 2071
rect 50582 2037 50616 2071
rect 50616 2037 50625 2071
rect 50573 2028 50625 2037
rect 50777 643 50829 652
rect 50777 609 50786 643
rect 50786 609 50820 643
rect 50820 609 50829 643
rect 50777 600 50829 609
rect 50981 847 51033 856
rect 50981 813 50990 847
rect 50990 813 51024 847
rect 51024 813 51033 847
rect 50981 804 51033 813
rect 51185 1051 51237 1060
rect 51185 1017 51194 1051
rect 51194 1017 51228 1051
rect 51228 1017 51237 1051
rect 51185 1008 51237 1017
rect 51389 1255 51441 1264
rect 51389 1221 51398 1255
rect 51398 1221 51432 1255
rect 51432 1221 51441 1255
rect 51389 1212 51441 1221
rect 51593 1459 51645 1468
rect 51593 1425 51602 1459
rect 51602 1425 51636 1459
rect 51636 1425 51645 1459
rect 51593 1416 51645 1425
rect 51797 1663 51849 1672
rect 51797 1629 51806 1663
rect 51806 1629 51840 1663
rect 51840 1629 51849 1663
rect 51797 1620 51849 1629
rect 52001 1867 52053 1876
rect 52001 1833 52010 1867
rect 52010 1833 52044 1867
rect 52044 1833 52053 1867
rect 52001 1824 52053 1833
rect 52205 2071 52257 2080
rect 52205 2037 52214 2071
rect 52214 2037 52248 2071
rect 52248 2037 52257 2071
rect 52205 2028 52257 2037
rect 68 382 120 434
rect 272 382 324 434
rect 476 382 528 434
rect 680 382 732 434
rect 884 382 936 434
rect 1088 382 1140 434
rect 1292 382 1344 434
rect 1496 382 1548 434
rect 1700 382 1752 434
rect 1904 382 1956 434
rect 2108 382 2160 434
rect 2312 382 2364 434
rect 2516 382 2568 434
rect 2720 382 2772 434
rect 2924 382 2976 434
rect 3128 382 3180 434
rect 3332 382 3384 434
rect 3536 382 3588 434
rect 3740 382 3792 434
rect 3944 382 3996 434
rect 4148 382 4200 434
rect 4352 382 4404 434
rect 4556 382 4608 434
rect 4760 382 4812 434
rect 4964 382 5016 434
rect 5168 382 5220 434
rect 5372 382 5424 434
rect 5576 382 5628 434
rect 5780 382 5832 434
rect 5984 382 6036 434
rect 6188 382 6240 434
rect 6392 382 6444 434
rect 6596 382 6648 434
rect 6800 382 6852 434
rect 7004 382 7056 434
rect 7208 382 7260 434
rect 7412 382 7464 434
rect 7616 382 7668 434
rect 7820 382 7872 434
rect 8024 382 8076 434
rect 8228 382 8280 434
rect 8432 382 8484 434
rect 8636 382 8688 434
rect 8840 382 8892 434
rect 9044 382 9096 434
rect 9248 382 9300 434
rect 9452 382 9504 434
rect 9656 382 9708 434
rect 9860 382 9912 434
rect 10064 382 10116 434
rect 10268 382 10320 434
rect 10472 382 10524 434
rect 10676 382 10728 434
rect 10880 382 10932 434
rect 11084 382 11136 434
rect 11288 382 11340 434
rect 11492 382 11544 434
rect 11696 382 11748 434
rect 11900 382 11952 434
rect 12104 382 12156 434
rect 12308 382 12360 434
rect 12512 382 12564 434
rect 12716 382 12768 434
rect 12920 382 12972 434
rect 13124 382 13176 434
rect 13328 382 13380 434
rect 13532 382 13584 434
rect 13736 382 13788 434
rect 13940 382 13992 434
rect 14144 382 14196 434
rect 14348 382 14400 434
rect 14552 382 14604 434
rect 14756 382 14808 434
rect 14960 382 15012 434
rect 15164 382 15216 434
rect 15368 382 15420 434
rect 15572 382 15624 434
rect 15776 382 15828 434
rect 15980 382 16032 434
rect 16184 382 16236 434
rect 16388 382 16440 434
rect 16592 382 16644 434
rect 16796 382 16848 434
rect 17000 382 17052 434
rect 17204 382 17256 434
rect 17408 382 17460 434
rect 17612 382 17664 434
rect 17816 382 17868 434
rect 18020 382 18072 434
rect 18224 382 18276 434
rect 18428 382 18480 434
rect 18632 382 18684 434
rect 18836 382 18888 434
rect 19040 382 19092 434
rect 19244 382 19296 434
rect 19448 382 19500 434
rect 19652 382 19704 434
rect 19856 382 19908 434
rect 20060 382 20112 434
rect 20264 382 20316 434
rect 20468 382 20520 434
rect 20672 382 20724 434
rect 20876 382 20928 434
rect 21080 382 21132 434
rect 21284 382 21336 434
rect 21488 382 21540 434
rect 21692 382 21744 434
rect 21896 382 21948 434
rect 22100 382 22152 434
rect 22304 382 22356 434
rect 22508 382 22560 434
rect 22712 382 22764 434
rect 22916 382 22968 434
rect 23120 382 23172 434
rect 23324 382 23376 434
rect 23528 382 23580 434
rect 23732 382 23784 434
rect 23936 382 23988 434
rect 24140 382 24192 434
rect 24344 382 24396 434
rect 24548 382 24600 434
rect 24752 382 24804 434
rect 24956 382 25008 434
rect 25160 382 25212 434
rect 25364 382 25416 434
rect 25568 382 25620 434
rect 25772 382 25824 434
rect 25976 382 26028 434
rect 26180 382 26232 434
rect 26384 382 26436 434
rect 26588 382 26640 434
rect 26792 382 26844 434
rect 26996 382 27048 434
rect 27200 382 27252 434
rect 27404 382 27456 434
rect 27608 382 27660 434
rect 27812 382 27864 434
rect 28016 382 28068 434
rect 28220 382 28272 434
rect 28424 382 28476 434
rect 28628 382 28680 434
rect 28832 382 28884 434
rect 29036 382 29088 434
rect 29240 382 29292 434
rect 29444 382 29496 434
rect 29648 382 29700 434
rect 29852 382 29904 434
rect 30056 382 30108 434
rect 30260 382 30312 434
rect 30464 382 30516 434
rect 30668 382 30720 434
rect 30872 382 30924 434
rect 31076 382 31128 434
rect 31280 382 31332 434
rect 31484 382 31536 434
rect 31688 382 31740 434
rect 31892 382 31944 434
rect 32096 382 32148 434
rect 32300 382 32352 434
rect 32504 382 32556 434
rect 32708 382 32760 434
rect 32912 382 32964 434
rect 33116 382 33168 434
rect 33320 382 33372 434
rect 33524 382 33576 434
rect 33728 382 33780 434
rect 33932 382 33984 434
rect 34136 382 34188 434
rect 34340 382 34392 434
rect 34544 382 34596 434
rect 34748 382 34800 434
rect 34952 382 35004 434
rect 35156 382 35208 434
rect 35360 382 35412 434
rect 35564 382 35616 434
rect 35768 382 35820 434
rect 35972 382 36024 434
rect 36176 382 36228 434
rect 36380 382 36432 434
rect 36584 382 36636 434
rect 36788 382 36840 434
rect 36992 382 37044 434
rect 37196 382 37248 434
rect 37400 382 37452 434
rect 37604 382 37656 434
rect 37808 382 37860 434
rect 38012 382 38064 434
rect 38216 382 38268 434
rect 38420 382 38472 434
rect 38624 382 38676 434
rect 38828 382 38880 434
rect 39032 382 39084 434
rect 39236 382 39288 434
rect 39440 382 39492 434
rect 39644 382 39696 434
rect 39848 382 39900 434
rect 40052 382 40104 434
rect 40256 382 40308 434
rect 40460 382 40512 434
rect 40664 382 40716 434
rect 40868 382 40920 434
rect 41072 382 41124 434
rect 41276 382 41328 434
rect 41480 382 41532 434
rect 41684 382 41736 434
rect 41888 382 41940 434
rect 42092 382 42144 434
rect 42296 382 42348 434
rect 42500 382 42552 434
rect 42704 382 42756 434
rect 42908 382 42960 434
rect 43112 382 43164 434
rect 43316 382 43368 434
rect 43520 382 43572 434
rect 43724 382 43776 434
rect 43928 382 43980 434
rect 44132 382 44184 434
rect 44336 382 44388 434
rect 44540 382 44592 434
rect 44744 382 44796 434
rect 44948 382 45000 434
rect 45152 382 45204 434
rect 45356 382 45408 434
rect 45560 382 45612 434
rect 45764 382 45816 434
rect 45968 382 46020 434
rect 46172 382 46224 434
rect 46376 382 46428 434
rect 46580 382 46632 434
rect 46784 382 46836 434
rect 46988 382 47040 434
rect 47192 382 47244 434
rect 47396 382 47448 434
rect 47600 382 47652 434
rect 47804 382 47856 434
rect 48008 382 48060 434
rect 48212 382 48264 434
rect 48416 382 48468 434
rect 48620 382 48672 434
rect 48824 382 48876 434
rect 49028 382 49080 434
rect 49232 382 49284 434
rect 49436 382 49488 434
rect 49640 382 49692 434
rect 49844 382 49896 434
rect 50048 382 50100 434
rect 50252 382 50304 434
rect 50456 382 50508 434
rect 50660 382 50712 434
rect 50864 382 50916 434
rect 51068 382 51120 434
rect 51272 382 51324 434
rect 51476 382 51528 434
rect 51680 382 51732 434
rect 51884 382 51936 434
rect 52088 382 52140 434
<< metal2 >>
rect 26 3020 52264 3026
rect 26 2968 178 3020
rect 230 2968 382 3020
rect 434 2968 586 3020
rect 638 2968 790 3020
rect 842 2968 994 3020
rect 1046 2968 1198 3020
rect 1250 2968 1402 3020
rect 1454 2968 1606 3020
rect 1658 2968 1810 3020
rect 1862 2968 2014 3020
rect 2066 2968 2218 3020
rect 2270 2968 2422 3020
rect 2474 2968 2626 3020
rect 2678 2968 2830 3020
rect 2882 2968 3034 3020
rect 3086 2968 3238 3020
rect 3290 2968 3442 3020
rect 3494 2968 3646 3020
rect 3698 2968 3850 3020
rect 3902 2968 4054 3020
rect 4106 2968 4258 3020
rect 4310 2968 4462 3020
rect 4514 2968 4666 3020
rect 4718 2968 4870 3020
rect 4922 2968 5074 3020
rect 5126 2968 5278 3020
rect 5330 2968 5482 3020
rect 5534 2968 5686 3020
rect 5738 2968 5890 3020
rect 5942 2968 6094 3020
rect 6146 2968 6298 3020
rect 6350 2968 6502 3020
rect 6554 2968 6706 3020
rect 6758 2968 6910 3020
rect 6962 2968 7114 3020
rect 7166 2968 7318 3020
rect 7370 2968 7522 3020
rect 7574 2968 7726 3020
rect 7778 2968 7930 3020
rect 7982 2968 8134 3020
rect 8186 2968 8338 3020
rect 8390 2968 8542 3020
rect 8594 2968 8746 3020
rect 8798 2968 8950 3020
rect 9002 2968 9154 3020
rect 9206 2968 9358 3020
rect 9410 2968 9562 3020
rect 9614 2968 9766 3020
rect 9818 2968 9970 3020
rect 10022 2968 10174 3020
rect 10226 2968 10378 3020
rect 10430 2968 10582 3020
rect 10634 2968 10786 3020
rect 10838 2968 10990 3020
rect 11042 2968 11194 3020
rect 11246 2968 11398 3020
rect 11450 2968 11602 3020
rect 11654 2968 11806 3020
rect 11858 2968 12010 3020
rect 12062 2968 12214 3020
rect 12266 2968 12418 3020
rect 12470 2968 12622 3020
rect 12674 2968 12826 3020
rect 12878 2968 13030 3020
rect 13082 2968 13234 3020
rect 13286 2968 13438 3020
rect 13490 2968 13642 3020
rect 13694 2968 13846 3020
rect 13898 2968 14050 3020
rect 14102 2968 14254 3020
rect 14306 2968 14458 3020
rect 14510 2968 14662 3020
rect 14714 2968 14866 3020
rect 14918 2968 15070 3020
rect 15122 2968 15274 3020
rect 15326 2968 15478 3020
rect 15530 2968 15682 3020
rect 15734 2968 15886 3020
rect 15938 2968 16090 3020
rect 16142 2968 16294 3020
rect 16346 2968 16498 3020
rect 16550 2968 16702 3020
rect 16754 2968 16906 3020
rect 16958 2968 17110 3020
rect 17162 2968 17314 3020
rect 17366 2968 17518 3020
rect 17570 2968 17722 3020
rect 17774 2968 17926 3020
rect 17978 2968 18130 3020
rect 18182 2968 18334 3020
rect 18386 2968 18538 3020
rect 18590 2968 18742 3020
rect 18794 2968 18946 3020
rect 18998 2968 19150 3020
rect 19202 2968 19354 3020
rect 19406 2968 19558 3020
rect 19610 2968 19762 3020
rect 19814 2968 19966 3020
rect 20018 2968 20170 3020
rect 20222 2968 20374 3020
rect 20426 2968 20578 3020
rect 20630 2968 20782 3020
rect 20834 2968 20986 3020
rect 21038 2968 21190 3020
rect 21242 2968 21394 3020
rect 21446 2968 21598 3020
rect 21650 2968 21802 3020
rect 21854 2968 22006 3020
rect 22058 2968 22210 3020
rect 22262 2968 22414 3020
rect 22466 2968 22618 3020
rect 22670 2968 22822 3020
rect 22874 2968 23026 3020
rect 23078 2968 23230 3020
rect 23282 2968 23434 3020
rect 23486 2968 23638 3020
rect 23690 2968 23842 3020
rect 23894 2968 24046 3020
rect 24098 2968 24250 3020
rect 24302 2968 24454 3020
rect 24506 2968 24658 3020
rect 24710 2968 24862 3020
rect 24914 2968 25066 3020
rect 25118 2968 25270 3020
rect 25322 2968 25474 3020
rect 25526 2968 25678 3020
rect 25730 2968 25882 3020
rect 25934 2968 26086 3020
rect 26138 2968 26290 3020
rect 26342 2968 26494 3020
rect 26546 2968 26698 3020
rect 26750 2968 26902 3020
rect 26954 2968 27106 3020
rect 27158 2968 27310 3020
rect 27362 2968 27514 3020
rect 27566 2968 27718 3020
rect 27770 2968 27922 3020
rect 27974 2968 28126 3020
rect 28178 2968 28330 3020
rect 28382 2968 28534 3020
rect 28586 2968 28738 3020
rect 28790 2968 28942 3020
rect 28994 2968 29146 3020
rect 29198 2968 29350 3020
rect 29402 2968 29554 3020
rect 29606 2968 29758 3020
rect 29810 2968 29962 3020
rect 30014 2968 30166 3020
rect 30218 2968 30370 3020
rect 30422 2968 30574 3020
rect 30626 2968 30778 3020
rect 30830 2968 30982 3020
rect 31034 2968 31186 3020
rect 31238 2968 31390 3020
rect 31442 2968 31594 3020
rect 31646 2968 31798 3020
rect 31850 2968 32002 3020
rect 32054 2968 32206 3020
rect 32258 2968 32410 3020
rect 32462 2968 32614 3020
rect 32666 2968 32818 3020
rect 32870 2968 33022 3020
rect 33074 2968 33226 3020
rect 33278 2968 33430 3020
rect 33482 2968 33634 3020
rect 33686 2968 33838 3020
rect 33890 2968 34042 3020
rect 34094 2968 34246 3020
rect 34298 2968 34450 3020
rect 34502 2968 34654 3020
rect 34706 2968 34858 3020
rect 34910 2968 35062 3020
rect 35114 2968 35266 3020
rect 35318 2968 35470 3020
rect 35522 2968 35674 3020
rect 35726 2968 35878 3020
rect 35930 2968 36082 3020
rect 36134 2968 36286 3020
rect 36338 2968 36490 3020
rect 36542 2968 36694 3020
rect 36746 2968 36898 3020
rect 36950 2968 37102 3020
rect 37154 2968 37306 3020
rect 37358 2968 37510 3020
rect 37562 2968 37714 3020
rect 37766 2968 37918 3020
rect 37970 2968 38122 3020
rect 38174 2968 38326 3020
rect 38378 2968 38530 3020
rect 38582 2968 38734 3020
rect 38786 2968 38938 3020
rect 38990 2968 39142 3020
rect 39194 2968 39346 3020
rect 39398 2968 39550 3020
rect 39602 2968 39754 3020
rect 39806 2968 39958 3020
rect 40010 2968 40162 3020
rect 40214 2968 40366 3020
rect 40418 2968 40570 3020
rect 40622 2968 40774 3020
rect 40826 2968 40978 3020
rect 41030 2968 41182 3020
rect 41234 2968 41386 3020
rect 41438 2968 41590 3020
rect 41642 2968 41794 3020
rect 41846 2968 41998 3020
rect 42050 2968 42202 3020
rect 42254 2968 42406 3020
rect 42458 2968 42610 3020
rect 42662 2968 42814 3020
rect 42866 2968 43018 3020
rect 43070 2968 43222 3020
rect 43274 2968 43426 3020
rect 43478 2968 43630 3020
rect 43682 2968 43834 3020
rect 43886 2968 44038 3020
rect 44090 2968 44242 3020
rect 44294 2968 44446 3020
rect 44498 2968 44650 3020
rect 44702 2968 44854 3020
rect 44906 2968 45058 3020
rect 45110 2968 45262 3020
rect 45314 2968 45466 3020
rect 45518 2968 45670 3020
rect 45722 2968 45874 3020
rect 45926 2968 46078 3020
rect 46130 2968 46282 3020
rect 46334 2968 46486 3020
rect 46538 2968 46690 3020
rect 46742 2968 46894 3020
rect 46946 2968 47098 3020
rect 47150 2968 47302 3020
rect 47354 2968 47506 3020
rect 47558 2968 47710 3020
rect 47762 2968 47914 3020
rect 47966 2968 48118 3020
rect 48170 2968 48322 3020
rect 48374 2968 48526 3020
rect 48578 2968 48730 3020
rect 48782 2968 48934 3020
rect 48986 2968 49138 3020
rect 49190 2968 49342 3020
rect 49394 2968 49546 3020
rect 49598 2968 49750 3020
rect 49802 2968 49954 3020
rect 50006 2968 50158 3020
rect 50210 2968 50362 3020
rect 50414 2968 50566 3020
rect 50618 2968 50770 3020
rect 50822 2968 50974 3020
rect 51026 2968 51178 3020
rect 51230 2968 51382 3020
rect 51434 2968 51586 3020
rect 51638 2968 51790 3020
rect 51842 2968 51994 3020
rect 52046 2968 52198 3020
rect 52250 2968 52264 3020
rect 26 2962 52264 2968
rect 1607 2068 1613 2080
rect 0 2040 1613 2068
rect 1607 2028 1613 2040
rect 1665 2068 1671 2080
rect 3239 2068 3245 2080
rect 1665 2040 3245 2068
rect 1665 2028 1671 2040
rect 3239 2028 3245 2040
rect 3297 2068 3303 2080
rect 4871 2068 4877 2080
rect 3297 2040 4877 2068
rect 3297 2028 3303 2040
rect 4871 2028 4877 2040
rect 4929 2068 4935 2080
rect 6503 2068 6509 2080
rect 4929 2040 6509 2068
rect 4929 2028 4935 2040
rect 6503 2028 6509 2040
rect 6561 2068 6567 2080
rect 8135 2068 8141 2080
rect 6561 2040 8141 2068
rect 6561 2028 6567 2040
rect 8135 2028 8141 2040
rect 8193 2068 8199 2080
rect 9767 2068 9773 2080
rect 8193 2040 9773 2068
rect 8193 2028 8199 2040
rect 9767 2028 9773 2040
rect 9825 2068 9831 2080
rect 11399 2068 11405 2080
rect 9825 2040 11405 2068
rect 9825 2028 9831 2040
rect 11399 2028 11405 2040
rect 11457 2068 11463 2080
rect 13031 2068 13037 2080
rect 11457 2040 13037 2068
rect 11457 2028 11463 2040
rect 13031 2028 13037 2040
rect 13089 2068 13095 2080
rect 14663 2068 14669 2080
rect 13089 2040 14669 2068
rect 13089 2028 13095 2040
rect 14663 2028 14669 2040
rect 14721 2068 14727 2080
rect 16295 2068 16301 2080
rect 14721 2040 16301 2068
rect 14721 2028 14727 2040
rect 16295 2028 16301 2040
rect 16353 2068 16359 2080
rect 17927 2068 17933 2080
rect 16353 2040 17933 2068
rect 16353 2028 16359 2040
rect 17927 2028 17933 2040
rect 17985 2068 17991 2080
rect 19559 2068 19565 2080
rect 17985 2040 19565 2068
rect 17985 2028 17991 2040
rect 19559 2028 19565 2040
rect 19617 2068 19623 2080
rect 21191 2068 21197 2080
rect 19617 2040 21197 2068
rect 19617 2028 19623 2040
rect 21191 2028 21197 2040
rect 21249 2068 21255 2080
rect 22823 2068 22829 2080
rect 21249 2040 22829 2068
rect 21249 2028 21255 2040
rect 22823 2028 22829 2040
rect 22881 2068 22887 2080
rect 24455 2068 24461 2080
rect 22881 2040 24461 2068
rect 22881 2028 22887 2040
rect 24455 2028 24461 2040
rect 24513 2068 24519 2080
rect 26087 2068 26093 2080
rect 24513 2040 26093 2068
rect 24513 2028 24519 2040
rect 26087 2028 26093 2040
rect 26145 2068 26151 2080
rect 27719 2068 27725 2080
rect 26145 2040 27725 2068
rect 26145 2028 26151 2040
rect 27719 2028 27725 2040
rect 27777 2068 27783 2080
rect 29351 2068 29357 2080
rect 27777 2040 29357 2068
rect 27777 2028 27783 2040
rect 29351 2028 29357 2040
rect 29409 2068 29415 2080
rect 30983 2068 30989 2080
rect 29409 2040 30989 2068
rect 29409 2028 29415 2040
rect 30983 2028 30989 2040
rect 31041 2068 31047 2080
rect 32615 2068 32621 2080
rect 31041 2040 32621 2068
rect 31041 2028 31047 2040
rect 32615 2028 32621 2040
rect 32673 2068 32679 2080
rect 34247 2068 34253 2080
rect 32673 2040 34253 2068
rect 32673 2028 32679 2040
rect 34247 2028 34253 2040
rect 34305 2068 34311 2080
rect 35879 2068 35885 2080
rect 34305 2040 35885 2068
rect 34305 2028 34311 2040
rect 35879 2028 35885 2040
rect 35937 2068 35943 2080
rect 37511 2068 37517 2080
rect 35937 2040 37517 2068
rect 35937 2028 35943 2040
rect 37511 2028 37517 2040
rect 37569 2068 37575 2080
rect 39143 2068 39149 2080
rect 37569 2040 39149 2068
rect 37569 2028 37575 2040
rect 39143 2028 39149 2040
rect 39201 2068 39207 2080
rect 40775 2068 40781 2080
rect 39201 2040 40781 2068
rect 39201 2028 39207 2040
rect 40775 2028 40781 2040
rect 40833 2068 40839 2080
rect 42407 2068 42413 2080
rect 40833 2040 42413 2068
rect 40833 2028 40839 2040
rect 42407 2028 42413 2040
rect 42465 2068 42471 2080
rect 44039 2068 44045 2080
rect 42465 2040 44045 2068
rect 42465 2028 42471 2040
rect 44039 2028 44045 2040
rect 44097 2068 44103 2080
rect 45671 2068 45677 2080
rect 44097 2040 45677 2068
rect 44097 2028 44103 2040
rect 45671 2028 45677 2040
rect 45729 2068 45735 2080
rect 47303 2068 47309 2080
rect 45729 2040 47309 2068
rect 45729 2028 45735 2040
rect 47303 2028 47309 2040
rect 47361 2068 47367 2080
rect 48935 2068 48941 2080
rect 47361 2040 48941 2068
rect 47361 2028 47367 2040
rect 48935 2028 48941 2040
rect 48993 2068 48999 2080
rect 50567 2068 50573 2080
rect 48993 2040 50573 2068
rect 48993 2028 48999 2040
rect 50567 2028 50573 2040
rect 50625 2068 50631 2080
rect 52199 2068 52205 2080
rect 50625 2040 52205 2068
rect 50625 2028 50631 2040
rect 52199 2028 52205 2040
rect 52257 2028 52263 2080
rect 1403 1864 1409 1876
rect 0 1836 1409 1864
rect 1403 1824 1409 1836
rect 1461 1864 1467 1876
rect 3035 1864 3041 1876
rect 1461 1836 3041 1864
rect 1461 1824 1467 1836
rect 3035 1824 3041 1836
rect 3093 1864 3099 1876
rect 4667 1864 4673 1876
rect 3093 1836 4673 1864
rect 3093 1824 3099 1836
rect 4667 1824 4673 1836
rect 4725 1864 4731 1876
rect 6299 1864 6305 1876
rect 4725 1836 6305 1864
rect 4725 1824 4731 1836
rect 6299 1824 6305 1836
rect 6357 1864 6363 1876
rect 7931 1864 7937 1876
rect 6357 1836 7937 1864
rect 6357 1824 6363 1836
rect 7931 1824 7937 1836
rect 7989 1864 7995 1876
rect 9563 1864 9569 1876
rect 7989 1836 9569 1864
rect 7989 1824 7995 1836
rect 9563 1824 9569 1836
rect 9621 1864 9627 1876
rect 11195 1864 11201 1876
rect 9621 1836 11201 1864
rect 9621 1824 9627 1836
rect 11195 1824 11201 1836
rect 11253 1864 11259 1876
rect 12827 1864 12833 1876
rect 11253 1836 12833 1864
rect 11253 1824 11259 1836
rect 12827 1824 12833 1836
rect 12885 1864 12891 1876
rect 14459 1864 14465 1876
rect 12885 1836 14465 1864
rect 12885 1824 12891 1836
rect 14459 1824 14465 1836
rect 14517 1864 14523 1876
rect 16091 1864 16097 1876
rect 14517 1836 16097 1864
rect 14517 1824 14523 1836
rect 16091 1824 16097 1836
rect 16149 1864 16155 1876
rect 17723 1864 17729 1876
rect 16149 1836 17729 1864
rect 16149 1824 16155 1836
rect 17723 1824 17729 1836
rect 17781 1864 17787 1876
rect 19355 1864 19361 1876
rect 17781 1836 19361 1864
rect 17781 1824 17787 1836
rect 19355 1824 19361 1836
rect 19413 1864 19419 1876
rect 20987 1864 20993 1876
rect 19413 1836 20993 1864
rect 19413 1824 19419 1836
rect 20987 1824 20993 1836
rect 21045 1864 21051 1876
rect 22619 1864 22625 1876
rect 21045 1836 22625 1864
rect 21045 1824 21051 1836
rect 22619 1824 22625 1836
rect 22677 1864 22683 1876
rect 24251 1864 24257 1876
rect 22677 1836 24257 1864
rect 22677 1824 22683 1836
rect 24251 1824 24257 1836
rect 24309 1864 24315 1876
rect 25883 1864 25889 1876
rect 24309 1836 25889 1864
rect 24309 1824 24315 1836
rect 25883 1824 25889 1836
rect 25941 1864 25947 1876
rect 27515 1864 27521 1876
rect 25941 1836 27521 1864
rect 25941 1824 25947 1836
rect 27515 1824 27521 1836
rect 27573 1864 27579 1876
rect 29147 1864 29153 1876
rect 27573 1836 29153 1864
rect 27573 1824 27579 1836
rect 29147 1824 29153 1836
rect 29205 1864 29211 1876
rect 30779 1864 30785 1876
rect 29205 1836 30785 1864
rect 29205 1824 29211 1836
rect 30779 1824 30785 1836
rect 30837 1864 30843 1876
rect 32411 1864 32417 1876
rect 30837 1836 32417 1864
rect 30837 1824 30843 1836
rect 32411 1824 32417 1836
rect 32469 1864 32475 1876
rect 34043 1864 34049 1876
rect 32469 1836 34049 1864
rect 32469 1824 32475 1836
rect 34043 1824 34049 1836
rect 34101 1864 34107 1876
rect 35675 1864 35681 1876
rect 34101 1836 35681 1864
rect 34101 1824 34107 1836
rect 35675 1824 35681 1836
rect 35733 1864 35739 1876
rect 37307 1864 37313 1876
rect 35733 1836 37313 1864
rect 35733 1824 35739 1836
rect 37307 1824 37313 1836
rect 37365 1864 37371 1876
rect 38939 1864 38945 1876
rect 37365 1836 38945 1864
rect 37365 1824 37371 1836
rect 38939 1824 38945 1836
rect 38997 1864 39003 1876
rect 40571 1864 40577 1876
rect 38997 1836 40577 1864
rect 38997 1824 39003 1836
rect 40571 1824 40577 1836
rect 40629 1864 40635 1876
rect 42203 1864 42209 1876
rect 40629 1836 42209 1864
rect 40629 1824 40635 1836
rect 42203 1824 42209 1836
rect 42261 1864 42267 1876
rect 43835 1864 43841 1876
rect 42261 1836 43841 1864
rect 42261 1824 42267 1836
rect 43835 1824 43841 1836
rect 43893 1864 43899 1876
rect 45467 1864 45473 1876
rect 43893 1836 45473 1864
rect 43893 1824 43899 1836
rect 45467 1824 45473 1836
rect 45525 1864 45531 1876
rect 47099 1864 47105 1876
rect 45525 1836 47105 1864
rect 45525 1824 45531 1836
rect 47099 1824 47105 1836
rect 47157 1864 47163 1876
rect 48731 1864 48737 1876
rect 47157 1836 48737 1864
rect 47157 1824 47163 1836
rect 48731 1824 48737 1836
rect 48789 1864 48795 1876
rect 50363 1864 50369 1876
rect 48789 1836 50369 1864
rect 48789 1824 48795 1836
rect 50363 1824 50369 1836
rect 50421 1864 50427 1876
rect 51995 1864 52001 1876
rect 50421 1836 52001 1864
rect 50421 1824 50427 1836
rect 51995 1824 52001 1836
rect 52053 1864 52059 1876
rect 52053 1836 52224 1864
rect 52053 1824 52059 1836
rect 1199 1660 1205 1672
rect 0 1632 1205 1660
rect 1199 1620 1205 1632
rect 1257 1660 1263 1672
rect 2831 1660 2837 1672
rect 1257 1632 2837 1660
rect 1257 1620 1263 1632
rect 2831 1620 2837 1632
rect 2889 1660 2895 1672
rect 4463 1660 4469 1672
rect 2889 1632 4469 1660
rect 2889 1620 2895 1632
rect 4463 1620 4469 1632
rect 4521 1660 4527 1672
rect 6095 1660 6101 1672
rect 4521 1632 6101 1660
rect 4521 1620 4527 1632
rect 6095 1620 6101 1632
rect 6153 1660 6159 1672
rect 7727 1660 7733 1672
rect 6153 1632 7733 1660
rect 6153 1620 6159 1632
rect 7727 1620 7733 1632
rect 7785 1660 7791 1672
rect 9359 1660 9365 1672
rect 7785 1632 9365 1660
rect 7785 1620 7791 1632
rect 9359 1620 9365 1632
rect 9417 1660 9423 1672
rect 10991 1660 10997 1672
rect 9417 1632 10997 1660
rect 9417 1620 9423 1632
rect 10991 1620 10997 1632
rect 11049 1660 11055 1672
rect 12623 1660 12629 1672
rect 11049 1632 12629 1660
rect 11049 1620 11055 1632
rect 12623 1620 12629 1632
rect 12681 1660 12687 1672
rect 14255 1660 14261 1672
rect 12681 1632 14261 1660
rect 12681 1620 12687 1632
rect 14255 1620 14261 1632
rect 14313 1660 14319 1672
rect 15887 1660 15893 1672
rect 14313 1632 15893 1660
rect 14313 1620 14319 1632
rect 15887 1620 15893 1632
rect 15945 1660 15951 1672
rect 17519 1660 17525 1672
rect 15945 1632 17525 1660
rect 15945 1620 15951 1632
rect 17519 1620 17525 1632
rect 17577 1660 17583 1672
rect 19151 1660 19157 1672
rect 17577 1632 19157 1660
rect 17577 1620 17583 1632
rect 19151 1620 19157 1632
rect 19209 1660 19215 1672
rect 20783 1660 20789 1672
rect 19209 1632 20789 1660
rect 19209 1620 19215 1632
rect 20783 1620 20789 1632
rect 20841 1660 20847 1672
rect 22415 1660 22421 1672
rect 20841 1632 22421 1660
rect 20841 1620 20847 1632
rect 22415 1620 22421 1632
rect 22473 1660 22479 1672
rect 24047 1660 24053 1672
rect 22473 1632 24053 1660
rect 22473 1620 22479 1632
rect 24047 1620 24053 1632
rect 24105 1660 24111 1672
rect 25679 1660 25685 1672
rect 24105 1632 25685 1660
rect 24105 1620 24111 1632
rect 25679 1620 25685 1632
rect 25737 1660 25743 1672
rect 27311 1660 27317 1672
rect 25737 1632 27317 1660
rect 25737 1620 25743 1632
rect 27311 1620 27317 1632
rect 27369 1660 27375 1672
rect 28943 1660 28949 1672
rect 27369 1632 28949 1660
rect 27369 1620 27375 1632
rect 28943 1620 28949 1632
rect 29001 1660 29007 1672
rect 30575 1660 30581 1672
rect 29001 1632 30581 1660
rect 29001 1620 29007 1632
rect 30575 1620 30581 1632
rect 30633 1660 30639 1672
rect 32207 1660 32213 1672
rect 30633 1632 32213 1660
rect 30633 1620 30639 1632
rect 32207 1620 32213 1632
rect 32265 1660 32271 1672
rect 33839 1660 33845 1672
rect 32265 1632 33845 1660
rect 32265 1620 32271 1632
rect 33839 1620 33845 1632
rect 33897 1660 33903 1672
rect 35471 1660 35477 1672
rect 33897 1632 35477 1660
rect 33897 1620 33903 1632
rect 35471 1620 35477 1632
rect 35529 1660 35535 1672
rect 37103 1660 37109 1672
rect 35529 1632 37109 1660
rect 35529 1620 35535 1632
rect 37103 1620 37109 1632
rect 37161 1660 37167 1672
rect 38735 1660 38741 1672
rect 37161 1632 38741 1660
rect 37161 1620 37167 1632
rect 38735 1620 38741 1632
rect 38793 1660 38799 1672
rect 40367 1660 40373 1672
rect 38793 1632 40373 1660
rect 38793 1620 38799 1632
rect 40367 1620 40373 1632
rect 40425 1660 40431 1672
rect 41999 1660 42005 1672
rect 40425 1632 42005 1660
rect 40425 1620 40431 1632
rect 41999 1620 42005 1632
rect 42057 1660 42063 1672
rect 43631 1660 43637 1672
rect 42057 1632 43637 1660
rect 42057 1620 42063 1632
rect 43631 1620 43637 1632
rect 43689 1660 43695 1672
rect 45263 1660 45269 1672
rect 43689 1632 45269 1660
rect 43689 1620 43695 1632
rect 45263 1620 45269 1632
rect 45321 1660 45327 1672
rect 46895 1660 46901 1672
rect 45321 1632 46901 1660
rect 45321 1620 45327 1632
rect 46895 1620 46901 1632
rect 46953 1660 46959 1672
rect 48527 1660 48533 1672
rect 46953 1632 48533 1660
rect 46953 1620 46959 1632
rect 48527 1620 48533 1632
rect 48585 1660 48591 1672
rect 50159 1660 50165 1672
rect 48585 1632 50165 1660
rect 48585 1620 48591 1632
rect 50159 1620 50165 1632
rect 50217 1660 50223 1672
rect 51791 1660 51797 1672
rect 50217 1632 51797 1660
rect 50217 1620 50223 1632
rect 51791 1620 51797 1632
rect 51849 1660 51855 1672
rect 51849 1632 52224 1660
rect 51849 1620 51855 1632
rect 995 1456 1001 1468
rect 0 1428 1001 1456
rect 995 1416 1001 1428
rect 1053 1456 1059 1468
rect 2627 1456 2633 1468
rect 1053 1428 2633 1456
rect 1053 1416 1059 1428
rect 2627 1416 2633 1428
rect 2685 1456 2691 1468
rect 4259 1456 4265 1468
rect 2685 1428 4265 1456
rect 2685 1416 2691 1428
rect 4259 1416 4265 1428
rect 4317 1456 4323 1468
rect 5891 1456 5897 1468
rect 4317 1428 5897 1456
rect 4317 1416 4323 1428
rect 5891 1416 5897 1428
rect 5949 1456 5955 1468
rect 7523 1456 7529 1468
rect 5949 1428 7529 1456
rect 5949 1416 5955 1428
rect 7523 1416 7529 1428
rect 7581 1456 7587 1468
rect 9155 1456 9161 1468
rect 7581 1428 9161 1456
rect 7581 1416 7587 1428
rect 9155 1416 9161 1428
rect 9213 1456 9219 1468
rect 10787 1456 10793 1468
rect 9213 1428 10793 1456
rect 9213 1416 9219 1428
rect 10787 1416 10793 1428
rect 10845 1456 10851 1468
rect 12419 1456 12425 1468
rect 10845 1428 12425 1456
rect 10845 1416 10851 1428
rect 12419 1416 12425 1428
rect 12477 1456 12483 1468
rect 14051 1456 14057 1468
rect 12477 1428 14057 1456
rect 12477 1416 12483 1428
rect 14051 1416 14057 1428
rect 14109 1456 14115 1468
rect 15683 1456 15689 1468
rect 14109 1428 15689 1456
rect 14109 1416 14115 1428
rect 15683 1416 15689 1428
rect 15741 1456 15747 1468
rect 17315 1456 17321 1468
rect 15741 1428 17321 1456
rect 15741 1416 15747 1428
rect 17315 1416 17321 1428
rect 17373 1456 17379 1468
rect 18947 1456 18953 1468
rect 17373 1428 18953 1456
rect 17373 1416 17379 1428
rect 18947 1416 18953 1428
rect 19005 1456 19011 1468
rect 20579 1456 20585 1468
rect 19005 1428 20585 1456
rect 19005 1416 19011 1428
rect 20579 1416 20585 1428
rect 20637 1456 20643 1468
rect 22211 1456 22217 1468
rect 20637 1428 22217 1456
rect 20637 1416 20643 1428
rect 22211 1416 22217 1428
rect 22269 1456 22275 1468
rect 23843 1456 23849 1468
rect 22269 1428 23849 1456
rect 22269 1416 22275 1428
rect 23843 1416 23849 1428
rect 23901 1456 23907 1468
rect 25475 1456 25481 1468
rect 23901 1428 25481 1456
rect 23901 1416 23907 1428
rect 25475 1416 25481 1428
rect 25533 1456 25539 1468
rect 27107 1456 27113 1468
rect 25533 1428 27113 1456
rect 25533 1416 25539 1428
rect 27107 1416 27113 1428
rect 27165 1456 27171 1468
rect 28739 1456 28745 1468
rect 27165 1428 28745 1456
rect 27165 1416 27171 1428
rect 28739 1416 28745 1428
rect 28797 1456 28803 1468
rect 30371 1456 30377 1468
rect 28797 1428 30377 1456
rect 28797 1416 28803 1428
rect 30371 1416 30377 1428
rect 30429 1456 30435 1468
rect 32003 1456 32009 1468
rect 30429 1428 32009 1456
rect 30429 1416 30435 1428
rect 32003 1416 32009 1428
rect 32061 1456 32067 1468
rect 33635 1456 33641 1468
rect 32061 1428 33641 1456
rect 32061 1416 32067 1428
rect 33635 1416 33641 1428
rect 33693 1456 33699 1468
rect 35267 1456 35273 1468
rect 33693 1428 35273 1456
rect 33693 1416 33699 1428
rect 35267 1416 35273 1428
rect 35325 1456 35331 1468
rect 36899 1456 36905 1468
rect 35325 1428 36905 1456
rect 35325 1416 35331 1428
rect 36899 1416 36905 1428
rect 36957 1456 36963 1468
rect 38531 1456 38537 1468
rect 36957 1428 38537 1456
rect 36957 1416 36963 1428
rect 38531 1416 38537 1428
rect 38589 1456 38595 1468
rect 40163 1456 40169 1468
rect 38589 1428 40169 1456
rect 38589 1416 38595 1428
rect 40163 1416 40169 1428
rect 40221 1456 40227 1468
rect 41795 1456 41801 1468
rect 40221 1428 41801 1456
rect 40221 1416 40227 1428
rect 41795 1416 41801 1428
rect 41853 1456 41859 1468
rect 43427 1456 43433 1468
rect 41853 1428 43433 1456
rect 41853 1416 41859 1428
rect 43427 1416 43433 1428
rect 43485 1456 43491 1468
rect 45059 1456 45065 1468
rect 43485 1428 45065 1456
rect 43485 1416 43491 1428
rect 45059 1416 45065 1428
rect 45117 1456 45123 1468
rect 46691 1456 46697 1468
rect 45117 1428 46697 1456
rect 45117 1416 45123 1428
rect 46691 1416 46697 1428
rect 46749 1456 46755 1468
rect 48323 1456 48329 1468
rect 46749 1428 48329 1456
rect 46749 1416 46755 1428
rect 48323 1416 48329 1428
rect 48381 1456 48387 1468
rect 49955 1456 49961 1468
rect 48381 1428 49961 1456
rect 48381 1416 48387 1428
rect 49955 1416 49961 1428
rect 50013 1456 50019 1468
rect 51587 1456 51593 1468
rect 50013 1428 51593 1456
rect 50013 1416 50019 1428
rect 51587 1416 51593 1428
rect 51645 1456 51651 1468
rect 51645 1428 52224 1456
rect 51645 1416 51651 1428
rect 791 1252 797 1264
rect 0 1224 797 1252
rect 791 1212 797 1224
rect 849 1252 855 1264
rect 2423 1252 2429 1264
rect 849 1224 2429 1252
rect 849 1212 855 1224
rect 2423 1212 2429 1224
rect 2481 1252 2487 1264
rect 4055 1252 4061 1264
rect 2481 1224 4061 1252
rect 2481 1212 2487 1224
rect 4055 1212 4061 1224
rect 4113 1252 4119 1264
rect 5687 1252 5693 1264
rect 4113 1224 5693 1252
rect 4113 1212 4119 1224
rect 5687 1212 5693 1224
rect 5745 1252 5751 1264
rect 7319 1252 7325 1264
rect 5745 1224 7325 1252
rect 5745 1212 5751 1224
rect 7319 1212 7325 1224
rect 7377 1252 7383 1264
rect 8951 1252 8957 1264
rect 7377 1224 8957 1252
rect 7377 1212 7383 1224
rect 8951 1212 8957 1224
rect 9009 1252 9015 1264
rect 10583 1252 10589 1264
rect 9009 1224 10589 1252
rect 9009 1212 9015 1224
rect 10583 1212 10589 1224
rect 10641 1252 10647 1264
rect 12215 1252 12221 1264
rect 10641 1224 12221 1252
rect 10641 1212 10647 1224
rect 12215 1212 12221 1224
rect 12273 1252 12279 1264
rect 13847 1252 13853 1264
rect 12273 1224 13853 1252
rect 12273 1212 12279 1224
rect 13847 1212 13853 1224
rect 13905 1252 13911 1264
rect 15479 1252 15485 1264
rect 13905 1224 15485 1252
rect 13905 1212 13911 1224
rect 15479 1212 15485 1224
rect 15537 1252 15543 1264
rect 17111 1252 17117 1264
rect 15537 1224 17117 1252
rect 15537 1212 15543 1224
rect 17111 1212 17117 1224
rect 17169 1252 17175 1264
rect 18743 1252 18749 1264
rect 17169 1224 18749 1252
rect 17169 1212 17175 1224
rect 18743 1212 18749 1224
rect 18801 1252 18807 1264
rect 20375 1252 20381 1264
rect 18801 1224 20381 1252
rect 18801 1212 18807 1224
rect 20375 1212 20381 1224
rect 20433 1252 20439 1264
rect 22007 1252 22013 1264
rect 20433 1224 22013 1252
rect 20433 1212 20439 1224
rect 22007 1212 22013 1224
rect 22065 1252 22071 1264
rect 23639 1252 23645 1264
rect 22065 1224 23645 1252
rect 22065 1212 22071 1224
rect 23639 1212 23645 1224
rect 23697 1252 23703 1264
rect 25271 1252 25277 1264
rect 23697 1224 25277 1252
rect 23697 1212 23703 1224
rect 25271 1212 25277 1224
rect 25329 1252 25335 1264
rect 26903 1252 26909 1264
rect 25329 1224 26909 1252
rect 25329 1212 25335 1224
rect 26903 1212 26909 1224
rect 26961 1252 26967 1264
rect 28535 1252 28541 1264
rect 26961 1224 28541 1252
rect 26961 1212 26967 1224
rect 28535 1212 28541 1224
rect 28593 1252 28599 1264
rect 30167 1252 30173 1264
rect 28593 1224 30173 1252
rect 28593 1212 28599 1224
rect 30167 1212 30173 1224
rect 30225 1252 30231 1264
rect 31799 1252 31805 1264
rect 30225 1224 31805 1252
rect 30225 1212 30231 1224
rect 31799 1212 31805 1224
rect 31857 1252 31863 1264
rect 33431 1252 33437 1264
rect 31857 1224 33437 1252
rect 31857 1212 31863 1224
rect 33431 1212 33437 1224
rect 33489 1252 33495 1264
rect 35063 1252 35069 1264
rect 33489 1224 35069 1252
rect 33489 1212 33495 1224
rect 35063 1212 35069 1224
rect 35121 1252 35127 1264
rect 36695 1252 36701 1264
rect 35121 1224 36701 1252
rect 35121 1212 35127 1224
rect 36695 1212 36701 1224
rect 36753 1252 36759 1264
rect 38327 1252 38333 1264
rect 36753 1224 38333 1252
rect 36753 1212 36759 1224
rect 38327 1212 38333 1224
rect 38385 1252 38391 1264
rect 39959 1252 39965 1264
rect 38385 1224 39965 1252
rect 38385 1212 38391 1224
rect 39959 1212 39965 1224
rect 40017 1252 40023 1264
rect 41591 1252 41597 1264
rect 40017 1224 41597 1252
rect 40017 1212 40023 1224
rect 41591 1212 41597 1224
rect 41649 1252 41655 1264
rect 43223 1252 43229 1264
rect 41649 1224 43229 1252
rect 41649 1212 41655 1224
rect 43223 1212 43229 1224
rect 43281 1252 43287 1264
rect 44855 1252 44861 1264
rect 43281 1224 44861 1252
rect 43281 1212 43287 1224
rect 44855 1212 44861 1224
rect 44913 1252 44919 1264
rect 46487 1252 46493 1264
rect 44913 1224 46493 1252
rect 44913 1212 44919 1224
rect 46487 1212 46493 1224
rect 46545 1252 46551 1264
rect 48119 1252 48125 1264
rect 46545 1224 48125 1252
rect 46545 1212 46551 1224
rect 48119 1212 48125 1224
rect 48177 1252 48183 1264
rect 49751 1252 49757 1264
rect 48177 1224 49757 1252
rect 48177 1212 48183 1224
rect 49751 1212 49757 1224
rect 49809 1252 49815 1264
rect 51383 1252 51389 1264
rect 49809 1224 51389 1252
rect 49809 1212 49815 1224
rect 51383 1212 51389 1224
rect 51441 1252 51447 1264
rect 51441 1224 52224 1252
rect 51441 1212 51447 1224
rect 587 1048 593 1060
rect 0 1020 593 1048
rect 587 1008 593 1020
rect 645 1048 651 1060
rect 2219 1048 2225 1060
rect 645 1020 2225 1048
rect 645 1008 651 1020
rect 2219 1008 2225 1020
rect 2277 1048 2283 1060
rect 3851 1048 3857 1060
rect 2277 1020 3857 1048
rect 2277 1008 2283 1020
rect 3851 1008 3857 1020
rect 3909 1048 3915 1060
rect 5483 1048 5489 1060
rect 3909 1020 5489 1048
rect 3909 1008 3915 1020
rect 5483 1008 5489 1020
rect 5541 1048 5547 1060
rect 7115 1048 7121 1060
rect 5541 1020 7121 1048
rect 5541 1008 5547 1020
rect 7115 1008 7121 1020
rect 7173 1048 7179 1060
rect 8747 1048 8753 1060
rect 7173 1020 8753 1048
rect 7173 1008 7179 1020
rect 8747 1008 8753 1020
rect 8805 1048 8811 1060
rect 10379 1048 10385 1060
rect 8805 1020 10385 1048
rect 8805 1008 8811 1020
rect 10379 1008 10385 1020
rect 10437 1048 10443 1060
rect 12011 1048 12017 1060
rect 10437 1020 12017 1048
rect 10437 1008 10443 1020
rect 12011 1008 12017 1020
rect 12069 1048 12075 1060
rect 13643 1048 13649 1060
rect 12069 1020 13649 1048
rect 12069 1008 12075 1020
rect 13643 1008 13649 1020
rect 13701 1048 13707 1060
rect 15275 1048 15281 1060
rect 13701 1020 15281 1048
rect 13701 1008 13707 1020
rect 15275 1008 15281 1020
rect 15333 1048 15339 1060
rect 16907 1048 16913 1060
rect 15333 1020 16913 1048
rect 15333 1008 15339 1020
rect 16907 1008 16913 1020
rect 16965 1048 16971 1060
rect 18539 1048 18545 1060
rect 16965 1020 18545 1048
rect 16965 1008 16971 1020
rect 18539 1008 18545 1020
rect 18597 1048 18603 1060
rect 20171 1048 20177 1060
rect 18597 1020 20177 1048
rect 18597 1008 18603 1020
rect 20171 1008 20177 1020
rect 20229 1048 20235 1060
rect 21803 1048 21809 1060
rect 20229 1020 21809 1048
rect 20229 1008 20235 1020
rect 21803 1008 21809 1020
rect 21861 1048 21867 1060
rect 23435 1048 23441 1060
rect 21861 1020 23441 1048
rect 21861 1008 21867 1020
rect 23435 1008 23441 1020
rect 23493 1048 23499 1060
rect 25067 1048 25073 1060
rect 23493 1020 25073 1048
rect 23493 1008 23499 1020
rect 25067 1008 25073 1020
rect 25125 1048 25131 1060
rect 26699 1048 26705 1060
rect 25125 1020 26705 1048
rect 25125 1008 25131 1020
rect 26699 1008 26705 1020
rect 26757 1048 26763 1060
rect 28331 1048 28337 1060
rect 26757 1020 28337 1048
rect 26757 1008 26763 1020
rect 28331 1008 28337 1020
rect 28389 1048 28395 1060
rect 29963 1048 29969 1060
rect 28389 1020 29969 1048
rect 28389 1008 28395 1020
rect 29963 1008 29969 1020
rect 30021 1048 30027 1060
rect 31595 1048 31601 1060
rect 30021 1020 31601 1048
rect 30021 1008 30027 1020
rect 31595 1008 31601 1020
rect 31653 1048 31659 1060
rect 33227 1048 33233 1060
rect 31653 1020 33233 1048
rect 31653 1008 31659 1020
rect 33227 1008 33233 1020
rect 33285 1048 33291 1060
rect 34859 1048 34865 1060
rect 33285 1020 34865 1048
rect 33285 1008 33291 1020
rect 34859 1008 34865 1020
rect 34917 1048 34923 1060
rect 36491 1048 36497 1060
rect 34917 1020 36497 1048
rect 34917 1008 34923 1020
rect 36491 1008 36497 1020
rect 36549 1048 36555 1060
rect 38123 1048 38129 1060
rect 36549 1020 38129 1048
rect 36549 1008 36555 1020
rect 38123 1008 38129 1020
rect 38181 1048 38187 1060
rect 39755 1048 39761 1060
rect 38181 1020 39761 1048
rect 38181 1008 38187 1020
rect 39755 1008 39761 1020
rect 39813 1048 39819 1060
rect 41387 1048 41393 1060
rect 39813 1020 41393 1048
rect 39813 1008 39819 1020
rect 41387 1008 41393 1020
rect 41445 1048 41451 1060
rect 43019 1048 43025 1060
rect 41445 1020 43025 1048
rect 41445 1008 41451 1020
rect 43019 1008 43025 1020
rect 43077 1048 43083 1060
rect 44651 1048 44657 1060
rect 43077 1020 44657 1048
rect 43077 1008 43083 1020
rect 44651 1008 44657 1020
rect 44709 1048 44715 1060
rect 46283 1048 46289 1060
rect 44709 1020 46289 1048
rect 44709 1008 44715 1020
rect 46283 1008 46289 1020
rect 46341 1048 46347 1060
rect 47915 1048 47921 1060
rect 46341 1020 47921 1048
rect 46341 1008 46347 1020
rect 47915 1008 47921 1020
rect 47973 1048 47979 1060
rect 49547 1048 49553 1060
rect 47973 1020 49553 1048
rect 47973 1008 47979 1020
rect 49547 1008 49553 1020
rect 49605 1048 49611 1060
rect 51179 1048 51185 1060
rect 49605 1020 51185 1048
rect 49605 1008 49611 1020
rect 51179 1008 51185 1020
rect 51237 1048 51243 1060
rect 51237 1020 52224 1048
rect 51237 1008 51243 1020
rect 383 844 389 856
rect 0 816 389 844
rect 383 804 389 816
rect 441 844 447 856
rect 2015 844 2021 856
rect 441 816 2021 844
rect 441 804 447 816
rect 2015 804 2021 816
rect 2073 844 2079 856
rect 3647 844 3653 856
rect 2073 816 3653 844
rect 2073 804 2079 816
rect 3647 804 3653 816
rect 3705 844 3711 856
rect 5279 844 5285 856
rect 3705 816 5285 844
rect 3705 804 3711 816
rect 5279 804 5285 816
rect 5337 844 5343 856
rect 6911 844 6917 856
rect 5337 816 6917 844
rect 5337 804 5343 816
rect 6911 804 6917 816
rect 6969 844 6975 856
rect 8543 844 8549 856
rect 6969 816 8549 844
rect 6969 804 6975 816
rect 8543 804 8549 816
rect 8601 844 8607 856
rect 10175 844 10181 856
rect 8601 816 10181 844
rect 8601 804 8607 816
rect 10175 804 10181 816
rect 10233 844 10239 856
rect 11807 844 11813 856
rect 10233 816 11813 844
rect 10233 804 10239 816
rect 11807 804 11813 816
rect 11865 844 11871 856
rect 13439 844 13445 856
rect 11865 816 13445 844
rect 11865 804 11871 816
rect 13439 804 13445 816
rect 13497 844 13503 856
rect 15071 844 15077 856
rect 13497 816 15077 844
rect 13497 804 13503 816
rect 15071 804 15077 816
rect 15129 844 15135 856
rect 16703 844 16709 856
rect 15129 816 16709 844
rect 15129 804 15135 816
rect 16703 804 16709 816
rect 16761 844 16767 856
rect 18335 844 18341 856
rect 16761 816 18341 844
rect 16761 804 16767 816
rect 18335 804 18341 816
rect 18393 844 18399 856
rect 19967 844 19973 856
rect 18393 816 19973 844
rect 18393 804 18399 816
rect 19967 804 19973 816
rect 20025 844 20031 856
rect 21599 844 21605 856
rect 20025 816 21605 844
rect 20025 804 20031 816
rect 21599 804 21605 816
rect 21657 844 21663 856
rect 23231 844 23237 856
rect 21657 816 23237 844
rect 21657 804 21663 816
rect 23231 804 23237 816
rect 23289 844 23295 856
rect 24863 844 24869 856
rect 23289 816 24869 844
rect 23289 804 23295 816
rect 24863 804 24869 816
rect 24921 844 24927 856
rect 26495 844 26501 856
rect 24921 816 26501 844
rect 24921 804 24927 816
rect 26495 804 26501 816
rect 26553 844 26559 856
rect 28127 844 28133 856
rect 26553 816 28133 844
rect 26553 804 26559 816
rect 28127 804 28133 816
rect 28185 844 28191 856
rect 29759 844 29765 856
rect 28185 816 29765 844
rect 28185 804 28191 816
rect 29759 804 29765 816
rect 29817 844 29823 856
rect 31391 844 31397 856
rect 29817 816 31397 844
rect 29817 804 29823 816
rect 31391 804 31397 816
rect 31449 844 31455 856
rect 33023 844 33029 856
rect 31449 816 33029 844
rect 31449 804 31455 816
rect 33023 804 33029 816
rect 33081 844 33087 856
rect 34655 844 34661 856
rect 33081 816 34661 844
rect 33081 804 33087 816
rect 34655 804 34661 816
rect 34713 844 34719 856
rect 36287 844 36293 856
rect 34713 816 36293 844
rect 34713 804 34719 816
rect 36287 804 36293 816
rect 36345 844 36351 856
rect 37919 844 37925 856
rect 36345 816 37925 844
rect 36345 804 36351 816
rect 37919 804 37925 816
rect 37977 844 37983 856
rect 39551 844 39557 856
rect 37977 816 39557 844
rect 37977 804 37983 816
rect 39551 804 39557 816
rect 39609 844 39615 856
rect 41183 844 41189 856
rect 39609 816 41189 844
rect 39609 804 39615 816
rect 41183 804 41189 816
rect 41241 844 41247 856
rect 42815 844 42821 856
rect 41241 816 42821 844
rect 41241 804 41247 816
rect 42815 804 42821 816
rect 42873 844 42879 856
rect 44447 844 44453 856
rect 42873 816 44453 844
rect 42873 804 42879 816
rect 44447 804 44453 816
rect 44505 844 44511 856
rect 46079 844 46085 856
rect 44505 816 46085 844
rect 44505 804 44511 816
rect 46079 804 46085 816
rect 46137 844 46143 856
rect 47711 844 47717 856
rect 46137 816 47717 844
rect 46137 804 46143 816
rect 47711 804 47717 816
rect 47769 844 47775 856
rect 49343 844 49349 856
rect 47769 816 49349 844
rect 47769 804 47775 816
rect 49343 804 49349 816
rect 49401 844 49407 856
rect 50975 844 50981 856
rect 49401 816 50981 844
rect 49401 804 49407 816
rect 50975 804 50981 816
rect 51033 844 51039 856
rect 51033 816 52224 844
rect 51033 804 51039 816
rect 179 640 185 652
rect 0 612 185 640
rect 179 600 185 612
rect 237 640 243 652
rect 1811 640 1817 652
rect 237 612 1817 640
rect 237 600 243 612
rect 1811 600 1817 612
rect 1869 640 1875 652
rect 3443 640 3449 652
rect 1869 612 3449 640
rect 1869 600 1875 612
rect 3443 600 3449 612
rect 3501 640 3507 652
rect 5075 640 5081 652
rect 3501 612 5081 640
rect 3501 600 3507 612
rect 5075 600 5081 612
rect 5133 640 5139 652
rect 6707 640 6713 652
rect 5133 612 6713 640
rect 5133 600 5139 612
rect 6707 600 6713 612
rect 6765 640 6771 652
rect 8339 640 8345 652
rect 6765 612 8345 640
rect 6765 600 6771 612
rect 8339 600 8345 612
rect 8397 640 8403 652
rect 9971 640 9977 652
rect 8397 612 9977 640
rect 8397 600 8403 612
rect 9971 600 9977 612
rect 10029 640 10035 652
rect 11603 640 11609 652
rect 10029 612 11609 640
rect 10029 600 10035 612
rect 11603 600 11609 612
rect 11661 640 11667 652
rect 13235 640 13241 652
rect 11661 612 13241 640
rect 11661 600 11667 612
rect 13235 600 13241 612
rect 13293 640 13299 652
rect 14867 640 14873 652
rect 13293 612 14873 640
rect 13293 600 13299 612
rect 14867 600 14873 612
rect 14925 640 14931 652
rect 16499 640 16505 652
rect 14925 612 16505 640
rect 14925 600 14931 612
rect 16499 600 16505 612
rect 16557 640 16563 652
rect 18131 640 18137 652
rect 16557 612 18137 640
rect 16557 600 16563 612
rect 18131 600 18137 612
rect 18189 640 18195 652
rect 19763 640 19769 652
rect 18189 612 19769 640
rect 18189 600 18195 612
rect 19763 600 19769 612
rect 19821 640 19827 652
rect 21395 640 21401 652
rect 19821 612 21401 640
rect 19821 600 19827 612
rect 21395 600 21401 612
rect 21453 640 21459 652
rect 23027 640 23033 652
rect 21453 612 23033 640
rect 21453 600 21459 612
rect 23027 600 23033 612
rect 23085 640 23091 652
rect 24659 640 24665 652
rect 23085 612 24665 640
rect 23085 600 23091 612
rect 24659 600 24665 612
rect 24717 640 24723 652
rect 26291 640 26297 652
rect 24717 612 26297 640
rect 24717 600 24723 612
rect 26291 600 26297 612
rect 26349 640 26355 652
rect 27923 640 27929 652
rect 26349 612 27929 640
rect 26349 600 26355 612
rect 27923 600 27929 612
rect 27981 640 27987 652
rect 29555 640 29561 652
rect 27981 612 29561 640
rect 27981 600 27987 612
rect 29555 600 29561 612
rect 29613 640 29619 652
rect 31187 640 31193 652
rect 29613 612 31193 640
rect 29613 600 29619 612
rect 31187 600 31193 612
rect 31245 640 31251 652
rect 32819 640 32825 652
rect 31245 612 32825 640
rect 31245 600 31251 612
rect 32819 600 32825 612
rect 32877 640 32883 652
rect 34451 640 34457 652
rect 32877 612 34457 640
rect 32877 600 32883 612
rect 34451 600 34457 612
rect 34509 640 34515 652
rect 36083 640 36089 652
rect 34509 612 36089 640
rect 34509 600 34515 612
rect 36083 600 36089 612
rect 36141 640 36147 652
rect 37715 640 37721 652
rect 36141 612 37721 640
rect 36141 600 36147 612
rect 37715 600 37721 612
rect 37773 640 37779 652
rect 39347 640 39353 652
rect 37773 612 39353 640
rect 37773 600 37779 612
rect 39347 600 39353 612
rect 39405 640 39411 652
rect 40979 640 40985 652
rect 39405 612 40985 640
rect 39405 600 39411 612
rect 40979 600 40985 612
rect 41037 640 41043 652
rect 42611 640 42617 652
rect 41037 612 42617 640
rect 41037 600 41043 612
rect 42611 600 42617 612
rect 42669 640 42675 652
rect 44243 640 44249 652
rect 42669 612 44249 640
rect 42669 600 42675 612
rect 44243 600 44249 612
rect 44301 640 44307 652
rect 45875 640 45881 652
rect 44301 612 45881 640
rect 44301 600 44307 612
rect 45875 600 45881 612
rect 45933 640 45939 652
rect 47507 640 47513 652
rect 45933 612 47513 640
rect 45933 600 45939 612
rect 47507 600 47513 612
rect 47565 640 47571 652
rect 49139 640 49145 652
rect 47565 612 49145 640
rect 47565 600 47571 612
rect 49139 600 49145 612
rect 49197 640 49203 652
rect 50771 640 50777 652
rect 49197 612 50777 640
rect 49197 600 49203 612
rect 50771 600 50777 612
rect 50829 640 50835 652
rect 50829 612 52224 640
rect 50829 600 50835 612
rect 62 382 68 434
rect 120 422 126 434
rect 266 422 272 434
rect 120 394 272 422
rect 120 382 126 394
rect 266 382 272 394
rect 324 422 330 434
rect 470 422 476 434
rect 324 394 476 422
rect 324 382 330 394
rect 470 382 476 394
rect 528 422 534 434
rect 674 422 680 434
rect 528 394 680 422
rect 528 382 534 394
rect 674 382 680 394
rect 732 422 738 434
rect 878 422 884 434
rect 732 394 884 422
rect 732 382 738 394
rect 878 382 884 394
rect 936 422 942 434
rect 1082 422 1088 434
rect 936 394 1088 422
rect 936 382 942 394
rect 1082 382 1088 394
rect 1140 422 1146 434
rect 1286 422 1292 434
rect 1140 394 1292 422
rect 1140 382 1146 394
rect 1286 382 1292 394
rect 1344 422 1350 434
rect 1490 422 1496 434
rect 1344 394 1496 422
rect 1344 382 1350 394
rect 1490 382 1496 394
rect 1548 382 1554 434
rect 1694 382 1700 434
rect 1752 422 1758 434
rect 1898 422 1904 434
rect 1752 394 1904 422
rect 1752 382 1758 394
rect 1898 382 1904 394
rect 1956 422 1962 434
rect 2102 422 2108 434
rect 1956 394 2108 422
rect 1956 382 1962 394
rect 2102 382 2108 394
rect 2160 422 2166 434
rect 2306 422 2312 434
rect 2160 394 2312 422
rect 2160 382 2166 394
rect 2306 382 2312 394
rect 2364 422 2370 434
rect 2510 422 2516 434
rect 2364 394 2516 422
rect 2364 382 2370 394
rect 2510 382 2516 394
rect 2568 422 2574 434
rect 2714 422 2720 434
rect 2568 394 2720 422
rect 2568 382 2574 394
rect 2714 382 2720 394
rect 2772 422 2778 434
rect 2918 422 2924 434
rect 2772 394 2924 422
rect 2772 382 2778 394
rect 2918 382 2924 394
rect 2976 422 2982 434
rect 3122 422 3128 434
rect 2976 394 3128 422
rect 2976 382 2982 394
rect 3122 382 3128 394
rect 3180 382 3186 434
rect 3326 382 3332 434
rect 3384 422 3390 434
rect 3530 422 3536 434
rect 3384 394 3536 422
rect 3384 382 3390 394
rect 3530 382 3536 394
rect 3588 422 3594 434
rect 3734 422 3740 434
rect 3588 394 3740 422
rect 3588 382 3594 394
rect 3734 382 3740 394
rect 3792 422 3798 434
rect 3938 422 3944 434
rect 3792 394 3944 422
rect 3792 382 3798 394
rect 3938 382 3944 394
rect 3996 422 4002 434
rect 4142 422 4148 434
rect 3996 394 4148 422
rect 3996 382 4002 394
rect 4142 382 4148 394
rect 4200 422 4206 434
rect 4346 422 4352 434
rect 4200 394 4352 422
rect 4200 382 4206 394
rect 4346 382 4352 394
rect 4404 422 4410 434
rect 4550 422 4556 434
rect 4404 394 4556 422
rect 4404 382 4410 394
rect 4550 382 4556 394
rect 4608 422 4614 434
rect 4754 422 4760 434
rect 4608 394 4760 422
rect 4608 382 4614 394
rect 4754 382 4760 394
rect 4812 382 4818 434
rect 4958 382 4964 434
rect 5016 422 5022 434
rect 5162 422 5168 434
rect 5016 394 5168 422
rect 5016 382 5022 394
rect 5162 382 5168 394
rect 5220 422 5226 434
rect 5366 422 5372 434
rect 5220 394 5372 422
rect 5220 382 5226 394
rect 5366 382 5372 394
rect 5424 422 5430 434
rect 5570 422 5576 434
rect 5424 394 5576 422
rect 5424 382 5430 394
rect 5570 382 5576 394
rect 5628 422 5634 434
rect 5774 422 5780 434
rect 5628 394 5780 422
rect 5628 382 5634 394
rect 5774 382 5780 394
rect 5832 422 5838 434
rect 5978 422 5984 434
rect 5832 394 5984 422
rect 5832 382 5838 394
rect 5978 382 5984 394
rect 6036 422 6042 434
rect 6182 422 6188 434
rect 6036 394 6188 422
rect 6036 382 6042 394
rect 6182 382 6188 394
rect 6240 422 6246 434
rect 6386 422 6392 434
rect 6240 394 6392 422
rect 6240 382 6246 394
rect 6386 382 6392 394
rect 6444 382 6450 434
rect 6590 382 6596 434
rect 6648 422 6654 434
rect 6794 422 6800 434
rect 6648 394 6800 422
rect 6648 382 6654 394
rect 6794 382 6800 394
rect 6852 422 6858 434
rect 6998 422 7004 434
rect 6852 394 7004 422
rect 6852 382 6858 394
rect 6998 382 7004 394
rect 7056 422 7062 434
rect 7202 422 7208 434
rect 7056 394 7208 422
rect 7056 382 7062 394
rect 7202 382 7208 394
rect 7260 422 7266 434
rect 7406 422 7412 434
rect 7260 394 7412 422
rect 7260 382 7266 394
rect 7406 382 7412 394
rect 7464 422 7470 434
rect 7610 422 7616 434
rect 7464 394 7616 422
rect 7464 382 7470 394
rect 7610 382 7616 394
rect 7668 422 7674 434
rect 7814 422 7820 434
rect 7668 394 7820 422
rect 7668 382 7674 394
rect 7814 382 7820 394
rect 7872 422 7878 434
rect 8018 422 8024 434
rect 7872 394 8024 422
rect 7872 382 7878 394
rect 8018 382 8024 394
rect 8076 382 8082 434
rect 8222 382 8228 434
rect 8280 422 8286 434
rect 8426 422 8432 434
rect 8280 394 8432 422
rect 8280 382 8286 394
rect 8426 382 8432 394
rect 8484 422 8490 434
rect 8630 422 8636 434
rect 8484 394 8636 422
rect 8484 382 8490 394
rect 8630 382 8636 394
rect 8688 422 8694 434
rect 8834 422 8840 434
rect 8688 394 8840 422
rect 8688 382 8694 394
rect 8834 382 8840 394
rect 8892 422 8898 434
rect 9038 422 9044 434
rect 8892 394 9044 422
rect 8892 382 8898 394
rect 9038 382 9044 394
rect 9096 422 9102 434
rect 9242 422 9248 434
rect 9096 394 9248 422
rect 9096 382 9102 394
rect 9242 382 9248 394
rect 9300 422 9306 434
rect 9446 422 9452 434
rect 9300 394 9452 422
rect 9300 382 9306 394
rect 9446 382 9452 394
rect 9504 422 9510 434
rect 9650 422 9656 434
rect 9504 394 9656 422
rect 9504 382 9510 394
rect 9650 382 9656 394
rect 9708 382 9714 434
rect 9854 382 9860 434
rect 9912 422 9918 434
rect 10058 422 10064 434
rect 9912 394 10064 422
rect 9912 382 9918 394
rect 10058 382 10064 394
rect 10116 422 10122 434
rect 10262 422 10268 434
rect 10116 394 10268 422
rect 10116 382 10122 394
rect 10262 382 10268 394
rect 10320 422 10326 434
rect 10466 422 10472 434
rect 10320 394 10472 422
rect 10320 382 10326 394
rect 10466 382 10472 394
rect 10524 422 10530 434
rect 10670 422 10676 434
rect 10524 394 10676 422
rect 10524 382 10530 394
rect 10670 382 10676 394
rect 10728 422 10734 434
rect 10874 422 10880 434
rect 10728 394 10880 422
rect 10728 382 10734 394
rect 10874 382 10880 394
rect 10932 422 10938 434
rect 11078 422 11084 434
rect 10932 394 11084 422
rect 10932 382 10938 394
rect 11078 382 11084 394
rect 11136 422 11142 434
rect 11282 422 11288 434
rect 11136 394 11288 422
rect 11136 382 11142 394
rect 11282 382 11288 394
rect 11340 382 11346 434
rect 11486 382 11492 434
rect 11544 422 11550 434
rect 11690 422 11696 434
rect 11544 394 11696 422
rect 11544 382 11550 394
rect 11690 382 11696 394
rect 11748 422 11754 434
rect 11894 422 11900 434
rect 11748 394 11900 422
rect 11748 382 11754 394
rect 11894 382 11900 394
rect 11952 422 11958 434
rect 12098 422 12104 434
rect 11952 394 12104 422
rect 11952 382 11958 394
rect 12098 382 12104 394
rect 12156 422 12162 434
rect 12302 422 12308 434
rect 12156 394 12308 422
rect 12156 382 12162 394
rect 12302 382 12308 394
rect 12360 422 12366 434
rect 12506 422 12512 434
rect 12360 394 12512 422
rect 12360 382 12366 394
rect 12506 382 12512 394
rect 12564 422 12570 434
rect 12710 422 12716 434
rect 12564 394 12716 422
rect 12564 382 12570 394
rect 12710 382 12716 394
rect 12768 422 12774 434
rect 12914 422 12920 434
rect 12768 394 12920 422
rect 12768 382 12774 394
rect 12914 382 12920 394
rect 12972 382 12978 434
rect 13118 382 13124 434
rect 13176 422 13182 434
rect 13322 422 13328 434
rect 13176 394 13328 422
rect 13176 382 13182 394
rect 13322 382 13328 394
rect 13380 422 13386 434
rect 13526 422 13532 434
rect 13380 394 13532 422
rect 13380 382 13386 394
rect 13526 382 13532 394
rect 13584 422 13590 434
rect 13730 422 13736 434
rect 13584 394 13736 422
rect 13584 382 13590 394
rect 13730 382 13736 394
rect 13788 422 13794 434
rect 13934 422 13940 434
rect 13788 394 13940 422
rect 13788 382 13794 394
rect 13934 382 13940 394
rect 13992 422 13998 434
rect 14138 422 14144 434
rect 13992 394 14144 422
rect 13992 382 13998 394
rect 14138 382 14144 394
rect 14196 422 14202 434
rect 14342 422 14348 434
rect 14196 394 14348 422
rect 14196 382 14202 394
rect 14342 382 14348 394
rect 14400 422 14406 434
rect 14546 422 14552 434
rect 14400 394 14552 422
rect 14400 382 14406 394
rect 14546 382 14552 394
rect 14604 382 14610 434
rect 14750 382 14756 434
rect 14808 422 14814 434
rect 14954 422 14960 434
rect 14808 394 14960 422
rect 14808 382 14814 394
rect 14954 382 14960 394
rect 15012 422 15018 434
rect 15158 422 15164 434
rect 15012 394 15164 422
rect 15012 382 15018 394
rect 15158 382 15164 394
rect 15216 422 15222 434
rect 15362 422 15368 434
rect 15216 394 15368 422
rect 15216 382 15222 394
rect 15362 382 15368 394
rect 15420 422 15426 434
rect 15566 422 15572 434
rect 15420 394 15572 422
rect 15420 382 15426 394
rect 15566 382 15572 394
rect 15624 422 15630 434
rect 15770 422 15776 434
rect 15624 394 15776 422
rect 15624 382 15630 394
rect 15770 382 15776 394
rect 15828 422 15834 434
rect 15974 422 15980 434
rect 15828 394 15980 422
rect 15828 382 15834 394
rect 15974 382 15980 394
rect 16032 422 16038 434
rect 16178 422 16184 434
rect 16032 394 16184 422
rect 16032 382 16038 394
rect 16178 382 16184 394
rect 16236 382 16242 434
rect 16382 382 16388 434
rect 16440 422 16446 434
rect 16586 422 16592 434
rect 16440 394 16592 422
rect 16440 382 16446 394
rect 16586 382 16592 394
rect 16644 422 16650 434
rect 16790 422 16796 434
rect 16644 394 16796 422
rect 16644 382 16650 394
rect 16790 382 16796 394
rect 16848 422 16854 434
rect 16994 422 17000 434
rect 16848 394 17000 422
rect 16848 382 16854 394
rect 16994 382 17000 394
rect 17052 422 17058 434
rect 17198 422 17204 434
rect 17052 394 17204 422
rect 17052 382 17058 394
rect 17198 382 17204 394
rect 17256 422 17262 434
rect 17402 422 17408 434
rect 17256 394 17408 422
rect 17256 382 17262 394
rect 17402 382 17408 394
rect 17460 422 17466 434
rect 17606 422 17612 434
rect 17460 394 17612 422
rect 17460 382 17466 394
rect 17606 382 17612 394
rect 17664 422 17670 434
rect 17810 422 17816 434
rect 17664 394 17816 422
rect 17664 382 17670 394
rect 17810 382 17816 394
rect 17868 382 17874 434
rect 18014 382 18020 434
rect 18072 422 18078 434
rect 18218 422 18224 434
rect 18072 394 18224 422
rect 18072 382 18078 394
rect 18218 382 18224 394
rect 18276 422 18282 434
rect 18422 422 18428 434
rect 18276 394 18428 422
rect 18276 382 18282 394
rect 18422 382 18428 394
rect 18480 422 18486 434
rect 18626 422 18632 434
rect 18480 394 18632 422
rect 18480 382 18486 394
rect 18626 382 18632 394
rect 18684 422 18690 434
rect 18830 422 18836 434
rect 18684 394 18836 422
rect 18684 382 18690 394
rect 18830 382 18836 394
rect 18888 422 18894 434
rect 19034 422 19040 434
rect 18888 394 19040 422
rect 18888 382 18894 394
rect 19034 382 19040 394
rect 19092 422 19098 434
rect 19238 422 19244 434
rect 19092 394 19244 422
rect 19092 382 19098 394
rect 19238 382 19244 394
rect 19296 422 19302 434
rect 19442 422 19448 434
rect 19296 394 19448 422
rect 19296 382 19302 394
rect 19442 382 19448 394
rect 19500 382 19506 434
rect 19646 382 19652 434
rect 19704 422 19710 434
rect 19850 422 19856 434
rect 19704 394 19856 422
rect 19704 382 19710 394
rect 19850 382 19856 394
rect 19908 422 19914 434
rect 20054 422 20060 434
rect 19908 394 20060 422
rect 19908 382 19914 394
rect 20054 382 20060 394
rect 20112 422 20118 434
rect 20258 422 20264 434
rect 20112 394 20264 422
rect 20112 382 20118 394
rect 20258 382 20264 394
rect 20316 422 20322 434
rect 20462 422 20468 434
rect 20316 394 20468 422
rect 20316 382 20322 394
rect 20462 382 20468 394
rect 20520 422 20526 434
rect 20666 422 20672 434
rect 20520 394 20672 422
rect 20520 382 20526 394
rect 20666 382 20672 394
rect 20724 422 20730 434
rect 20870 422 20876 434
rect 20724 394 20876 422
rect 20724 382 20730 394
rect 20870 382 20876 394
rect 20928 422 20934 434
rect 21074 422 21080 434
rect 20928 394 21080 422
rect 20928 382 20934 394
rect 21074 382 21080 394
rect 21132 382 21138 434
rect 21278 382 21284 434
rect 21336 422 21342 434
rect 21482 422 21488 434
rect 21336 394 21488 422
rect 21336 382 21342 394
rect 21482 382 21488 394
rect 21540 422 21546 434
rect 21686 422 21692 434
rect 21540 394 21692 422
rect 21540 382 21546 394
rect 21686 382 21692 394
rect 21744 422 21750 434
rect 21890 422 21896 434
rect 21744 394 21896 422
rect 21744 382 21750 394
rect 21890 382 21896 394
rect 21948 422 21954 434
rect 22094 422 22100 434
rect 21948 394 22100 422
rect 21948 382 21954 394
rect 22094 382 22100 394
rect 22152 422 22158 434
rect 22298 422 22304 434
rect 22152 394 22304 422
rect 22152 382 22158 394
rect 22298 382 22304 394
rect 22356 422 22362 434
rect 22502 422 22508 434
rect 22356 394 22508 422
rect 22356 382 22362 394
rect 22502 382 22508 394
rect 22560 422 22566 434
rect 22706 422 22712 434
rect 22560 394 22712 422
rect 22560 382 22566 394
rect 22706 382 22712 394
rect 22764 382 22770 434
rect 22910 382 22916 434
rect 22968 422 22974 434
rect 23114 422 23120 434
rect 22968 394 23120 422
rect 22968 382 22974 394
rect 23114 382 23120 394
rect 23172 422 23178 434
rect 23318 422 23324 434
rect 23172 394 23324 422
rect 23172 382 23178 394
rect 23318 382 23324 394
rect 23376 422 23382 434
rect 23522 422 23528 434
rect 23376 394 23528 422
rect 23376 382 23382 394
rect 23522 382 23528 394
rect 23580 422 23586 434
rect 23726 422 23732 434
rect 23580 394 23732 422
rect 23580 382 23586 394
rect 23726 382 23732 394
rect 23784 422 23790 434
rect 23930 422 23936 434
rect 23784 394 23936 422
rect 23784 382 23790 394
rect 23930 382 23936 394
rect 23988 422 23994 434
rect 24134 422 24140 434
rect 23988 394 24140 422
rect 23988 382 23994 394
rect 24134 382 24140 394
rect 24192 422 24198 434
rect 24338 422 24344 434
rect 24192 394 24344 422
rect 24192 382 24198 394
rect 24338 382 24344 394
rect 24396 382 24402 434
rect 24542 382 24548 434
rect 24600 422 24606 434
rect 24746 422 24752 434
rect 24600 394 24752 422
rect 24600 382 24606 394
rect 24746 382 24752 394
rect 24804 422 24810 434
rect 24950 422 24956 434
rect 24804 394 24956 422
rect 24804 382 24810 394
rect 24950 382 24956 394
rect 25008 422 25014 434
rect 25154 422 25160 434
rect 25008 394 25160 422
rect 25008 382 25014 394
rect 25154 382 25160 394
rect 25212 422 25218 434
rect 25358 422 25364 434
rect 25212 394 25364 422
rect 25212 382 25218 394
rect 25358 382 25364 394
rect 25416 422 25422 434
rect 25562 422 25568 434
rect 25416 394 25568 422
rect 25416 382 25422 394
rect 25562 382 25568 394
rect 25620 422 25626 434
rect 25766 422 25772 434
rect 25620 394 25772 422
rect 25620 382 25626 394
rect 25766 382 25772 394
rect 25824 422 25830 434
rect 25970 422 25976 434
rect 25824 394 25976 422
rect 25824 382 25830 394
rect 25970 382 25976 394
rect 26028 382 26034 434
rect 26174 382 26180 434
rect 26232 422 26238 434
rect 26378 422 26384 434
rect 26232 394 26384 422
rect 26232 382 26238 394
rect 26378 382 26384 394
rect 26436 422 26442 434
rect 26582 422 26588 434
rect 26436 394 26588 422
rect 26436 382 26442 394
rect 26582 382 26588 394
rect 26640 422 26646 434
rect 26786 422 26792 434
rect 26640 394 26792 422
rect 26640 382 26646 394
rect 26786 382 26792 394
rect 26844 422 26850 434
rect 26990 422 26996 434
rect 26844 394 26996 422
rect 26844 382 26850 394
rect 26990 382 26996 394
rect 27048 422 27054 434
rect 27194 422 27200 434
rect 27048 394 27200 422
rect 27048 382 27054 394
rect 27194 382 27200 394
rect 27252 422 27258 434
rect 27398 422 27404 434
rect 27252 394 27404 422
rect 27252 382 27258 394
rect 27398 382 27404 394
rect 27456 422 27462 434
rect 27602 422 27608 434
rect 27456 394 27608 422
rect 27456 382 27462 394
rect 27602 382 27608 394
rect 27660 382 27666 434
rect 27806 382 27812 434
rect 27864 422 27870 434
rect 28010 422 28016 434
rect 27864 394 28016 422
rect 27864 382 27870 394
rect 28010 382 28016 394
rect 28068 422 28074 434
rect 28214 422 28220 434
rect 28068 394 28220 422
rect 28068 382 28074 394
rect 28214 382 28220 394
rect 28272 422 28278 434
rect 28418 422 28424 434
rect 28272 394 28424 422
rect 28272 382 28278 394
rect 28418 382 28424 394
rect 28476 422 28482 434
rect 28622 422 28628 434
rect 28476 394 28628 422
rect 28476 382 28482 394
rect 28622 382 28628 394
rect 28680 422 28686 434
rect 28826 422 28832 434
rect 28680 394 28832 422
rect 28680 382 28686 394
rect 28826 382 28832 394
rect 28884 422 28890 434
rect 29030 422 29036 434
rect 28884 394 29036 422
rect 28884 382 28890 394
rect 29030 382 29036 394
rect 29088 422 29094 434
rect 29234 422 29240 434
rect 29088 394 29240 422
rect 29088 382 29094 394
rect 29234 382 29240 394
rect 29292 382 29298 434
rect 29438 382 29444 434
rect 29496 422 29502 434
rect 29642 422 29648 434
rect 29496 394 29648 422
rect 29496 382 29502 394
rect 29642 382 29648 394
rect 29700 422 29706 434
rect 29846 422 29852 434
rect 29700 394 29852 422
rect 29700 382 29706 394
rect 29846 382 29852 394
rect 29904 422 29910 434
rect 30050 422 30056 434
rect 29904 394 30056 422
rect 29904 382 29910 394
rect 30050 382 30056 394
rect 30108 422 30114 434
rect 30254 422 30260 434
rect 30108 394 30260 422
rect 30108 382 30114 394
rect 30254 382 30260 394
rect 30312 422 30318 434
rect 30458 422 30464 434
rect 30312 394 30464 422
rect 30312 382 30318 394
rect 30458 382 30464 394
rect 30516 422 30522 434
rect 30662 422 30668 434
rect 30516 394 30668 422
rect 30516 382 30522 394
rect 30662 382 30668 394
rect 30720 422 30726 434
rect 30866 422 30872 434
rect 30720 394 30872 422
rect 30720 382 30726 394
rect 30866 382 30872 394
rect 30924 382 30930 434
rect 31070 382 31076 434
rect 31128 422 31134 434
rect 31274 422 31280 434
rect 31128 394 31280 422
rect 31128 382 31134 394
rect 31274 382 31280 394
rect 31332 422 31338 434
rect 31478 422 31484 434
rect 31332 394 31484 422
rect 31332 382 31338 394
rect 31478 382 31484 394
rect 31536 422 31542 434
rect 31682 422 31688 434
rect 31536 394 31688 422
rect 31536 382 31542 394
rect 31682 382 31688 394
rect 31740 422 31746 434
rect 31886 422 31892 434
rect 31740 394 31892 422
rect 31740 382 31746 394
rect 31886 382 31892 394
rect 31944 422 31950 434
rect 32090 422 32096 434
rect 31944 394 32096 422
rect 31944 382 31950 394
rect 32090 382 32096 394
rect 32148 422 32154 434
rect 32294 422 32300 434
rect 32148 394 32300 422
rect 32148 382 32154 394
rect 32294 382 32300 394
rect 32352 422 32358 434
rect 32498 422 32504 434
rect 32352 394 32504 422
rect 32352 382 32358 394
rect 32498 382 32504 394
rect 32556 382 32562 434
rect 32702 382 32708 434
rect 32760 422 32766 434
rect 32906 422 32912 434
rect 32760 394 32912 422
rect 32760 382 32766 394
rect 32906 382 32912 394
rect 32964 422 32970 434
rect 33110 422 33116 434
rect 32964 394 33116 422
rect 32964 382 32970 394
rect 33110 382 33116 394
rect 33168 422 33174 434
rect 33314 422 33320 434
rect 33168 394 33320 422
rect 33168 382 33174 394
rect 33314 382 33320 394
rect 33372 422 33378 434
rect 33518 422 33524 434
rect 33372 394 33524 422
rect 33372 382 33378 394
rect 33518 382 33524 394
rect 33576 422 33582 434
rect 33722 422 33728 434
rect 33576 394 33728 422
rect 33576 382 33582 394
rect 33722 382 33728 394
rect 33780 422 33786 434
rect 33926 422 33932 434
rect 33780 394 33932 422
rect 33780 382 33786 394
rect 33926 382 33932 394
rect 33984 422 33990 434
rect 34130 422 34136 434
rect 33984 394 34136 422
rect 33984 382 33990 394
rect 34130 382 34136 394
rect 34188 382 34194 434
rect 34334 382 34340 434
rect 34392 422 34398 434
rect 34538 422 34544 434
rect 34392 394 34544 422
rect 34392 382 34398 394
rect 34538 382 34544 394
rect 34596 422 34602 434
rect 34742 422 34748 434
rect 34596 394 34748 422
rect 34596 382 34602 394
rect 34742 382 34748 394
rect 34800 422 34806 434
rect 34946 422 34952 434
rect 34800 394 34952 422
rect 34800 382 34806 394
rect 34946 382 34952 394
rect 35004 422 35010 434
rect 35150 422 35156 434
rect 35004 394 35156 422
rect 35004 382 35010 394
rect 35150 382 35156 394
rect 35208 422 35214 434
rect 35354 422 35360 434
rect 35208 394 35360 422
rect 35208 382 35214 394
rect 35354 382 35360 394
rect 35412 422 35418 434
rect 35558 422 35564 434
rect 35412 394 35564 422
rect 35412 382 35418 394
rect 35558 382 35564 394
rect 35616 422 35622 434
rect 35762 422 35768 434
rect 35616 394 35768 422
rect 35616 382 35622 394
rect 35762 382 35768 394
rect 35820 382 35826 434
rect 35966 382 35972 434
rect 36024 422 36030 434
rect 36170 422 36176 434
rect 36024 394 36176 422
rect 36024 382 36030 394
rect 36170 382 36176 394
rect 36228 422 36234 434
rect 36374 422 36380 434
rect 36228 394 36380 422
rect 36228 382 36234 394
rect 36374 382 36380 394
rect 36432 422 36438 434
rect 36578 422 36584 434
rect 36432 394 36584 422
rect 36432 382 36438 394
rect 36578 382 36584 394
rect 36636 422 36642 434
rect 36782 422 36788 434
rect 36636 394 36788 422
rect 36636 382 36642 394
rect 36782 382 36788 394
rect 36840 422 36846 434
rect 36986 422 36992 434
rect 36840 394 36992 422
rect 36840 382 36846 394
rect 36986 382 36992 394
rect 37044 422 37050 434
rect 37190 422 37196 434
rect 37044 394 37196 422
rect 37044 382 37050 394
rect 37190 382 37196 394
rect 37248 422 37254 434
rect 37394 422 37400 434
rect 37248 394 37400 422
rect 37248 382 37254 394
rect 37394 382 37400 394
rect 37452 382 37458 434
rect 37598 382 37604 434
rect 37656 422 37662 434
rect 37802 422 37808 434
rect 37656 394 37808 422
rect 37656 382 37662 394
rect 37802 382 37808 394
rect 37860 422 37866 434
rect 38006 422 38012 434
rect 37860 394 38012 422
rect 37860 382 37866 394
rect 38006 382 38012 394
rect 38064 422 38070 434
rect 38210 422 38216 434
rect 38064 394 38216 422
rect 38064 382 38070 394
rect 38210 382 38216 394
rect 38268 422 38274 434
rect 38414 422 38420 434
rect 38268 394 38420 422
rect 38268 382 38274 394
rect 38414 382 38420 394
rect 38472 422 38478 434
rect 38618 422 38624 434
rect 38472 394 38624 422
rect 38472 382 38478 394
rect 38618 382 38624 394
rect 38676 422 38682 434
rect 38822 422 38828 434
rect 38676 394 38828 422
rect 38676 382 38682 394
rect 38822 382 38828 394
rect 38880 422 38886 434
rect 39026 422 39032 434
rect 38880 394 39032 422
rect 38880 382 38886 394
rect 39026 382 39032 394
rect 39084 382 39090 434
rect 39230 382 39236 434
rect 39288 422 39294 434
rect 39434 422 39440 434
rect 39288 394 39440 422
rect 39288 382 39294 394
rect 39434 382 39440 394
rect 39492 422 39498 434
rect 39638 422 39644 434
rect 39492 394 39644 422
rect 39492 382 39498 394
rect 39638 382 39644 394
rect 39696 422 39702 434
rect 39842 422 39848 434
rect 39696 394 39848 422
rect 39696 382 39702 394
rect 39842 382 39848 394
rect 39900 422 39906 434
rect 40046 422 40052 434
rect 39900 394 40052 422
rect 39900 382 39906 394
rect 40046 382 40052 394
rect 40104 422 40110 434
rect 40250 422 40256 434
rect 40104 394 40256 422
rect 40104 382 40110 394
rect 40250 382 40256 394
rect 40308 422 40314 434
rect 40454 422 40460 434
rect 40308 394 40460 422
rect 40308 382 40314 394
rect 40454 382 40460 394
rect 40512 422 40518 434
rect 40658 422 40664 434
rect 40512 394 40664 422
rect 40512 382 40518 394
rect 40658 382 40664 394
rect 40716 382 40722 434
rect 40862 382 40868 434
rect 40920 422 40926 434
rect 41066 422 41072 434
rect 40920 394 41072 422
rect 40920 382 40926 394
rect 41066 382 41072 394
rect 41124 422 41130 434
rect 41270 422 41276 434
rect 41124 394 41276 422
rect 41124 382 41130 394
rect 41270 382 41276 394
rect 41328 422 41334 434
rect 41474 422 41480 434
rect 41328 394 41480 422
rect 41328 382 41334 394
rect 41474 382 41480 394
rect 41532 422 41538 434
rect 41678 422 41684 434
rect 41532 394 41684 422
rect 41532 382 41538 394
rect 41678 382 41684 394
rect 41736 422 41742 434
rect 41882 422 41888 434
rect 41736 394 41888 422
rect 41736 382 41742 394
rect 41882 382 41888 394
rect 41940 422 41946 434
rect 42086 422 42092 434
rect 41940 394 42092 422
rect 41940 382 41946 394
rect 42086 382 42092 394
rect 42144 422 42150 434
rect 42290 422 42296 434
rect 42144 394 42296 422
rect 42144 382 42150 394
rect 42290 382 42296 394
rect 42348 382 42354 434
rect 42494 382 42500 434
rect 42552 422 42558 434
rect 42698 422 42704 434
rect 42552 394 42704 422
rect 42552 382 42558 394
rect 42698 382 42704 394
rect 42756 422 42762 434
rect 42902 422 42908 434
rect 42756 394 42908 422
rect 42756 382 42762 394
rect 42902 382 42908 394
rect 42960 422 42966 434
rect 43106 422 43112 434
rect 42960 394 43112 422
rect 42960 382 42966 394
rect 43106 382 43112 394
rect 43164 422 43170 434
rect 43310 422 43316 434
rect 43164 394 43316 422
rect 43164 382 43170 394
rect 43310 382 43316 394
rect 43368 422 43374 434
rect 43514 422 43520 434
rect 43368 394 43520 422
rect 43368 382 43374 394
rect 43514 382 43520 394
rect 43572 422 43578 434
rect 43718 422 43724 434
rect 43572 394 43724 422
rect 43572 382 43578 394
rect 43718 382 43724 394
rect 43776 422 43782 434
rect 43922 422 43928 434
rect 43776 394 43928 422
rect 43776 382 43782 394
rect 43922 382 43928 394
rect 43980 382 43986 434
rect 44126 382 44132 434
rect 44184 422 44190 434
rect 44330 422 44336 434
rect 44184 394 44336 422
rect 44184 382 44190 394
rect 44330 382 44336 394
rect 44388 422 44394 434
rect 44534 422 44540 434
rect 44388 394 44540 422
rect 44388 382 44394 394
rect 44534 382 44540 394
rect 44592 422 44598 434
rect 44738 422 44744 434
rect 44592 394 44744 422
rect 44592 382 44598 394
rect 44738 382 44744 394
rect 44796 422 44802 434
rect 44942 422 44948 434
rect 44796 394 44948 422
rect 44796 382 44802 394
rect 44942 382 44948 394
rect 45000 422 45006 434
rect 45146 422 45152 434
rect 45000 394 45152 422
rect 45000 382 45006 394
rect 45146 382 45152 394
rect 45204 422 45210 434
rect 45350 422 45356 434
rect 45204 394 45356 422
rect 45204 382 45210 394
rect 45350 382 45356 394
rect 45408 422 45414 434
rect 45554 422 45560 434
rect 45408 394 45560 422
rect 45408 382 45414 394
rect 45554 382 45560 394
rect 45612 382 45618 434
rect 45758 382 45764 434
rect 45816 422 45822 434
rect 45962 422 45968 434
rect 45816 394 45968 422
rect 45816 382 45822 394
rect 45962 382 45968 394
rect 46020 422 46026 434
rect 46166 422 46172 434
rect 46020 394 46172 422
rect 46020 382 46026 394
rect 46166 382 46172 394
rect 46224 422 46230 434
rect 46370 422 46376 434
rect 46224 394 46376 422
rect 46224 382 46230 394
rect 46370 382 46376 394
rect 46428 422 46434 434
rect 46574 422 46580 434
rect 46428 394 46580 422
rect 46428 382 46434 394
rect 46574 382 46580 394
rect 46632 422 46638 434
rect 46778 422 46784 434
rect 46632 394 46784 422
rect 46632 382 46638 394
rect 46778 382 46784 394
rect 46836 422 46842 434
rect 46982 422 46988 434
rect 46836 394 46988 422
rect 46836 382 46842 394
rect 46982 382 46988 394
rect 47040 422 47046 434
rect 47186 422 47192 434
rect 47040 394 47192 422
rect 47040 382 47046 394
rect 47186 382 47192 394
rect 47244 382 47250 434
rect 47390 382 47396 434
rect 47448 422 47454 434
rect 47594 422 47600 434
rect 47448 394 47600 422
rect 47448 382 47454 394
rect 47594 382 47600 394
rect 47652 422 47658 434
rect 47798 422 47804 434
rect 47652 394 47804 422
rect 47652 382 47658 394
rect 47798 382 47804 394
rect 47856 422 47862 434
rect 48002 422 48008 434
rect 47856 394 48008 422
rect 47856 382 47862 394
rect 48002 382 48008 394
rect 48060 422 48066 434
rect 48206 422 48212 434
rect 48060 394 48212 422
rect 48060 382 48066 394
rect 48206 382 48212 394
rect 48264 422 48270 434
rect 48410 422 48416 434
rect 48264 394 48416 422
rect 48264 382 48270 394
rect 48410 382 48416 394
rect 48468 422 48474 434
rect 48614 422 48620 434
rect 48468 394 48620 422
rect 48468 382 48474 394
rect 48614 382 48620 394
rect 48672 422 48678 434
rect 48818 422 48824 434
rect 48672 394 48824 422
rect 48672 382 48678 394
rect 48818 382 48824 394
rect 48876 382 48882 434
rect 49022 382 49028 434
rect 49080 422 49086 434
rect 49226 422 49232 434
rect 49080 394 49232 422
rect 49080 382 49086 394
rect 49226 382 49232 394
rect 49284 422 49290 434
rect 49430 422 49436 434
rect 49284 394 49436 422
rect 49284 382 49290 394
rect 49430 382 49436 394
rect 49488 422 49494 434
rect 49634 422 49640 434
rect 49488 394 49640 422
rect 49488 382 49494 394
rect 49634 382 49640 394
rect 49692 422 49698 434
rect 49838 422 49844 434
rect 49692 394 49844 422
rect 49692 382 49698 394
rect 49838 382 49844 394
rect 49896 422 49902 434
rect 50042 422 50048 434
rect 49896 394 50048 422
rect 49896 382 49902 394
rect 50042 382 50048 394
rect 50100 422 50106 434
rect 50246 422 50252 434
rect 50100 394 50252 422
rect 50100 382 50106 394
rect 50246 382 50252 394
rect 50304 422 50310 434
rect 50450 422 50456 434
rect 50304 394 50456 422
rect 50304 382 50310 394
rect 50450 382 50456 394
rect 50508 382 50514 434
rect 50654 382 50660 434
rect 50712 422 50718 434
rect 50858 422 50864 434
rect 50712 394 50864 422
rect 50712 382 50718 394
rect 50858 382 50864 394
rect 50916 422 50922 434
rect 51062 422 51068 434
rect 50916 394 51068 422
rect 50916 382 50922 394
rect 51062 382 51068 394
rect 51120 422 51126 434
rect 51266 422 51272 434
rect 51120 394 51272 422
rect 51120 382 51126 394
rect 51266 382 51272 394
rect 51324 422 51330 434
rect 51470 422 51476 434
rect 51324 394 51476 422
rect 51324 382 51330 394
rect 51470 382 51476 394
rect 51528 422 51534 434
rect 51674 422 51680 434
rect 51528 394 51680 422
rect 51528 382 51534 394
rect 51674 382 51680 394
rect 51732 422 51738 434
rect 51878 422 51884 434
rect 51732 394 51884 422
rect 51732 382 51738 394
rect 51878 382 51884 394
rect 51936 422 51942 434
rect 52082 422 52088 434
rect 51936 394 52088 422
rect 51936 382 51942 394
rect 52082 382 52088 394
rect 52140 382 52146 434
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_0
timestamp 1581449089
transform 1 0 52020 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_1
timestamp 1581449089
transform 1 0 51816 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_2
timestamp 1581449089
transform 1 0 51612 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_3
timestamp 1581449089
transform 1 0 51408 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_4
timestamp 1581449089
transform 1 0 51204 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_5
timestamp 1581449089
transform 1 0 51000 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_6
timestamp 1581449089
transform 1 0 50796 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_7
timestamp 1581449089
transform 1 0 50592 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_8
timestamp 1581449089
transform 1 0 50388 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_9
timestamp 1581449089
transform 1 0 50184 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_10
timestamp 1581449089
transform 1 0 49980 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_11
timestamp 1581449089
transform 1 0 49776 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_12
timestamp 1581449089
transform 1 0 49572 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_13
timestamp 1581449089
transform 1 0 49368 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_14
timestamp 1581449089
transform 1 0 49164 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_15
timestamp 1581449089
transform 1 0 48960 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_16
timestamp 1581449089
transform 1 0 48756 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_17
timestamp 1581449089
transform 1 0 48552 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_18
timestamp 1581449089
transform 1 0 48348 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_19
timestamp 1581449089
transform 1 0 48144 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_20
timestamp 1581449089
transform 1 0 47940 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_21
timestamp 1581449089
transform 1 0 47736 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_22
timestamp 1581449089
transform 1 0 47532 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_23
timestamp 1581449089
transform 1 0 47328 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_24
timestamp 1581449089
transform 1 0 47124 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_25
timestamp 1581449089
transform 1 0 46920 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_26
timestamp 1581449089
transform 1 0 46716 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_27
timestamp 1581449089
transform 1 0 46512 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_28
timestamp 1581449089
transform 1 0 46308 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_29
timestamp 1581449089
transform 1 0 46104 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_30
timestamp 1581449089
transform 1 0 45900 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_31
timestamp 1581449089
transform 1 0 45696 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_32
timestamp 1581449089
transform 1 0 45492 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_33
timestamp 1581449089
transform 1 0 45288 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_34
timestamp 1581449089
transform 1 0 45084 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_35
timestamp 1581449089
transform 1 0 44880 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_36
timestamp 1581449089
transform 1 0 44676 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_37
timestamp 1581449089
transform 1 0 44472 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_38
timestamp 1581449089
transform 1 0 44268 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_39
timestamp 1581449089
transform 1 0 44064 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_40
timestamp 1581449089
transform 1 0 43860 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_41
timestamp 1581449089
transform 1 0 43656 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_42
timestamp 1581449089
transform 1 0 43452 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_43
timestamp 1581449089
transform 1 0 43248 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_44
timestamp 1581449089
transform 1 0 43044 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_45
timestamp 1581449089
transform 1 0 42840 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_46
timestamp 1581449089
transform 1 0 42636 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_47
timestamp 1581449089
transform 1 0 42432 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_48
timestamp 1581449089
transform 1 0 42228 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_49
timestamp 1581449089
transform 1 0 42024 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_50
timestamp 1581449089
transform 1 0 41820 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_51
timestamp 1581449089
transform 1 0 41616 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_52
timestamp 1581449089
transform 1 0 41412 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_53
timestamp 1581449089
transform 1 0 41208 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_54
timestamp 1581449089
transform 1 0 41004 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_55
timestamp 1581449089
transform 1 0 40800 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_56
timestamp 1581449089
transform 1 0 40596 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_57
timestamp 1581449089
transform 1 0 40392 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_58
timestamp 1581449089
transform 1 0 40188 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_59
timestamp 1581449089
transform 1 0 39984 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_60
timestamp 1581449089
transform 1 0 39780 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_61
timestamp 1581449089
transform 1 0 39576 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_62
timestamp 1581449089
transform 1 0 39372 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_63
timestamp 1581449089
transform 1 0 39168 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_64
timestamp 1581449089
transform 1 0 38964 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_65
timestamp 1581449089
transform 1 0 38760 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_66
timestamp 1581449089
transform 1 0 38556 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_67
timestamp 1581449089
transform 1 0 38352 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_68
timestamp 1581449089
transform 1 0 38148 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_69
timestamp 1581449089
transform 1 0 37944 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_70
timestamp 1581449089
transform 1 0 37740 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_71
timestamp 1581449089
transform 1 0 37536 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_72
timestamp 1581449089
transform 1 0 37332 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_73
timestamp 1581449089
transform 1 0 37128 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_74
timestamp 1581449089
transform 1 0 36924 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_75
timestamp 1581449089
transform 1 0 36720 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_76
timestamp 1581449089
transform 1 0 36516 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_77
timestamp 1581449089
transform 1 0 36312 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_78
timestamp 1581449089
transform 1 0 36108 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_79
timestamp 1581449089
transform 1 0 35904 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_80
timestamp 1581449089
transform 1 0 35700 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_81
timestamp 1581449089
transform 1 0 35496 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_82
timestamp 1581449089
transform 1 0 35292 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_83
timestamp 1581449089
transform 1 0 35088 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_84
timestamp 1581449089
transform 1 0 34884 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_85
timestamp 1581449089
transform 1 0 34680 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_86
timestamp 1581449089
transform 1 0 34476 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_87
timestamp 1581449089
transform 1 0 34272 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_88
timestamp 1581449089
transform 1 0 34068 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_89
timestamp 1581449089
transform 1 0 33864 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_90
timestamp 1581449089
transform 1 0 33660 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_91
timestamp 1581449089
transform 1 0 33456 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_92
timestamp 1581449089
transform 1 0 33252 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_93
timestamp 1581449089
transform 1 0 33048 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_94
timestamp 1581449089
transform 1 0 32844 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_95
timestamp 1581449089
transform 1 0 32640 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_96
timestamp 1581449089
transform 1 0 32436 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_97
timestamp 1581449089
transform 1 0 32232 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_98
timestamp 1581449089
transform 1 0 32028 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_99
timestamp 1581449089
transform 1 0 31824 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_100
timestamp 1581449089
transform 1 0 31620 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_101
timestamp 1581449089
transform 1 0 31416 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_102
timestamp 1581449089
transform 1 0 31212 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_103
timestamp 1581449089
transform 1 0 31008 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_104
timestamp 1581449089
transform 1 0 30804 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_105
timestamp 1581449089
transform 1 0 30600 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_106
timestamp 1581449089
transform 1 0 30396 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_107
timestamp 1581449089
transform 1 0 30192 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_108
timestamp 1581449089
transform 1 0 29988 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_109
timestamp 1581449089
transform 1 0 29784 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_110
timestamp 1581449089
transform 1 0 29580 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_111
timestamp 1581449089
transform 1 0 29376 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_112
timestamp 1581449089
transform 1 0 29172 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_113
timestamp 1581449089
transform 1 0 28968 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_114
timestamp 1581449089
transform 1 0 28764 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_115
timestamp 1581449089
transform 1 0 28560 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_116
timestamp 1581449089
transform 1 0 28356 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_117
timestamp 1581449089
transform 1 0 28152 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_118
timestamp 1581449089
transform 1 0 27948 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_119
timestamp 1581449089
transform 1 0 27744 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_120
timestamp 1581449089
transform 1 0 27540 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_121
timestamp 1581449089
transform 1 0 27336 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_122
timestamp 1581449089
transform 1 0 27132 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_123
timestamp 1581449089
transform 1 0 26928 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_124
timestamp 1581449089
transform 1 0 26724 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_125
timestamp 1581449089
transform 1 0 26520 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_126
timestamp 1581449089
transform 1 0 26316 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_127
timestamp 1581449089
transform 1 0 26112 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_128
timestamp 1581449089
transform 1 0 25908 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_129
timestamp 1581449089
transform 1 0 25704 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_130
timestamp 1581449089
transform 1 0 25500 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_131
timestamp 1581449089
transform 1 0 25296 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_132
timestamp 1581449089
transform 1 0 25092 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_133
timestamp 1581449089
transform 1 0 24888 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_134
timestamp 1581449089
transform 1 0 24684 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_135
timestamp 1581449089
transform 1 0 24480 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_136
timestamp 1581449089
transform 1 0 24276 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_137
timestamp 1581449089
transform 1 0 24072 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_138
timestamp 1581449089
transform 1 0 23868 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_139
timestamp 1581449089
transform 1 0 23664 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_140
timestamp 1581449089
transform 1 0 23460 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_141
timestamp 1581449089
transform 1 0 23256 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_142
timestamp 1581449089
transform 1 0 23052 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_143
timestamp 1581449089
transform 1 0 22848 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_144
timestamp 1581449089
transform 1 0 22644 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_145
timestamp 1581449089
transform 1 0 22440 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_146
timestamp 1581449089
transform 1 0 22236 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_147
timestamp 1581449089
transform 1 0 22032 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_148
timestamp 1581449089
transform 1 0 21828 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_149
timestamp 1581449089
transform 1 0 21624 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_150
timestamp 1581449089
transform 1 0 21420 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_151
timestamp 1581449089
transform 1 0 21216 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_152
timestamp 1581449089
transform 1 0 21012 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_153
timestamp 1581449089
transform 1 0 20808 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_154
timestamp 1581449089
transform 1 0 20604 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_155
timestamp 1581449089
transform 1 0 20400 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_156
timestamp 1581449089
transform 1 0 20196 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_157
timestamp 1581449089
transform 1 0 19992 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_158
timestamp 1581449089
transform 1 0 19788 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_159
timestamp 1581449089
transform 1 0 19584 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_160
timestamp 1581449089
transform 1 0 19380 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_161
timestamp 1581449089
transform 1 0 19176 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_162
timestamp 1581449089
transform 1 0 18972 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_163
timestamp 1581449089
transform 1 0 18768 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_164
timestamp 1581449089
transform 1 0 18564 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_165
timestamp 1581449089
transform 1 0 18360 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_166
timestamp 1581449089
transform 1 0 18156 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_167
timestamp 1581449089
transform 1 0 17952 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_168
timestamp 1581449089
transform 1 0 17748 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_169
timestamp 1581449089
transform 1 0 17544 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_170
timestamp 1581449089
transform 1 0 17340 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_171
timestamp 1581449089
transform 1 0 17136 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_172
timestamp 1581449089
transform 1 0 16932 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_173
timestamp 1581449089
transform 1 0 16728 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_174
timestamp 1581449089
transform 1 0 16524 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_175
timestamp 1581449089
transform 1 0 16320 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_176
timestamp 1581449089
transform 1 0 16116 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_177
timestamp 1581449089
transform 1 0 15912 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_178
timestamp 1581449089
transform 1 0 15708 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_179
timestamp 1581449089
transform 1 0 15504 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_180
timestamp 1581449089
transform 1 0 15300 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_181
timestamp 1581449089
transform 1 0 15096 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_182
timestamp 1581449089
transform 1 0 14892 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_183
timestamp 1581449089
transform 1 0 14688 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_184
timestamp 1581449089
transform 1 0 14484 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_185
timestamp 1581449089
transform 1 0 14280 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_186
timestamp 1581449089
transform 1 0 14076 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_187
timestamp 1581449089
transform 1 0 13872 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_188
timestamp 1581449089
transform 1 0 13668 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_189
timestamp 1581449089
transform 1 0 13464 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_190
timestamp 1581449089
transform 1 0 13260 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_191
timestamp 1581449089
transform 1 0 13056 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_192
timestamp 1581449089
transform 1 0 12852 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_193
timestamp 1581449089
transform 1 0 12648 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_194
timestamp 1581449089
transform 1 0 12444 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_195
timestamp 1581449089
transform 1 0 12240 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_196
timestamp 1581449089
transform 1 0 12036 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_197
timestamp 1581449089
transform 1 0 11832 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_198
timestamp 1581449089
transform 1 0 11628 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_199
timestamp 1581449089
transform 1 0 11424 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_200
timestamp 1581449089
transform 1 0 11220 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_201
timestamp 1581449089
transform 1 0 11016 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_202
timestamp 1581449089
transform 1 0 10812 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_203
timestamp 1581449089
transform 1 0 10608 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_204
timestamp 1581449089
transform 1 0 10404 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_205
timestamp 1581449089
transform 1 0 10200 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_206
timestamp 1581449089
transform 1 0 9996 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_207
timestamp 1581449089
transform 1 0 9792 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_208
timestamp 1581449089
transform 1 0 9588 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_209
timestamp 1581449089
transform 1 0 9384 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_210
timestamp 1581449089
transform 1 0 9180 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_211
timestamp 1581449089
transform 1 0 8976 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_212
timestamp 1581449089
transform 1 0 8772 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_213
timestamp 1581449089
transform 1 0 8568 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_214
timestamp 1581449089
transform 1 0 8364 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_215
timestamp 1581449089
transform 1 0 8160 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_216
timestamp 1581449089
transform 1 0 7956 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_217
timestamp 1581449089
transform 1 0 7752 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_218
timestamp 1581449089
transform 1 0 7548 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_219
timestamp 1581449089
transform 1 0 7344 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_220
timestamp 1581449089
transform 1 0 7140 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_221
timestamp 1581449089
transform 1 0 6936 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_222
timestamp 1581449089
transform 1 0 6732 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_223
timestamp 1581449089
transform 1 0 6528 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_224
timestamp 1581449089
transform 1 0 6324 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_225
timestamp 1581449089
transform 1 0 6120 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_226
timestamp 1581449089
transform 1 0 5916 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_227
timestamp 1581449089
transform 1 0 5712 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_228
timestamp 1581449089
transform 1 0 5508 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_229
timestamp 1581449089
transform 1 0 5304 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_230
timestamp 1581449089
transform 1 0 5100 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_231
timestamp 1581449089
transform 1 0 4896 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_232
timestamp 1581449089
transform 1 0 4692 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_233
timestamp 1581449089
transform 1 0 4488 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_234
timestamp 1581449089
transform 1 0 4284 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_235
timestamp 1581449089
transform 1 0 4080 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_236
timestamp 1581449089
transform 1 0 3876 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_237
timestamp 1581449089
transform 1 0 3672 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_238
timestamp 1581449089
transform 1 0 3468 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_239
timestamp 1581449089
transform 1 0 3264 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_240
timestamp 1581449089
transform 1 0 3060 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_241
timestamp 1581449089
transform 1 0 2856 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_242
timestamp 1581449089
transform 1 0 2652 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_243
timestamp 1581449089
transform 1 0 2448 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_244
timestamp 1581449089
transform 1 0 2244 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_245
timestamp 1581449089
transform 1 0 2040 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_246
timestamp 1581449089
transform 1 0 1836 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_247
timestamp 1581449089
transform 1 0 1632 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_248
timestamp 1581449089
transform 1 0 1428 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_249
timestamp 1581449089
transform 1 0 1224 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_250
timestamp 1581449089
transform 1 0 1020 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_251
timestamp 1581449089
transform 1 0 816 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_252
timestamp 1581449089
transform 1 0 612 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_253
timestamp 1581449089
transform 1 0 408 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_254
timestamp 1581449089
transform 1 0 204 0 1 2244
box 1 0 255 817
use sky130_rom_krom_rom_column_mux  sky130_rom_krom_rom_column_mux_255
timestamp 1581449089
transform 1 0 0 0 1 2244
box 1 0 255 817
<< labels >>
rlabel metal2 s 0 612 52224 640 4 sel_0
port 3 nsew
rlabel metal2 s 0 816 52224 844 4 sel_1
port 5 nsew
rlabel metal2 s 0 1020 52224 1048 4 sel_2
port 7 nsew
rlabel metal2 s 0 1224 52224 1252 4 sel_3
port 9 nsew
rlabel metal2 s 0 1428 52224 1456 4 sel_4
port 11 nsew
rlabel metal2 s 0 1632 52224 1660 4 sel_5
port 13 nsew
rlabel metal2 s 0 1836 52224 1864 4 sel_6
port 15 nsew
rlabel metal2 s 0 2040 52224 2068 4 sel_7
port 17 nsew
rlabel metal1 s 80 408 108 2244 4 bl_out_0
port 19 nsew
rlabel metal1 s 1712 408 1740 2244 4 bl_out_1
port 21 nsew
rlabel metal1 s 3344 408 3372 2244 4 bl_out_2
port 23 nsew
rlabel metal1 s 4976 408 5004 2244 4 bl_out_3
port 25 nsew
rlabel metal1 s 6608 408 6636 2244 4 bl_out_4
port 27 nsew
rlabel metal1 s 8240 408 8268 2244 4 bl_out_5
port 29 nsew
rlabel metal1 s 9872 408 9900 2244 4 bl_out_6
port 31 nsew
rlabel metal1 s 11504 408 11532 2244 4 bl_out_7
port 33 nsew
rlabel metal1 s 13136 408 13164 2244 4 bl_out_8
port 35 nsew
rlabel metal1 s 14768 408 14796 2244 4 bl_out_9
port 37 nsew
rlabel metal1 s 16400 408 16428 2244 4 bl_out_10
port 39 nsew
rlabel metal1 s 18032 408 18060 2244 4 bl_out_11
port 41 nsew
rlabel metal1 s 19664 408 19692 2244 4 bl_out_12
port 43 nsew
rlabel metal1 s 21296 408 21324 2244 4 bl_out_13
port 45 nsew
rlabel metal1 s 22928 408 22956 2244 4 bl_out_14
port 47 nsew
rlabel metal1 s 24560 408 24588 2244 4 bl_out_15
port 49 nsew
rlabel metal1 s 26192 408 26220 2244 4 bl_out_16
port 51 nsew
rlabel metal1 s 27824 408 27852 2244 4 bl_out_17
port 53 nsew
rlabel metal1 s 29456 408 29484 2244 4 bl_out_18
port 55 nsew
rlabel metal1 s 31088 408 31116 2244 4 bl_out_19
port 57 nsew
rlabel metal1 s 32720 408 32748 2244 4 bl_out_20
port 59 nsew
rlabel metal1 s 34352 408 34380 2244 4 bl_out_21
port 61 nsew
rlabel metal1 s 35984 408 36012 2244 4 bl_out_22
port 63 nsew
rlabel metal1 s 37616 408 37644 2244 4 bl_out_23
port 65 nsew
rlabel metal1 s 39248 408 39276 2244 4 bl_out_24
port 67 nsew
rlabel metal1 s 40880 408 40908 2244 4 bl_out_25
port 69 nsew
rlabel metal1 s 42512 408 42540 2244 4 bl_out_26
port 71 nsew
rlabel metal1 s 44144 408 44172 2244 4 bl_out_27
port 73 nsew
rlabel metal1 s 45776 408 45804 2244 4 bl_out_28
port 75 nsew
rlabel metal1 s 47408 408 47436 2244 4 bl_out_29
port 77 nsew
rlabel metal1 s 49040 408 49068 2244 4 bl_out_30
port 79 nsew
rlabel metal1 s 50672 408 50700 2244 4 bl_out_31
port 81 nsew
rlabel metal2 s 26 2962 52264 3026 4 gnd
port 83 nsew
rlabel metal1 s 80 2874 108 3026 4 bl_0
port 85 nsew
rlabel metal1 s 284 2874 312 3026 4 bl_1
port 87 nsew
rlabel metal1 s 488 2874 516 3026 4 bl_2
port 89 nsew
rlabel metal1 s 692 2874 720 3026 4 bl_3
port 91 nsew
rlabel metal1 s 896 2874 924 3026 4 bl_4
port 93 nsew
rlabel metal1 s 1100 2874 1128 3026 4 bl_5
port 95 nsew
rlabel metal1 s 1304 2874 1332 3026 4 bl_6
port 97 nsew
rlabel metal1 s 1508 2874 1536 3026 4 bl_7
port 99 nsew
rlabel metal1 s 1712 2874 1740 3026 4 bl_8
port 101 nsew
rlabel metal1 s 1916 2874 1944 3026 4 bl_9
port 103 nsew
rlabel metal1 s 2120 2874 2148 3026 4 bl_10
port 105 nsew
rlabel metal1 s 2324 2874 2352 3026 4 bl_11
port 107 nsew
rlabel metal1 s 2528 2874 2556 3026 4 bl_12
port 109 nsew
rlabel metal1 s 2732 2874 2760 3026 4 bl_13
port 111 nsew
rlabel metal1 s 2936 2874 2964 3026 4 bl_14
port 113 nsew
rlabel metal1 s 3140 2874 3168 3026 4 bl_15
port 115 nsew
rlabel metal1 s 3344 2874 3372 3026 4 bl_16
port 117 nsew
rlabel metal1 s 3548 2874 3576 3026 4 bl_17
port 119 nsew
rlabel metal1 s 3752 2874 3780 3026 4 bl_18
port 121 nsew
rlabel metal1 s 3956 2874 3984 3026 4 bl_19
port 123 nsew
rlabel metal1 s 4160 2874 4188 3026 4 bl_20
port 125 nsew
rlabel metal1 s 4364 2874 4392 3026 4 bl_21
port 127 nsew
rlabel metal1 s 4568 2874 4596 3026 4 bl_22
port 129 nsew
rlabel metal1 s 4772 2874 4800 3026 4 bl_23
port 131 nsew
rlabel metal1 s 4976 2874 5004 3026 4 bl_24
port 133 nsew
rlabel metal1 s 5180 2874 5208 3026 4 bl_25
port 135 nsew
rlabel metal1 s 5384 2874 5412 3026 4 bl_26
port 137 nsew
rlabel metal1 s 5588 2874 5616 3026 4 bl_27
port 139 nsew
rlabel metal1 s 5792 2874 5820 3026 4 bl_28
port 141 nsew
rlabel metal1 s 5996 2874 6024 3026 4 bl_29
port 143 nsew
rlabel metal1 s 6200 2874 6228 3026 4 bl_30
port 145 nsew
rlabel metal1 s 6404 2874 6432 3026 4 bl_31
port 147 nsew
rlabel metal1 s 6608 2874 6636 3026 4 bl_32
port 149 nsew
rlabel metal1 s 6812 2874 6840 3026 4 bl_33
port 151 nsew
rlabel metal1 s 7016 2874 7044 3026 4 bl_34
port 153 nsew
rlabel metal1 s 7220 2874 7248 3026 4 bl_35
port 155 nsew
rlabel metal1 s 7424 2874 7452 3026 4 bl_36
port 157 nsew
rlabel metal1 s 7628 2874 7656 3026 4 bl_37
port 159 nsew
rlabel metal1 s 7832 2874 7860 3026 4 bl_38
port 161 nsew
rlabel metal1 s 8036 2874 8064 3026 4 bl_39
port 163 nsew
rlabel metal1 s 8240 2874 8268 3026 4 bl_40
port 165 nsew
rlabel metal1 s 8444 2874 8472 3026 4 bl_41
port 167 nsew
rlabel metal1 s 8648 2874 8676 3026 4 bl_42
port 169 nsew
rlabel metal1 s 8852 2874 8880 3026 4 bl_43
port 171 nsew
rlabel metal1 s 9056 2874 9084 3026 4 bl_44
port 173 nsew
rlabel metal1 s 9260 2874 9288 3026 4 bl_45
port 175 nsew
rlabel metal1 s 9464 2874 9492 3026 4 bl_46
port 177 nsew
rlabel metal1 s 9668 2874 9696 3026 4 bl_47
port 179 nsew
rlabel metal1 s 9872 2874 9900 3026 4 bl_48
port 181 nsew
rlabel metal1 s 10076 2874 10104 3026 4 bl_49
port 183 nsew
rlabel metal1 s 10280 2874 10308 3026 4 bl_50
port 185 nsew
rlabel metal1 s 10484 2874 10512 3026 4 bl_51
port 187 nsew
rlabel metal1 s 10688 2874 10716 3026 4 bl_52
port 189 nsew
rlabel metal1 s 10892 2874 10920 3026 4 bl_53
port 191 nsew
rlabel metal1 s 11096 2874 11124 3026 4 bl_54
port 193 nsew
rlabel metal1 s 11300 2874 11328 3026 4 bl_55
port 195 nsew
rlabel metal1 s 11504 2874 11532 3026 4 bl_56
port 197 nsew
rlabel metal1 s 11708 2874 11736 3026 4 bl_57
port 199 nsew
rlabel metal1 s 11912 2874 11940 3026 4 bl_58
port 201 nsew
rlabel metal1 s 12116 2874 12144 3026 4 bl_59
port 203 nsew
rlabel metal1 s 12320 2874 12348 3026 4 bl_60
port 205 nsew
rlabel metal1 s 12524 2874 12552 3026 4 bl_61
port 207 nsew
rlabel metal1 s 12728 2874 12756 3026 4 bl_62
port 209 nsew
rlabel metal1 s 12932 2874 12960 3026 4 bl_63
port 211 nsew
rlabel metal1 s 13136 2874 13164 3026 4 bl_64
port 213 nsew
rlabel metal1 s 13340 2874 13368 3026 4 bl_65
port 215 nsew
rlabel metal1 s 13544 2874 13572 3026 4 bl_66
port 217 nsew
rlabel metal1 s 13748 2874 13776 3026 4 bl_67
port 219 nsew
rlabel metal1 s 13952 2874 13980 3026 4 bl_68
port 221 nsew
rlabel metal1 s 14156 2874 14184 3026 4 bl_69
port 223 nsew
rlabel metal1 s 14360 2874 14388 3026 4 bl_70
port 225 nsew
rlabel metal1 s 14564 2874 14592 3026 4 bl_71
port 227 nsew
rlabel metal1 s 14768 2874 14796 3026 4 bl_72
port 229 nsew
rlabel metal1 s 14972 2874 15000 3026 4 bl_73
port 231 nsew
rlabel metal1 s 15176 2874 15204 3026 4 bl_74
port 233 nsew
rlabel metal1 s 15380 2874 15408 3026 4 bl_75
port 235 nsew
rlabel metal1 s 15584 2874 15612 3026 4 bl_76
port 237 nsew
rlabel metal1 s 15788 2874 15816 3026 4 bl_77
port 239 nsew
rlabel metal1 s 15992 2874 16020 3026 4 bl_78
port 241 nsew
rlabel metal1 s 16196 2874 16224 3026 4 bl_79
port 243 nsew
rlabel metal1 s 16400 2874 16428 3026 4 bl_80
port 245 nsew
rlabel metal1 s 16604 2874 16632 3026 4 bl_81
port 247 nsew
rlabel metal1 s 16808 2874 16836 3026 4 bl_82
port 249 nsew
rlabel metal1 s 17012 2874 17040 3026 4 bl_83
port 251 nsew
rlabel metal1 s 17216 2874 17244 3026 4 bl_84
port 253 nsew
rlabel metal1 s 17420 2874 17448 3026 4 bl_85
port 255 nsew
rlabel metal1 s 17624 2874 17652 3026 4 bl_86
port 257 nsew
rlabel metal1 s 17828 2874 17856 3026 4 bl_87
port 259 nsew
rlabel metal1 s 18032 2874 18060 3026 4 bl_88
port 261 nsew
rlabel metal1 s 18236 2874 18264 3026 4 bl_89
port 263 nsew
rlabel metal1 s 18440 2874 18468 3026 4 bl_90
port 265 nsew
rlabel metal1 s 18644 2874 18672 3026 4 bl_91
port 267 nsew
rlabel metal1 s 18848 2874 18876 3026 4 bl_92
port 269 nsew
rlabel metal1 s 19052 2874 19080 3026 4 bl_93
port 271 nsew
rlabel metal1 s 19256 2874 19284 3026 4 bl_94
port 273 nsew
rlabel metal1 s 19460 2874 19488 3026 4 bl_95
port 275 nsew
rlabel metal1 s 19664 2874 19692 3026 4 bl_96
port 277 nsew
rlabel metal1 s 19868 2874 19896 3026 4 bl_97
port 279 nsew
rlabel metal1 s 20072 2874 20100 3026 4 bl_98
port 281 nsew
rlabel metal1 s 20276 2874 20304 3026 4 bl_99
port 283 nsew
rlabel metal1 s 20480 2874 20508 3026 4 bl_100
port 285 nsew
rlabel metal1 s 20684 2874 20712 3026 4 bl_101
port 287 nsew
rlabel metal1 s 20888 2874 20916 3026 4 bl_102
port 289 nsew
rlabel metal1 s 21092 2874 21120 3026 4 bl_103
port 291 nsew
rlabel metal1 s 21296 2874 21324 3026 4 bl_104
port 293 nsew
rlabel metal1 s 21500 2874 21528 3026 4 bl_105
port 295 nsew
rlabel metal1 s 21704 2874 21732 3026 4 bl_106
port 297 nsew
rlabel metal1 s 21908 2874 21936 3026 4 bl_107
port 299 nsew
rlabel metal1 s 22112 2874 22140 3026 4 bl_108
port 301 nsew
rlabel metal1 s 22316 2874 22344 3026 4 bl_109
port 303 nsew
rlabel metal1 s 22520 2874 22548 3026 4 bl_110
port 305 nsew
rlabel metal1 s 22724 2874 22752 3026 4 bl_111
port 307 nsew
rlabel metal1 s 22928 2874 22956 3026 4 bl_112
port 309 nsew
rlabel metal1 s 23132 2874 23160 3026 4 bl_113
port 311 nsew
rlabel metal1 s 23336 2874 23364 3026 4 bl_114
port 313 nsew
rlabel metal1 s 23540 2874 23568 3026 4 bl_115
port 315 nsew
rlabel metal1 s 23744 2874 23772 3026 4 bl_116
port 317 nsew
rlabel metal1 s 23948 2874 23976 3026 4 bl_117
port 319 nsew
rlabel metal1 s 24152 2874 24180 3026 4 bl_118
port 321 nsew
rlabel metal1 s 24356 2874 24384 3026 4 bl_119
port 323 nsew
rlabel metal1 s 24560 2874 24588 3026 4 bl_120
port 325 nsew
rlabel metal1 s 24764 2874 24792 3026 4 bl_121
port 327 nsew
rlabel metal1 s 24968 2874 24996 3026 4 bl_122
port 329 nsew
rlabel metal1 s 25172 2874 25200 3026 4 bl_123
port 331 nsew
rlabel metal1 s 25376 2874 25404 3026 4 bl_124
port 333 nsew
rlabel metal1 s 25580 2874 25608 3026 4 bl_125
port 335 nsew
rlabel metal1 s 25784 2874 25812 3026 4 bl_126
port 337 nsew
rlabel metal1 s 25988 2874 26016 3026 4 bl_127
port 339 nsew
rlabel metal1 s 26192 2874 26220 3026 4 bl_128
port 341 nsew
rlabel metal1 s 26396 2874 26424 3026 4 bl_129
port 343 nsew
rlabel metal1 s 26600 2874 26628 3026 4 bl_130
port 345 nsew
rlabel metal1 s 26804 2874 26832 3026 4 bl_131
port 347 nsew
rlabel metal1 s 27008 2874 27036 3026 4 bl_132
port 349 nsew
rlabel metal1 s 27212 2874 27240 3026 4 bl_133
port 351 nsew
rlabel metal1 s 27416 2874 27444 3026 4 bl_134
port 353 nsew
rlabel metal1 s 27620 2874 27648 3026 4 bl_135
port 355 nsew
rlabel metal1 s 27824 2874 27852 3026 4 bl_136
port 357 nsew
rlabel metal1 s 28028 2874 28056 3026 4 bl_137
port 359 nsew
rlabel metal1 s 28232 2874 28260 3026 4 bl_138
port 361 nsew
rlabel metal1 s 28436 2874 28464 3026 4 bl_139
port 363 nsew
rlabel metal1 s 28640 2874 28668 3026 4 bl_140
port 365 nsew
rlabel metal1 s 28844 2874 28872 3026 4 bl_141
port 367 nsew
rlabel metal1 s 29048 2874 29076 3026 4 bl_142
port 369 nsew
rlabel metal1 s 29252 2874 29280 3026 4 bl_143
port 371 nsew
rlabel metal1 s 29456 2874 29484 3026 4 bl_144
port 373 nsew
rlabel metal1 s 29660 2874 29688 3026 4 bl_145
port 375 nsew
rlabel metal1 s 29864 2874 29892 3026 4 bl_146
port 377 nsew
rlabel metal1 s 30068 2874 30096 3026 4 bl_147
port 379 nsew
rlabel metal1 s 30272 2874 30300 3026 4 bl_148
port 381 nsew
rlabel metal1 s 30476 2874 30504 3026 4 bl_149
port 383 nsew
rlabel metal1 s 30680 2874 30708 3026 4 bl_150
port 385 nsew
rlabel metal1 s 30884 2874 30912 3026 4 bl_151
port 387 nsew
rlabel metal1 s 31088 2874 31116 3026 4 bl_152
port 389 nsew
rlabel metal1 s 31292 2874 31320 3026 4 bl_153
port 391 nsew
rlabel metal1 s 31496 2874 31524 3026 4 bl_154
port 393 nsew
rlabel metal1 s 31700 2874 31728 3026 4 bl_155
port 395 nsew
rlabel metal1 s 31904 2874 31932 3026 4 bl_156
port 397 nsew
rlabel metal1 s 32108 2874 32136 3026 4 bl_157
port 399 nsew
rlabel metal1 s 32312 2874 32340 3026 4 bl_158
port 401 nsew
rlabel metal1 s 32516 2874 32544 3026 4 bl_159
port 403 nsew
rlabel metal1 s 32720 2874 32748 3026 4 bl_160
port 405 nsew
rlabel metal1 s 32924 2874 32952 3026 4 bl_161
port 407 nsew
rlabel metal1 s 33128 2874 33156 3026 4 bl_162
port 409 nsew
rlabel metal1 s 33332 2874 33360 3026 4 bl_163
port 411 nsew
rlabel metal1 s 33536 2874 33564 3026 4 bl_164
port 413 nsew
rlabel metal1 s 33740 2874 33768 3026 4 bl_165
port 415 nsew
rlabel metal1 s 33944 2874 33972 3026 4 bl_166
port 417 nsew
rlabel metal1 s 34148 2874 34176 3026 4 bl_167
port 419 nsew
rlabel metal1 s 34352 2874 34380 3026 4 bl_168
port 421 nsew
rlabel metal1 s 34556 2874 34584 3026 4 bl_169
port 423 nsew
rlabel metal1 s 34760 2874 34788 3026 4 bl_170
port 425 nsew
rlabel metal1 s 34964 2874 34992 3026 4 bl_171
port 427 nsew
rlabel metal1 s 35168 2874 35196 3026 4 bl_172
port 429 nsew
rlabel metal1 s 35372 2874 35400 3026 4 bl_173
port 431 nsew
rlabel metal1 s 35576 2874 35604 3026 4 bl_174
port 433 nsew
rlabel metal1 s 35780 2874 35808 3026 4 bl_175
port 435 nsew
rlabel metal1 s 35984 2874 36012 3026 4 bl_176
port 437 nsew
rlabel metal1 s 36188 2874 36216 3026 4 bl_177
port 439 nsew
rlabel metal1 s 36392 2874 36420 3026 4 bl_178
port 441 nsew
rlabel metal1 s 36596 2874 36624 3026 4 bl_179
port 443 nsew
rlabel metal1 s 36800 2874 36828 3026 4 bl_180
port 445 nsew
rlabel metal1 s 37004 2874 37032 3026 4 bl_181
port 447 nsew
rlabel metal1 s 37208 2874 37236 3026 4 bl_182
port 449 nsew
rlabel metal1 s 37412 2874 37440 3026 4 bl_183
port 451 nsew
rlabel metal1 s 37616 2874 37644 3026 4 bl_184
port 453 nsew
rlabel metal1 s 37820 2874 37848 3026 4 bl_185
port 455 nsew
rlabel metal1 s 38024 2874 38052 3026 4 bl_186
port 457 nsew
rlabel metal1 s 38228 2874 38256 3026 4 bl_187
port 459 nsew
rlabel metal1 s 38432 2874 38460 3026 4 bl_188
port 461 nsew
rlabel metal1 s 38636 2874 38664 3026 4 bl_189
port 463 nsew
rlabel metal1 s 38840 2874 38868 3026 4 bl_190
port 465 nsew
rlabel metal1 s 39044 2874 39072 3026 4 bl_191
port 467 nsew
rlabel metal1 s 39248 2874 39276 3026 4 bl_192
port 469 nsew
rlabel metal1 s 39452 2874 39480 3026 4 bl_193
port 471 nsew
rlabel metal1 s 39656 2874 39684 3026 4 bl_194
port 473 nsew
rlabel metal1 s 39860 2874 39888 3026 4 bl_195
port 475 nsew
rlabel metal1 s 40064 2874 40092 3026 4 bl_196
port 477 nsew
rlabel metal1 s 40268 2874 40296 3026 4 bl_197
port 479 nsew
rlabel metal1 s 40472 2874 40500 3026 4 bl_198
port 481 nsew
rlabel metal1 s 40676 2874 40704 3026 4 bl_199
port 483 nsew
rlabel metal1 s 40880 2874 40908 3026 4 bl_200
port 485 nsew
rlabel metal1 s 41084 2874 41112 3026 4 bl_201
port 487 nsew
rlabel metal1 s 41288 2874 41316 3026 4 bl_202
port 489 nsew
rlabel metal1 s 41492 2874 41520 3026 4 bl_203
port 491 nsew
rlabel metal1 s 41696 2874 41724 3026 4 bl_204
port 493 nsew
rlabel metal1 s 41900 2874 41928 3026 4 bl_205
port 495 nsew
rlabel metal1 s 42104 2874 42132 3026 4 bl_206
port 497 nsew
rlabel metal1 s 42308 2874 42336 3026 4 bl_207
port 499 nsew
rlabel metal1 s 42512 2874 42540 3026 4 bl_208
port 501 nsew
rlabel metal1 s 42716 2874 42744 3026 4 bl_209
port 503 nsew
rlabel metal1 s 42920 2874 42948 3026 4 bl_210
port 505 nsew
rlabel metal1 s 43124 2874 43152 3026 4 bl_211
port 507 nsew
rlabel metal1 s 43328 2874 43356 3026 4 bl_212
port 509 nsew
rlabel metal1 s 43532 2874 43560 3026 4 bl_213
port 511 nsew
rlabel metal1 s 43736 2874 43764 3026 4 bl_214
port 513 nsew
rlabel metal1 s 43940 2874 43968 3026 4 bl_215
port 515 nsew
rlabel metal1 s 44144 2874 44172 3026 4 bl_216
port 517 nsew
rlabel metal1 s 44348 2874 44376 3026 4 bl_217
port 519 nsew
rlabel metal1 s 44552 2874 44580 3026 4 bl_218
port 521 nsew
rlabel metal1 s 44756 2874 44784 3026 4 bl_219
port 523 nsew
rlabel metal1 s 44960 2874 44988 3026 4 bl_220
port 525 nsew
rlabel metal1 s 45164 2874 45192 3026 4 bl_221
port 527 nsew
rlabel metal1 s 45368 2874 45396 3026 4 bl_222
port 529 nsew
rlabel metal1 s 45572 2874 45600 3026 4 bl_223
port 531 nsew
rlabel metal1 s 45776 2874 45804 3026 4 bl_224
port 533 nsew
rlabel metal1 s 45980 2874 46008 3026 4 bl_225
port 535 nsew
rlabel metal1 s 46184 2874 46212 3026 4 bl_226
port 537 nsew
rlabel metal1 s 46388 2874 46416 3026 4 bl_227
port 539 nsew
rlabel metal1 s 46592 2874 46620 3026 4 bl_228
port 541 nsew
rlabel metal1 s 46796 2874 46824 3026 4 bl_229
port 543 nsew
rlabel metal1 s 47000 2874 47028 3026 4 bl_230
port 545 nsew
rlabel metal1 s 47204 2874 47232 3026 4 bl_231
port 547 nsew
rlabel metal1 s 47408 2874 47436 3026 4 bl_232
port 549 nsew
rlabel metal1 s 47612 2874 47640 3026 4 bl_233
port 551 nsew
rlabel metal1 s 47816 2874 47844 3026 4 bl_234
port 553 nsew
rlabel metal1 s 48020 2874 48048 3026 4 bl_235
port 555 nsew
rlabel metal1 s 48224 2874 48252 3026 4 bl_236
port 557 nsew
rlabel metal1 s 48428 2874 48456 3026 4 bl_237
port 559 nsew
rlabel metal1 s 48632 2874 48660 3026 4 bl_238
port 561 nsew
rlabel metal1 s 48836 2874 48864 3026 4 bl_239
port 563 nsew
rlabel metal1 s 49040 2874 49068 3026 4 bl_240
port 565 nsew
rlabel metal1 s 49244 2874 49272 3026 4 bl_241
port 567 nsew
rlabel metal1 s 49448 2874 49476 3026 4 bl_242
port 569 nsew
rlabel metal1 s 49652 2874 49680 3026 4 bl_243
port 571 nsew
rlabel metal1 s 49856 2874 49884 3026 4 bl_244
port 573 nsew
rlabel metal1 s 50060 2874 50088 3026 4 bl_245
port 575 nsew
rlabel metal1 s 50264 2874 50292 3026 4 bl_246
port 577 nsew
rlabel metal1 s 50468 2874 50496 3026 4 bl_247
port 579 nsew
rlabel metal1 s 50672 2874 50700 3026 4 bl_248
port 581 nsew
rlabel metal1 s 50876 2874 50904 3026 4 bl_249
port 583 nsew
rlabel metal1 s 51080 2874 51108 3026 4 bl_250
port 585 nsew
rlabel metal1 s 51284 2874 51312 3026 4 bl_251
port 587 nsew
rlabel metal1 s 51488 2874 51516 3026 4 bl_252
port 589 nsew
rlabel metal1 s 51692 2874 51720 3026 4 bl_253
port 591 nsew
rlabel metal1 s 51896 2874 51924 3026 4 bl_254
port 593 nsew
rlabel metal1 s 52100 2874 52128 3026 4 bl_255
port 595 nsew
<< properties >>
string FIXED_BBOX 0 0 52224 2001
<< end >>
