magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1296 -1277 1674 3436
<< nwell >>
rect -36 1017 414 2176
<< pwell >>
rect 28 25 330 225
<< scnmos >>
rect 114 51 144 199
rect 214 51 244 199
<< scpmos >>
rect 114 1844 144 2068
rect 214 1844 244 2068
<< ndiff >>
rect 54 142 114 199
rect 54 108 62 142
rect 96 108 114 142
rect 54 51 114 108
rect 144 51 214 199
rect 244 142 304 199
rect 244 108 262 142
rect 296 108 304 142
rect 244 51 304 108
<< pdiff >>
rect 54 1973 114 2068
rect 54 1939 62 1973
rect 96 1939 114 1973
rect 54 1844 114 1939
rect 144 1973 214 2068
rect 144 1939 162 1973
rect 196 1939 214 1973
rect 144 1844 214 1939
rect 244 1973 304 2068
rect 244 1939 262 1973
rect 296 1939 304 1973
rect 244 1844 304 1939
<< ndiffc >>
rect 62 108 96 142
rect 262 108 296 142
<< pdiffc >>
rect 62 1939 96 1973
rect 162 1939 196 1973
rect 262 1939 296 1973
<< poly >>
rect 114 2068 144 2094
rect 214 2068 244 2094
rect 114 303 144 1844
rect 214 551 244 1844
rect 196 535 262 551
rect 196 501 212 535
rect 246 501 262 535
rect 196 485 262 501
rect 96 287 162 303
rect 96 253 112 287
rect 146 253 162 287
rect 96 237 162 253
rect 114 199 144 237
rect 214 199 244 485
rect 114 25 144 51
rect 214 25 244 51
<< polycont >>
rect 212 501 246 535
rect 112 253 146 287
<< locali >>
rect 0 2102 378 2136
rect 62 1973 96 2102
rect 62 1923 96 1939
rect 162 1973 196 1989
rect 162 1873 196 1939
rect 262 1973 296 2102
rect 262 1923 296 1939
rect 162 1839 364 1873
rect 212 535 246 551
rect 212 485 246 501
rect 112 287 146 303
rect 112 237 146 253
rect 330 243 364 1839
rect 262 209 364 243
rect 62 142 96 158
rect 62 17 96 108
rect 262 142 296 209
rect 262 92 296 108
rect 0 -17 378 17
<< labels >>
rlabel locali s 347 1856 347 1856 4 Z
port 1 nsew
rlabel locali s 189 0 189 0 4 gnd
port 2 nsew
rlabel locali s 189 2119 189 2119 4 vdd
port 3 nsew
rlabel locali s 129 270 129 270 4 A
port 4 nsew
rlabel locali s 229 518 229 518 4 B
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 378 1872
<< end >>
