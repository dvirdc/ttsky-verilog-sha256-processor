magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1299 -1216 7991 13973
<< locali >>
rect 3585 12339 3619 12355
rect 6679 12305 6713 12339
rect 3585 12289 3619 12305
rect 3585 12135 3619 12151
rect 6679 12101 6713 12135
rect 3585 12085 3619 12101
rect 3585 11827 3619 11843
rect 6679 11793 6713 11827
rect 3585 11777 3619 11793
rect 3585 11623 3619 11639
rect 6679 11589 6713 11623
rect 3585 11573 3619 11589
rect 3585 11419 3619 11435
rect 6679 11385 6713 11419
rect 3585 11369 3619 11385
rect 3585 11215 3619 11231
rect 6679 11181 6713 11215
rect 3585 11165 3619 11181
rect 3585 11011 3619 11027
rect 6679 10977 6713 11011
rect 3585 10961 3619 10977
rect 3585 10807 3619 10823
rect 6679 10773 6713 10807
rect 3585 10757 3619 10773
rect 3585 10603 3619 10619
rect 6679 10569 6713 10603
rect 3585 10553 3619 10569
rect 3585 10399 3619 10415
rect 6679 10365 6713 10399
rect 3585 10349 3619 10365
rect 3585 10091 3619 10107
rect 6679 10057 6713 10091
rect 3585 10041 3619 10057
rect 3585 9887 3619 9903
rect 6679 9853 6713 9887
rect 3585 9837 3619 9853
rect 3585 9683 3619 9699
rect 6679 9649 6713 9683
rect 3585 9633 3619 9649
rect 3585 9479 3619 9495
rect 6679 9445 6713 9479
rect 3585 9429 3619 9445
rect 3585 9275 3619 9291
rect 6679 9241 6713 9275
rect 3585 9225 3619 9241
rect 3585 9071 3619 9087
rect 6679 9037 6713 9071
rect 3585 9021 3619 9037
rect 3585 8867 3619 8883
rect 6679 8833 6713 8867
rect 3585 8817 3619 8833
rect 3585 8663 3619 8679
rect 6679 8629 6713 8663
rect 3585 8613 3619 8629
rect 3585 8355 3619 8371
rect 6679 8321 6713 8355
rect 3585 8305 3619 8321
rect 3585 8151 3619 8167
rect 6679 8117 6713 8151
rect 3585 8101 3619 8117
rect 3585 7947 3619 7963
rect 6679 7913 6713 7947
rect 3585 7897 3619 7913
rect 3585 7743 3619 7759
rect 6679 7709 6713 7743
rect 3585 7693 3619 7709
rect 3585 7539 3619 7555
rect 6679 7505 6713 7539
rect 3585 7489 3619 7505
rect 3585 7335 3619 7351
rect 6679 7301 6713 7335
rect 3585 7285 3619 7301
rect 3585 7131 3619 7147
rect 6679 7097 6713 7131
rect 3585 7081 3619 7097
rect 3585 6927 3619 6943
rect 6679 6893 6713 6927
rect 3585 6877 3619 6893
rect 3585 6619 3619 6635
rect 6679 6585 6713 6619
rect 3585 6569 3619 6585
rect 3585 6415 3619 6431
rect 6679 6381 6713 6415
rect 3585 6365 3619 6381
rect 3585 6211 3619 6227
rect 6679 6177 6713 6211
rect 3585 6161 3619 6177
rect 3585 6007 3619 6023
rect 6679 5973 6713 6007
rect 3585 5957 3619 5973
rect 3585 5803 3619 5819
rect 6679 5769 6713 5803
rect 3585 5753 3619 5769
rect 3585 5599 3619 5615
rect 6679 5565 6713 5599
rect 3585 5549 3619 5565
rect 3585 5395 3619 5411
rect 6679 5361 6713 5395
rect 3585 5345 3619 5361
rect 3585 5191 3619 5207
rect 6679 5157 6713 5191
rect 3585 5141 3619 5157
rect 3585 4883 3619 4899
rect 6679 4849 6713 4883
rect 3585 4833 3619 4849
rect 3585 4679 3619 4695
rect 6679 4645 6713 4679
rect 3585 4629 3619 4645
rect 3585 4475 3619 4491
rect 6679 4441 6713 4475
rect 3585 4425 3619 4441
rect 3585 4271 3619 4287
rect 6679 4237 6713 4271
rect 3585 4221 3619 4237
rect 3585 4067 3619 4083
rect 6679 4033 6713 4067
rect 3585 4017 3619 4033
rect 3585 3863 3619 3879
rect 6679 3829 6713 3863
rect 3585 3813 3619 3829
rect 3585 3659 3619 3675
rect 6679 3625 6713 3659
rect 3585 3609 3619 3625
rect 3585 3455 3619 3471
rect 6679 3421 6713 3455
rect 3585 3405 3619 3421
rect 321 60 387 94
rect 729 60 795 94
rect 1137 60 1203 94
rect 1545 60 1611 94
rect 1953 60 2019 94
rect 2361 60 2427 94
<< viali >>
rect 3585 12305 3619 12339
rect 3585 12101 3619 12135
rect 3585 11793 3619 11827
rect 3585 11589 3619 11623
rect 3585 11385 3619 11419
rect 3585 11181 3619 11215
rect 3585 10977 3619 11011
rect 3585 10773 3619 10807
rect 3585 10569 3619 10603
rect 3585 10365 3619 10399
rect 3585 10057 3619 10091
rect 3585 9853 3619 9887
rect 3585 9649 3619 9683
rect 3585 9445 3619 9479
rect 3585 9241 3619 9275
rect 3585 9037 3619 9071
rect 3585 8833 3619 8867
rect 3585 8629 3619 8663
rect 3585 8321 3619 8355
rect 3585 8117 3619 8151
rect 3585 7913 3619 7947
rect 3585 7709 3619 7743
rect 3585 7505 3619 7539
rect 3585 7301 3619 7335
rect 3585 7097 3619 7131
rect 3585 6893 3619 6927
rect 3585 6585 3619 6619
rect 3585 6381 3619 6415
rect 3585 6177 3619 6211
rect 3585 5973 3619 6007
rect 3585 5769 3619 5803
rect 3585 5565 3619 5599
rect 3585 5361 3619 5395
rect 3585 5157 3619 5191
rect 3585 4849 3619 4883
rect 3585 4645 3619 4679
rect 3585 4441 3619 4475
rect 3585 4237 3619 4271
rect 3585 4033 3619 4067
rect 3585 3829 3619 3863
rect 3585 3625 3619 3659
rect 3585 3421 3619 3455
<< metal1 >>
rect 3101 12685 3129 12713
rect 3709 12428 3737 12456
rect 4105 12428 4133 12456
rect 4715 12428 4743 12456
rect 5963 12428 5991 12456
rect 3573 12339 3631 12345
rect 3573 12336 3585 12339
rect 3483 12308 3585 12336
rect 3573 12305 3585 12308
rect 3619 12305 3631 12339
rect 3573 12299 3631 12305
rect 3573 12135 3631 12141
rect 3573 12132 3585 12135
rect 3483 12104 3585 12132
rect 3573 12101 3585 12104
rect 3619 12101 3631 12135
rect 3573 12095 3631 12101
rect 3573 11827 3631 11833
rect 3573 11824 3585 11827
rect 3483 11796 3585 11824
rect 3573 11793 3585 11796
rect 3619 11793 3631 11827
rect 3573 11787 3631 11793
rect 3573 11623 3631 11629
rect 3573 11620 3585 11623
rect 3483 11592 3585 11620
rect 3573 11589 3585 11592
rect 3619 11589 3631 11623
rect 3573 11583 3631 11589
rect 3573 11419 3631 11425
rect 3573 11416 3585 11419
rect 3483 11388 3585 11416
rect 3573 11385 3585 11388
rect 3619 11385 3631 11419
rect 3573 11379 3631 11385
rect 3573 11215 3631 11221
rect 3573 11212 3585 11215
rect 3483 11184 3585 11212
rect 3573 11181 3585 11184
rect 3619 11181 3631 11215
rect 3573 11175 3631 11181
rect 3573 11011 3631 11017
rect 3573 11008 3585 11011
rect 3483 10980 3585 11008
rect 3573 10977 3585 10980
rect 3619 10977 3631 11011
rect 3573 10971 3631 10977
rect 3573 10807 3631 10813
rect 3573 10804 3585 10807
rect 3483 10776 3585 10804
rect 3573 10773 3585 10776
rect 3619 10773 3631 10807
rect 3573 10767 3631 10773
rect 3573 10603 3631 10609
rect 3573 10600 3585 10603
rect 3483 10572 3585 10600
rect 3573 10569 3585 10572
rect 3619 10569 3631 10603
rect 3573 10563 3631 10569
rect 3573 10399 3631 10405
rect 3573 10396 3585 10399
rect 3483 10368 3585 10396
rect 3573 10365 3585 10368
rect 3619 10365 3631 10399
rect 3573 10359 3631 10365
rect 3573 10091 3631 10097
rect 3573 10088 3585 10091
rect 3483 10060 3585 10088
rect 3573 10057 3585 10060
rect 3619 10057 3631 10091
rect 3573 10051 3631 10057
rect 3573 9887 3631 9893
rect 3573 9884 3585 9887
rect 3483 9856 3585 9884
rect 3573 9853 3585 9856
rect 3619 9853 3631 9887
rect 3573 9847 3631 9853
rect 3573 9683 3631 9689
rect 3573 9680 3585 9683
rect 3483 9652 3585 9680
rect 3573 9649 3585 9652
rect 3619 9649 3631 9683
rect 3573 9643 3631 9649
rect 3573 9479 3631 9485
rect 3573 9476 3585 9479
rect 3483 9448 3585 9476
rect 3573 9445 3585 9448
rect 3619 9445 3631 9479
rect 3573 9439 3631 9445
rect 3573 9275 3631 9281
rect 3573 9272 3585 9275
rect 3483 9244 3585 9272
rect 3573 9241 3585 9244
rect 3619 9241 3631 9275
rect 3573 9235 3631 9241
rect 3573 9071 3631 9077
rect 3573 9068 3585 9071
rect 3483 9040 3585 9068
rect 3573 9037 3585 9040
rect 3619 9037 3631 9071
rect 3573 9031 3631 9037
rect 3573 8867 3631 8873
rect 3573 8864 3585 8867
rect 3483 8836 3585 8864
rect 3573 8833 3585 8836
rect 3619 8833 3631 8867
rect 3573 8827 3631 8833
rect 3573 8663 3631 8669
rect 3573 8660 3585 8663
rect 3483 8632 3585 8660
rect 3573 8629 3585 8632
rect 3619 8629 3631 8663
rect 3573 8623 3631 8629
rect 3573 8355 3631 8361
rect 3573 8352 3585 8355
rect 3483 8324 3585 8352
rect 3573 8321 3585 8324
rect 3619 8321 3631 8355
rect 3573 8315 3631 8321
rect 3573 8151 3631 8157
rect 3573 8148 3585 8151
rect 3483 8120 3585 8148
rect 3573 8117 3585 8120
rect 3619 8117 3631 8151
rect 3573 8111 3631 8117
rect 3573 7947 3631 7953
rect 3573 7944 3585 7947
rect 3483 7916 3585 7944
rect 3573 7913 3585 7916
rect 3619 7913 3631 7947
rect 3573 7907 3631 7913
rect 3573 7743 3631 7749
rect 3573 7740 3585 7743
rect 3483 7712 3585 7740
rect 3573 7709 3585 7712
rect 3619 7709 3631 7743
rect 3573 7703 3631 7709
rect 3573 7539 3631 7545
rect 3573 7536 3585 7539
rect 3483 7508 3585 7536
rect 3573 7505 3585 7508
rect 3619 7505 3631 7539
rect 3573 7499 3631 7505
rect 3573 7335 3631 7341
rect 3573 7332 3585 7335
rect 3483 7304 3585 7332
rect 3573 7301 3585 7304
rect 3619 7301 3631 7335
rect 3573 7295 3631 7301
rect 3573 7131 3631 7137
rect 3573 7128 3585 7131
rect 3483 7100 3585 7128
rect 3573 7097 3585 7100
rect 3619 7097 3631 7131
rect 3573 7091 3631 7097
rect 3573 6927 3631 6933
rect 3573 6924 3585 6927
rect 3483 6896 3585 6924
rect 3573 6893 3585 6896
rect 3619 6893 3631 6927
rect 3573 6887 3631 6893
rect 3573 6619 3631 6625
rect 3573 6616 3585 6619
rect 3483 6588 3585 6616
rect 3573 6585 3585 6588
rect 3619 6585 3631 6619
rect 3573 6579 3631 6585
rect 3573 6415 3631 6421
rect 3573 6412 3585 6415
rect 3483 6384 3585 6412
rect 3573 6381 3585 6384
rect 3619 6381 3631 6415
rect 3573 6375 3631 6381
rect 3573 6211 3631 6217
rect 3573 6208 3585 6211
rect 3483 6180 3585 6208
rect 3573 6177 3585 6180
rect 3619 6177 3631 6211
rect 3573 6171 3631 6177
rect 3573 6007 3631 6013
rect 3573 6004 3585 6007
rect 3483 5976 3585 6004
rect 3573 5973 3585 5976
rect 3619 5973 3631 6007
rect 3573 5967 3631 5973
rect 3573 5803 3631 5809
rect 3573 5800 3585 5803
rect 3483 5772 3585 5800
rect 3573 5769 3585 5772
rect 3619 5769 3631 5803
rect 3573 5763 3631 5769
rect 3573 5599 3631 5605
rect 3573 5596 3585 5599
rect 3483 5568 3585 5596
rect 3573 5565 3585 5568
rect 3619 5565 3631 5599
rect 3573 5559 3631 5565
rect 3573 5395 3631 5401
rect 3573 5392 3585 5395
rect 3483 5364 3585 5392
rect 3573 5361 3585 5364
rect 3619 5361 3631 5395
rect 3573 5355 3631 5361
rect 3573 5191 3631 5197
rect 3573 5188 3585 5191
rect 3483 5160 3585 5188
rect 3573 5157 3585 5160
rect 3619 5157 3631 5191
rect 3573 5151 3631 5157
rect 3573 4883 3631 4889
rect 3573 4880 3585 4883
rect 3483 4852 3585 4880
rect 3573 4849 3585 4852
rect 3619 4849 3631 4883
rect 3573 4843 3631 4849
rect 3573 4679 3631 4685
rect 3573 4676 3585 4679
rect 3483 4648 3585 4676
rect 3573 4645 3585 4648
rect 3619 4645 3631 4679
rect 3573 4639 3631 4645
rect 3573 4475 3631 4481
rect 3573 4472 3585 4475
rect 3483 4444 3585 4472
rect 3573 4441 3585 4444
rect 3619 4441 3631 4475
rect 3573 4435 3631 4441
rect 3573 4271 3631 4277
rect 3573 4268 3585 4271
rect 3483 4240 3585 4268
rect 3573 4237 3585 4240
rect 3619 4237 3631 4271
rect 3573 4231 3631 4237
rect 3573 4067 3631 4073
rect 3573 4064 3585 4067
rect 3483 4036 3585 4064
rect 3573 4033 3585 4036
rect 3619 4033 3631 4067
rect 3573 4027 3631 4033
rect 3573 3863 3631 3869
rect 3573 3860 3585 3863
rect 3483 3832 3585 3860
rect 3573 3829 3585 3832
rect 3619 3829 3631 3863
rect 3573 3823 3631 3829
rect 3573 3659 3631 3665
rect 3573 3656 3585 3659
rect 3483 3628 3585 3656
rect 3573 3625 3585 3628
rect 3619 3625 3631 3659
rect 3573 3619 3631 3625
rect 3573 3455 3631 3461
rect 3573 3452 3585 3455
rect 3483 3424 3585 3452
rect 3573 3421 3585 3424
rect 3619 3421 3631 3455
rect 3573 3415 3631 3421
rect 3709 3256 3737 3284
rect 4105 3256 4133 3284
rect 4715 3256 4743 3284
rect 5963 3256 5991 3284
rect 298 3199 304 3251
rect 356 3199 362 3251
rect 502 3199 508 3251
rect 560 3199 566 3251
rect 706 3199 712 3251
rect 764 3199 770 3251
rect 910 3199 916 3251
rect 968 3199 974 3251
rect 1114 3199 1120 3251
rect 1172 3199 1178 3251
rect 1318 3199 1324 3251
rect 1376 3199 1382 3251
rect 1522 3199 1528 3251
rect 1580 3199 1586 3251
rect 1726 3199 1732 3251
rect 1784 3199 1790 3251
rect 1930 3199 1936 3251
rect 1988 3199 1994 3251
rect 2134 3199 2140 3251
rect 2192 3199 2198 3251
rect 2338 3199 2344 3251
rect 2396 3199 2402 3251
rect 2542 3199 2548 3251
rect 2600 3199 2606 3251
rect 316 3138 344 3199
rect 298 3086 304 3138
rect 356 3086 362 3138
rect 438 3086 444 3138
rect 496 3126 502 3138
rect 520 3126 548 3199
rect 724 3138 752 3199
rect 496 3098 548 3126
rect 496 3086 502 3098
rect 706 3086 712 3138
rect 764 3086 770 3138
rect 846 3086 852 3138
rect 904 3126 910 3138
rect 928 3126 956 3199
rect 1132 3138 1160 3199
rect 904 3098 956 3126
rect 904 3086 910 3098
rect 1114 3086 1120 3138
rect 1172 3086 1178 3138
rect 1254 3086 1260 3138
rect 1312 3126 1318 3138
rect 1336 3126 1364 3199
rect 1540 3138 1568 3199
rect 1312 3098 1364 3126
rect 1312 3086 1318 3098
rect 1522 3086 1528 3138
rect 1580 3086 1586 3138
rect 1662 3086 1668 3138
rect 1720 3126 1726 3138
rect 1744 3126 1772 3199
rect 1948 3138 1976 3199
rect 1720 3098 1772 3126
rect 1720 3086 1726 3098
rect 1930 3086 1936 3138
rect 1988 3086 1994 3138
rect 2070 3086 2076 3138
rect 2128 3126 2134 3138
rect 2152 3126 2180 3199
rect 2356 3138 2384 3199
rect 2128 3098 2180 3126
rect 2128 3086 2134 3098
rect 2338 3086 2344 3138
rect 2396 3086 2402 3138
rect 2478 3086 2484 3138
rect 2536 3126 2542 3138
rect 2560 3126 2588 3199
rect 2536 3098 2588 3126
rect 2536 3086 2542 3098
rect 127 2833 155 2861
rect 2575 2408 2603 2436
rect 127 2160 2575 2188
rect 127 1881 155 1909
rect 2575 1456 2603 1484
rect 127 844 155 872
rect 2575 222 2603 250
<< via1 >>
rect 304 3199 356 3251
rect 508 3199 560 3251
rect 712 3199 764 3251
rect 916 3199 968 3251
rect 1120 3199 1172 3251
rect 1324 3199 1376 3251
rect 1528 3199 1580 3251
rect 1732 3199 1784 3251
rect 1936 3199 1988 3251
rect 2140 3199 2192 3251
rect 2344 3199 2396 3251
rect 2548 3199 2600 3251
rect 304 3086 356 3138
rect 444 3086 496 3138
rect 712 3086 764 3138
rect 852 3086 904 3138
rect 1120 3086 1172 3138
rect 1260 3086 1312 3138
rect 1528 3086 1580 3138
rect 1668 3086 1720 3138
rect 1936 3086 1988 3138
rect 2076 3086 2128 3138
rect 2344 3086 2396 3138
rect 2484 3086 2536 3138
<< metal2 >>
rect 304 3251 356 3257
rect 304 3193 356 3199
rect 508 3251 560 3257
rect 508 3193 560 3199
rect 712 3251 764 3257
rect 712 3193 764 3199
rect 916 3251 968 3257
rect 916 3193 968 3199
rect 1120 3251 1172 3257
rect 1120 3193 1172 3199
rect 1324 3251 1376 3257
rect 1324 3193 1376 3199
rect 1528 3251 1580 3257
rect 1528 3193 1580 3199
rect 1732 3251 1784 3257
rect 1732 3193 1784 3199
rect 1936 3251 1988 3257
rect 1936 3193 1988 3199
rect 2140 3251 2192 3257
rect 2140 3193 2192 3199
rect 2344 3251 2396 3257
rect 2344 3193 2396 3199
rect 2548 3251 2600 3257
rect 3101 3253 3129 3281
rect 3465 3204 3529 3232
rect 2548 3193 2600 3199
rect 304 3138 356 3144
rect 304 3080 356 3086
rect 444 3138 496 3144
rect 444 3080 496 3086
rect 712 3138 764 3144
rect 712 3080 764 3086
rect 852 3138 904 3144
rect 852 3080 904 3086
rect 1120 3138 1172 3144
rect 1120 3080 1172 3086
rect 1260 3138 1312 3144
rect 1260 3080 1312 3086
rect 1528 3138 1580 3144
rect 1528 3080 1580 3086
rect 1668 3138 1720 3144
rect 1668 3080 1720 3086
rect 1936 3138 1988 3144
rect 1936 3080 1988 3086
rect 2076 3138 2128 3144
rect 2076 3080 2128 3086
rect 2344 3138 2396 3144
rect 2344 3080 2396 3086
rect 2484 3138 2536 3144
rect 2484 3080 2536 3086
<< metal3 >>
rect -31 12415 29 12475
rect 2459 12415 2519 12475
rect -31 11903 29 11963
rect 2459 11903 2519 11963
rect -31 10167 29 10227
rect 2459 10167 2519 10227
rect -31 8431 29 8491
rect 2459 8431 2519 8491
rect -31 6695 29 6755
rect 2459 6695 2519 6755
rect -31 4959 29 5019
rect 2459 4959 2519 5019
rect -31 3223 29 3283
rect 2459 3223 2519 3283
use sky130_rom_krom_rom_address_control_array  sky130_rom_krom_rom_address_control_array_0
timestamp 1581321264
transform 1 0 127 0 1 0
box -48 44 2543 3128
use sky130_rom_krom_rom_row_decode_array  sky130_rom_krom_rom_row_decode_array_0
timestamp 1581321264
transform 0 -1 3497 1 0 3192
box -6 -84 9521 3536
use sky130_rom_krom_rom_row_decode_wordline_buffer  sky130_rom_krom_rom_row_decode_wordline_buffer_0
timestamp 1581321264
transform 1 0 3525 0 1 3250
box 44 -50 3206 9287
<< labels >>
rlabel metal1 s 127 2160 2575 2188 4 clk
port 3 nsew
rlabel locali s 6696 3438 6696 3438 4 wl_0
port 4 nsew
rlabel locali s 6696 3642 6696 3642 4 wl_1
port 5 nsew
rlabel locali s 6696 3846 6696 3846 4 wl_2
port 6 nsew
rlabel locali s 6696 4050 6696 4050 4 wl_3
port 7 nsew
rlabel locali s 6696 4254 6696 4254 4 wl_4
port 8 nsew
rlabel locali s 6696 4458 6696 4458 4 wl_5
port 9 nsew
rlabel locali s 6696 4662 6696 4662 4 wl_6
port 10 nsew
rlabel locali s 6696 4866 6696 4866 4 wl_7
port 11 nsew
rlabel locali s 6696 5174 6696 5174 4 wl_8
port 12 nsew
rlabel locali s 6696 5378 6696 5378 4 wl_9
port 13 nsew
rlabel locali s 6696 5582 6696 5582 4 wl_10
port 14 nsew
rlabel locali s 6696 5786 6696 5786 4 wl_11
port 15 nsew
rlabel locali s 6696 5990 6696 5990 4 wl_12
port 16 nsew
rlabel locali s 6696 6194 6696 6194 4 wl_13
port 17 nsew
rlabel locali s 6696 6398 6696 6398 4 wl_14
port 18 nsew
rlabel locali s 6696 6602 6696 6602 4 wl_15
port 19 nsew
rlabel locali s 6696 6910 6696 6910 4 wl_16
port 20 nsew
rlabel locali s 6696 7114 6696 7114 4 wl_17
port 21 nsew
rlabel locali s 6696 7318 6696 7318 4 wl_18
port 22 nsew
rlabel locali s 6696 7522 6696 7522 4 wl_19
port 23 nsew
rlabel locali s 6696 7726 6696 7726 4 wl_20
port 24 nsew
rlabel locali s 6696 7930 6696 7930 4 wl_21
port 25 nsew
rlabel locali s 6696 8134 6696 8134 4 wl_22
port 26 nsew
rlabel locali s 6696 8338 6696 8338 4 wl_23
port 27 nsew
rlabel locali s 6696 8646 6696 8646 4 wl_24
port 28 nsew
rlabel locali s 6696 8850 6696 8850 4 wl_25
port 29 nsew
rlabel locali s 6696 9054 6696 9054 4 wl_26
port 30 nsew
rlabel locali s 6696 9258 6696 9258 4 wl_27
port 31 nsew
rlabel locali s 6696 9462 6696 9462 4 wl_28
port 32 nsew
rlabel locali s 6696 9666 6696 9666 4 wl_29
port 33 nsew
rlabel locali s 6696 9870 6696 9870 4 wl_30
port 34 nsew
rlabel locali s 6696 10074 6696 10074 4 wl_31
port 35 nsew
rlabel locali s 6696 10382 6696 10382 4 wl_32
port 36 nsew
rlabel locali s 6696 10586 6696 10586 4 wl_33
port 37 nsew
rlabel locali s 6696 10790 6696 10790 4 wl_34
port 38 nsew
rlabel locali s 6696 10994 6696 10994 4 wl_35
port 39 nsew
rlabel locali s 6696 11198 6696 11198 4 wl_36
port 40 nsew
rlabel locali s 6696 11402 6696 11402 4 wl_37
port 41 nsew
rlabel locali s 6696 11606 6696 11606 4 wl_38
port 42 nsew
rlabel locali s 6696 11810 6696 11810 4 wl_39
port 43 nsew
rlabel locali s 6696 12118 6696 12118 4 wl_40
port 44 nsew
rlabel locali s 6696 12322 6696 12322 4 wl_41
port 45 nsew
rlabel metal2 s 3101 3253 3129 3281 4 precharge
port 47 nsew
rlabel metal1 s 3101 12685 3129 12713 4 precharge_r
port 49 nsew
rlabel locali s 354 77 354 77 4 A0
port 50 nsew
rlabel locali s 762 77 762 77 4 A1
port 51 nsew
rlabel locali s 1170 77 1170 77 4 A2
port 52 nsew
rlabel locali s 1578 77 1578 77 4 A3
port 53 nsew
rlabel locali s 1986 77 1986 77 4 A4
port 54 nsew
rlabel locali s 2394 77 2394 77 4 A5
port 55 nsew
rlabel metal2 s 3465 3204 3529 3232 4 vdd
port 57 nsew
rlabel metal1 s 127 2833 155 2861 4 vdd
port 57 nsew
rlabel metal1 s 5963 3256 5991 3284 4 vdd
port 57 nsew
rlabel metal1 s 5963 12428 5991 12456 4 vdd
port 57 nsew
rlabel metal1 s 4105 3256 4133 3284 4 vdd
port 57 nsew
rlabel metal1 s 127 1881 155 1909 4 vdd
port 57 nsew
rlabel metal1 s 4105 12428 4133 12456 4 vdd
port 57 nsew
rlabel metal1 s 127 844 155 872 4 vdd
port 57 nsew
rlabel metal3 s -31 8431 29 8491 4 gnd
port 59 nsew
rlabel metal3 s -31 4959 29 5019 4 gnd
port 59 nsew
rlabel metal3 s -31 12415 29 12475 4 gnd
port 59 nsew
rlabel metal3 s 2459 8431 2519 8491 4 gnd
port 59 nsew
rlabel metal1 s 3709 12428 3737 12456 4 gnd
port 59 nsew
rlabel metal1 s 2575 1456 2603 1484 4 gnd
port 59 nsew
rlabel metal1 s 2575 222 2603 250 4 gnd
port 59 nsew
rlabel metal3 s 2459 11903 2519 11963 4 gnd
port 59 nsew
rlabel metal3 s 2459 10167 2519 10227 4 gnd
port 59 nsew
rlabel metal3 s 2459 4959 2519 5019 4 gnd
port 59 nsew
rlabel metal1 s 4715 3256 4743 3284 4 gnd
port 59 nsew
rlabel metal1 s 4715 12428 4743 12456 4 gnd
port 59 nsew
rlabel metal3 s 2459 12415 2519 12475 4 gnd
port 59 nsew
rlabel metal1 s 2575 2408 2603 2436 4 gnd
port 59 nsew
rlabel metal1 s 3709 3256 3737 3284 4 gnd
port 59 nsew
rlabel metal3 s -31 11903 29 11963 4 gnd
port 59 nsew
rlabel metal3 s -31 6695 29 6755 4 gnd
port 59 nsew
rlabel metal3 s 2459 3223 2519 3283 4 gnd
port 59 nsew
rlabel metal3 s 2459 6695 2519 6755 4 gnd
port 59 nsew
rlabel metal3 s -31 3223 29 3283 4 gnd
port 59 nsew
rlabel metal3 s -31 10167 29 10227 4 gnd
port 59 nsew
<< properties >>
string FIXED_BBOX -31 0 6713 12713
<< end >>
