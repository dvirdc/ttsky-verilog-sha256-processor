magic
tech sky130A
magscale 1 2
timestamp 1581321264
<< checkpaint >>
rect -1216 -1310 3060 6283
<< nwell >>
rect 1162 4570 1330 4738
rect 1162 4262 1330 4430
rect 1162 3954 1330 4122
rect 1162 3646 1330 3814
rect 1162 3338 1330 3506
rect 1162 3030 1330 3198
rect 1162 2722 1330 2890
rect 1162 2414 1330 2582
rect 1162 2106 1330 2274
rect 1162 1798 1330 1966
rect 1162 1490 1330 1658
rect 1162 1182 1330 1350
rect 1162 874 1330 1042
rect 1162 566 1330 734
rect 1162 258 1330 426
rect 1162 -50 1330 118
<< pwell >>
rect 263 4603 397 4705
rect 263 4295 397 4397
rect 263 3987 397 4089
rect 263 3679 397 3781
rect 263 3371 397 3473
rect 263 3063 397 3165
rect 263 2755 397 2857
rect 263 2447 397 2549
rect 263 2139 397 2241
rect 263 1831 397 1933
rect 263 1523 397 1625
rect 263 1215 397 1317
rect 263 907 397 1009
rect 263 599 397 701
rect 263 291 397 393
rect 263 -17 397 85
<< psubdiff >>
rect 289 4671 371 4679
rect 289 4637 313 4671
rect 347 4637 371 4671
rect 289 4629 371 4637
rect 289 4363 371 4371
rect 289 4329 313 4363
rect 347 4329 371 4363
rect 289 4321 371 4329
rect 289 4055 371 4063
rect 289 4021 313 4055
rect 347 4021 371 4055
rect 289 4013 371 4021
rect 289 3747 371 3755
rect 289 3713 313 3747
rect 347 3713 371 3747
rect 289 3705 371 3713
rect 289 3439 371 3447
rect 289 3405 313 3439
rect 347 3405 371 3439
rect 289 3397 371 3405
rect 289 3131 371 3139
rect 289 3097 313 3131
rect 347 3097 371 3131
rect 289 3089 371 3097
rect 289 2823 371 2831
rect 289 2789 313 2823
rect 347 2789 371 2823
rect 289 2781 371 2789
rect 289 2515 371 2523
rect 289 2481 313 2515
rect 347 2481 371 2515
rect 289 2473 371 2481
rect 289 2207 371 2215
rect 289 2173 313 2207
rect 347 2173 371 2207
rect 289 2165 371 2173
rect 289 1899 371 1907
rect 289 1865 313 1899
rect 347 1865 371 1899
rect 289 1857 371 1865
rect 289 1591 371 1599
rect 289 1557 313 1591
rect 347 1557 371 1591
rect 289 1549 371 1557
rect 289 1283 371 1291
rect 289 1249 313 1283
rect 347 1249 371 1283
rect 289 1241 371 1249
rect 289 975 371 983
rect 289 941 313 975
rect 347 941 371 975
rect 289 933 371 941
rect 289 667 371 675
rect 289 633 313 667
rect 347 633 371 667
rect 289 625 371 633
rect 289 359 371 367
rect 289 325 313 359
rect 347 325 371 359
rect 289 317 371 325
rect 289 51 371 59
rect 289 17 313 51
rect 347 17 371 51
rect 289 9 371 17
<< nsubdiff >>
rect 1205 4671 1287 4679
rect 1205 4637 1229 4671
rect 1263 4637 1287 4671
rect 1205 4629 1287 4637
rect 1205 4363 1287 4371
rect 1205 4329 1229 4363
rect 1263 4329 1287 4363
rect 1205 4321 1287 4329
rect 1205 4055 1287 4063
rect 1205 4021 1229 4055
rect 1263 4021 1287 4055
rect 1205 4013 1287 4021
rect 1205 3747 1287 3755
rect 1205 3713 1229 3747
rect 1263 3713 1287 3747
rect 1205 3705 1287 3713
rect 1205 3439 1287 3447
rect 1205 3405 1229 3439
rect 1263 3405 1287 3439
rect 1205 3397 1287 3405
rect 1205 3131 1287 3139
rect 1205 3097 1229 3131
rect 1263 3097 1287 3131
rect 1205 3089 1287 3097
rect 1205 2823 1287 2831
rect 1205 2789 1229 2823
rect 1263 2789 1287 2823
rect 1205 2781 1287 2789
rect 1205 2515 1287 2523
rect 1205 2481 1229 2515
rect 1263 2481 1287 2515
rect 1205 2473 1287 2481
rect 1205 2207 1287 2215
rect 1205 2173 1229 2207
rect 1263 2173 1287 2207
rect 1205 2165 1287 2173
rect 1205 1899 1287 1907
rect 1205 1865 1229 1899
rect 1263 1865 1287 1899
rect 1205 1857 1287 1865
rect 1205 1591 1287 1599
rect 1205 1557 1229 1591
rect 1263 1557 1287 1591
rect 1205 1549 1287 1557
rect 1205 1283 1287 1291
rect 1205 1249 1229 1283
rect 1263 1249 1287 1283
rect 1205 1241 1287 1249
rect 1205 975 1287 983
rect 1205 941 1229 975
rect 1263 941 1287 975
rect 1205 933 1287 941
rect 1205 667 1287 675
rect 1205 633 1229 667
rect 1263 633 1287 667
rect 1205 625 1287 633
rect 1205 359 1287 367
rect 1205 325 1229 359
rect 1263 325 1287 359
rect 1205 317 1287 325
rect 1205 51 1287 59
rect 1205 17 1229 51
rect 1263 17 1287 51
rect 1205 9 1287 17
<< psubdiffcont >>
rect 313 4637 347 4671
rect 313 4329 347 4363
rect 313 4021 347 4055
rect 313 3713 347 3747
rect 313 3405 347 3439
rect 313 3097 347 3131
rect 313 2789 347 2823
rect 313 2481 347 2515
rect 313 2173 347 2207
rect 313 1865 347 1899
rect 313 1557 347 1591
rect 313 1249 347 1283
rect 313 941 347 975
rect 313 633 347 667
rect 313 325 347 359
rect 313 17 347 51
<< nsubdiffcont >>
rect 1229 4637 1263 4671
rect 1229 4329 1263 4363
rect 1229 4021 1263 4055
rect 1229 3713 1263 3747
rect 1229 3405 1263 3439
rect 1229 3097 1263 3131
rect 1229 2789 1263 2823
rect 1229 2481 1263 2515
rect 1229 2173 1263 2207
rect 1229 1865 1263 1899
rect 1229 1557 1263 1591
rect 1229 1249 1263 1283
rect 1229 941 1263 975
rect 1229 633 1263 667
rect 1229 325 1263 359
rect 1229 17 1263 51
<< locali >>
rect 60 4775 94 4841
rect 1748 4758 1782 4825
rect 297 4637 313 4671
rect 347 4637 363 4671
rect 1213 4637 1229 4671
rect 1263 4637 1279 4671
rect 60 4467 94 4533
rect 1748 4450 1782 4517
rect 297 4329 313 4363
rect 347 4329 363 4363
rect 1213 4329 1229 4363
rect 1263 4329 1279 4363
rect 60 4159 94 4225
rect 1748 4142 1782 4209
rect 297 4021 313 4055
rect 347 4021 363 4055
rect 1213 4021 1229 4055
rect 1263 4021 1279 4055
rect 60 3851 94 3917
rect 1748 3834 1782 3901
rect 297 3713 313 3747
rect 347 3713 363 3747
rect 1213 3713 1229 3747
rect 1263 3713 1279 3747
rect 60 3543 94 3609
rect 1748 3526 1782 3593
rect 297 3405 313 3439
rect 347 3405 363 3439
rect 1213 3405 1229 3439
rect 1263 3405 1279 3439
rect 60 3235 94 3301
rect 1748 3218 1782 3285
rect 297 3097 313 3131
rect 347 3097 363 3131
rect 1213 3097 1229 3131
rect 1263 3097 1279 3131
rect 60 2927 94 2993
rect 1748 2910 1782 2977
rect 297 2789 313 2823
rect 347 2789 363 2823
rect 1213 2789 1229 2823
rect 1263 2789 1279 2823
rect 60 2619 94 2685
rect 1748 2602 1782 2669
rect 297 2481 313 2515
rect 347 2481 363 2515
rect 1213 2481 1229 2515
rect 1263 2481 1279 2515
rect 60 2311 94 2377
rect 1748 2294 1782 2361
rect 297 2173 313 2207
rect 347 2173 363 2207
rect 1213 2173 1229 2207
rect 1263 2173 1279 2207
rect 60 2003 94 2069
rect 1748 1986 1782 2053
rect 297 1865 313 1899
rect 347 1865 363 1899
rect 1213 1865 1229 1899
rect 1263 1865 1279 1899
rect 60 1695 94 1761
rect 1748 1678 1782 1745
rect 297 1557 313 1591
rect 347 1557 363 1591
rect 1213 1557 1229 1591
rect 1263 1557 1279 1591
rect 60 1387 94 1453
rect 1748 1370 1782 1437
rect 297 1249 313 1283
rect 347 1249 363 1283
rect 1213 1249 1229 1283
rect 1263 1249 1279 1283
rect 60 1079 94 1145
rect 1748 1062 1782 1129
rect 297 941 313 975
rect 347 941 363 975
rect 1213 941 1229 975
rect 1263 941 1279 975
rect 60 771 94 837
rect 1748 754 1782 821
rect 297 633 313 667
rect 347 633 363 667
rect 1213 633 1229 667
rect 1263 633 1279 667
rect 60 463 94 529
rect 1748 446 1782 513
rect 297 325 313 359
rect 347 325 363 359
rect 1213 325 1229 359
rect 1263 325 1279 359
rect 60 155 94 221
rect 1748 138 1782 205
rect 297 17 313 51
rect 347 17 363 51
rect 1213 17 1229 51
rect 1263 17 1279 51
<< viali >>
rect 313 4637 347 4671
rect 1229 4637 1263 4671
rect 313 4329 347 4363
rect 1229 4329 1263 4363
rect 313 4021 347 4055
rect 1229 4021 1263 4055
rect 313 3713 347 3747
rect 1229 3713 1263 3747
rect 313 3405 347 3439
rect 1229 3405 1263 3439
rect 313 3097 347 3131
rect 1229 3097 1263 3131
rect 313 2789 347 2823
rect 1229 2789 1263 2823
rect 313 2481 347 2515
rect 1229 2481 1263 2515
rect 313 2173 347 2207
rect 1229 2173 1263 2207
rect 313 1865 347 1899
rect 1229 1865 1263 1899
rect 313 1557 347 1591
rect 1229 1557 1263 1591
rect 313 1249 347 1283
rect 1229 1249 1263 1283
rect 313 941 347 975
rect 1229 941 1263 975
rect 313 633 347 667
rect 1229 633 1263 667
rect 313 325 347 359
rect 1229 325 1263 359
rect 313 17 347 51
rect 1229 17 1263 51
<< metal1 >>
rect 316 4683 344 4942
rect 1232 4683 1260 4942
rect 307 4671 353 4683
rect 307 4637 313 4671
rect 347 4637 353 4671
rect 307 4625 353 4637
rect 1223 4671 1269 4683
rect 1223 4637 1229 4671
rect 1263 4637 1269 4671
rect 1223 4625 1269 4637
rect 316 4375 344 4625
rect 1232 4375 1260 4625
rect 307 4363 353 4375
rect 307 4329 313 4363
rect 347 4329 353 4363
rect 307 4317 353 4329
rect 1223 4363 1269 4375
rect 1223 4329 1229 4363
rect 1263 4329 1269 4363
rect 1223 4317 1269 4329
rect 316 4067 344 4317
rect 1232 4067 1260 4317
rect 307 4055 353 4067
rect 307 4021 313 4055
rect 347 4021 353 4055
rect 307 4009 353 4021
rect 1223 4055 1269 4067
rect 1223 4021 1229 4055
rect 1263 4021 1269 4055
rect 1223 4009 1269 4021
rect 316 3759 344 4009
rect 1232 3759 1260 4009
rect 307 3747 353 3759
rect 307 3713 313 3747
rect 347 3713 353 3747
rect 307 3701 353 3713
rect 1223 3747 1269 3759
rect 1223 3713 1229 3747
rect 1263 3713 1269 3747
rect 1223 3701 1269 3713
rect 316 3451 344 3701
rect 1232 3451 1260 3701
rect 307 3439 353 3451
rect 307 3405 313 3439
rect 347 3405 353 3439
rect 307 3393 353 3405
rect 1223 3439 1269 3451
rect 1223 3405 1229 3439
rect 1263 3405 1269 3439
rect 1223 3393 1269 3405
rect 316 3143 344 3393
rect 1232 3143 1260 3393
rect 307 3131 353 3143
rect 307 3097 313 3131
rect 347 3097 353 3131
rect 307 3085 353 3097
rect 1223 3131 1269 3143
rect 1223 3097 1229 3131
rect 1263 3097 1269 3131
rect 1223 3085 1269 3097
rect 316 2835 344 3085
rect 1232 2835 1260 3085
rect 307 2823 353 2835
rect 307 2789 313 2823
rect 347 2789 353 2823
rect 307 2777 353 2789
rect 1223 2823 1269 2835
rect 1223 2789 1229 2823
rect 1263 2789 1269 2823
rect 1223 2777 1269 2789
rect 316 2527 344 2777
rect 1232 2527 1260 2777
rect 307 2515 353 2527
rect 307 2481 313 2515
rect 347 2481 353 2515
rect 307 2469 353 2481
rect 1223 2515 1269 2527
rect 1223 2481 1229 2515
rect 1263 2481 1269 2515
rect 1223 2469 1269 2481
rect 316 2219 344 2469
rect 1232 2219 1260 2469
rect 307 2207 353 2219
rect 307 2173 313 2207
rect 347 2173 353 2207
rect 307 2161 353 2173
rect 1223 2207 1269 2219
rect 1223 2173 1229 2207
rect 1263 2173 1269 2207
rect 1223 2161 1269 2173
rect 316 1911 344 2161
rect 1232 1911 1260 2161
rect 307 1899 353 1911
rect 307 1865 313 1899
rect 347 1865 353 1899
rect 307 1853 353 1865
rect 1223 1899 1269 1911
rect 1223 1865 1229 1899
rect 1263 1865 1269 1899
rect 1223 1853 1269 1865
rect 316 1603 344 1853
rect 1232 1603 1260 1853
rect 307 1591 353 1603
rect 307 1557 313 1591
rect 347 1557 353 1591
rect 307 1545 353 1557
rect 1223 1591 1269 1603
rect 1223 1557 1229 1591
rect 1263 1557 1269 1591
rect 1223 1545 1269 1557
rect 316 1295 344 1545
rect 1232 1295 1260 1545
rect 307 1283 353 1295
rect 307 1249 313 1283
rect 347 1249 353 1283
rect 307 1237 353 1249
rect 1223 1283 1269 1295
rect 1223 1249 1229 1283
rect 1263 1249 1269 1283
rect 1223 1237 1269 1249
rect 316 987 344 1237
rect 1232 987 1260 1237
rect 307 975 353 987
rect 307 941 313 975
rect 347 941 353 975
rect 307 929 353 941
rect 1223 975 1269 987
rect 1223 941 1229 975
rect 1263 941 1269 975
rect 1223 929 1269 941
rect 316 679 344 929
rect 1232 679 1260 929
rect 307 667 353 679
rect 307 633 313 667
rect 347 633 353 667
rect 307 621 353 633
rect 1223 667 1269 679
rect 1223 633 1229 667
rect 1263 633 1269 667
rect 1223 621 1269 633
rect 316 371 344 621
rect 1232 371 1260 621
rect 307 359 353 371
rect 307 325 313 359
rect 347 325 353 359
rect 307 313 353 325
rect 1223 359 1269 371
rect 1223 325 1229 359
rect 1263 325 1269 359
rect 1223 313 1269 325
rect 316 63 344 313
rect 1232 63 1260 313
rect 307 51 353 63
rect 307 17 313 51
rect 347 17 353 51
rect 307 5 353 17
rect 1223 51 1269 63
rect 1223 17 1229 51
rect 1263 17 1269 51
rect 1223 5 1269 17
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_0
timestamp 1581321264
transform 1 0 0 0 1 4724
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_1
timestamp 1581321264
transform 1 0 0 0 1 4416
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_2
timestamp 1581321264
transform 1 0 0 0 1 4108
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_3
timestamp 1581321264
transform 1 0 0 0 1 3800
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_4
timestamp 1581321264
transform 1 0 0 0 1 3492
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_5
timestamp 1581321264
transform 1 0 0 0 1 3184
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_6
timestamp 1581321264
transform 1 0 0 0 1 2876
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_7
timestamp 1581321264
transform 1 0 0 0 1 2568
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_8
timestamp 1581321264
transform 1 0 0 0 1 2260
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_9
timestamp 1581321264
transform 1 0 0 0 1 1952
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_10
timestamp 1581321264
transform 1 0 0 0 1 1644
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_11
timestamp 1581321264
transform 1 0 0 0 1 1336
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_12
timestamp 1581321264
transform 1 0 0 0 1 1028
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_13
timestamp 1581321264
transform 1 0 0 0 1 720
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_14
timestamp 1581321264
transform 1 0 0 0 1 412
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_15
timestamp 1581321264
transform 1 0 0 0 1 104
box 44 -50 1800 299
<< labels >>
rlabel locali s 77 188 77 188 4 in_0
port 2 nsew
rlabel locali s 1765 188 1765 188 4 out_0
port 3 nsew
rlabel locali s 77 496 77 496 4 in_1
port 4 nsew
rlabel locali s 1765 496 1765 496 4 out_1
port 5 nsew
rlabel locali s 77 804 77 804 4 in_2
port 6 nsew
rlabel locali s 1765 804 1765 804 4 out_2
port 7 nsew
rlabel locali s 77 1112 77 1112 4 in_3
port 8 nsew
rlabel locali s 1765 1112 1765 1112 4 out_3
port 9 nsew
rlabel locali s 77 1420 77 1420 4 in_4
port 10 nsew
rlabel locali s 1765 1420 1765 1420 4 out_4
port 11 nsew
rlabel locali s 77 1728 77 1728 4 in_5
port 12 nsew
rlabel locali s 1765 1728 1765 1728 4 out_5
port 13 nsew
rlabel locali s 77 2036 77 2036 4 in_6
port 14 nsew
rlabel locali s 1765 2036 1765 2036 4 out_6
port 15 nsew
rlabel locali s 77 2344 77 2344 4 in_7
port 16 nsew
rlabel locali s 1765 2344 1765 2344 4 out_7
port 17 nsew
rlabel locali s 77 2652 77 2652 4 in_8
port 18 nsew
rlabel locali s 1765 2652 1765 2652 4 out_8
port 19 nsew
rlabel locali s 77 2960 77 2960 4 in_9
port 20 nsew
rlabel locali s 1765 2960 1765 2960 4 out_9
port 21 nsew
rlabel locali s 77 3268 77 3268 4 in_10
port 22 nsew
rlabel locali s 1765 3268 1765 3268 4 out_10
port 23 nsew
rlabel locali s 77 3576 77 3576 4 in_11
port 24 nsew
rlabel locali s 1765 3576 1765 3576 4 out_11
port 25 nsew
rlabel locali s 77 3884 77 3884 4 in_12
port 26 nsew
rlabel locali s 1765 3884 1765 3884 4 out_12
port 27 nsew
rlabel locali s 77 4192 77 4192 4 in_13
port 28 nsew
rlabel locali s 1765 4192 1765 4192 4 out_13
port 29 nsew
rlabel locali s 77 4500 77 4500 4 in_14
port 30 nsew
rlabel locali s 1765 4500 1765 4500 4 out_14
port 31 nsew
rlabel locali s 77 4808 77 4808 4 in_15
port 32 nsew
rlabel locali s 1765 4808 1765 4808 4 out_15
port 33 nsew
rlabel metal1 s 316 6 344 34 4 gnd
port 35 nsew
rlabel metal1 s 316 4914 344 4942 4 gnd
port 35 nsew
rlabel metal1 s 1232 6 1260 34 4 vdd
port 37 nsew
rlabel metal1 s 1232 4914 1260 4942 4 vdd
port 37 nsew
<< properties >>
string FIXED_BBOX 1162 -50 1330 0
<< end >>
