magic
tech sky130A
magscale 1 2
timestamp 1581365163
<< checkpaint >>
rect -1124 -1339 3139 53579
<< locali >>
rect 226 52071 260 52121
rect 1821 52071 1855 52137
rect 226 52037 297 52071
rect 226 51867 260 51917
rect 1821 51867 1855 51933
rect 226 51833 297 51867
rect 226 51663 260 51713
rect 1821 51663 1855 51729
rect 226 51629 297 51663
rect 226 51459 260 51509
rect 1821 51459 1855 51525
rect 226 51425 297 51459
rect 226 51255 260 51305
rect 1821 51255 1855 51321
rect 226 51221 297 51255
rect 226 51051 260 51101
rect 1821 51051 1855 51117
rect 226 51017 297 51051
rect 226 50847 260 50897
rect 1821 50847 1855 50913
rect 226 50813 297 50847
rect 226 50643 260 50693
rect 1821 50643 1855 50709
rect 226 50609 297 50643
rect 226 50439 260 50489
rect 1821 50439 1855 50505
rect 226 50405 297 50439
rect 226 50235 260 50285
rect 1821 50235 1855 50301
rect 226 50201 297 50235
rect 226 50031 260 50081
rect 1821 50031 1855 50097
rect 226 49997 297 50031
rect 226 49827 260 49877
rect 1821 49827 1855 49893
rect 226 49793 297 49827
rect 226 49623 260 49673
rect 1821 49623 1855 49689
rect 226 49589 297 49623
rect 226 49419 260 49469
rect 1821 49419 1855 49485
rect 226 49385 297 49419
rect 226 49215 260 49265
rect 1821 49215 1855 49281
rect 226 49181 297 49215
rect 226 49011 260 49061
rect 1821 49011 1855 49077
rect 226 48977 297 49011
rect 226 48807 260 48857
rect 1821 48807 1855 48873
rect 226 48773 297 48807
rect 226 48603 260 48653
rect 1821 48603 1855 48669
rect 226 48569 297 48603
rect 226 48399 260 48449
rect 1821 48399 1855 48465
rect 226 48365 297 48399
rect 226 48195 260 48245
rect 1821 48195 1855 48261
rect 226 48161 297 48195
rect 226 47991 260 48041
rect 1821 47991 1855 48057
rect 226 47957 297 47991
rect 226 47787 260 47837
rect 1821 47787 1855 47853
rect 226 47753 297 47787
rect 226 47583 260 47633
rect 1821 47583 1855 47649
rect 226 47549 297 47583
rect 226 47379 260 47429
rect 1821 47379 1855 47445
rect 226 47345 297 47379
rect 226 47175 260 47225
rect 1821 47175 1855 47241
rect 226 47141 297 47175
rect 226 46971 260 47021
rect 1821 46971 1855 47037
rect 226 46937 297 46971
rect 226 46767 260 46817
rect 1821 46767 1855 46833
rect 226 46733 297 46767
rect 226 46563 260 46613
rect 1821 46563 1855 46629
rect 226 46529 297 46563
rect 226 46359 260 46409
rect 1821 46359 1855 46425
rect 226 46325 297 46359
rect 226 46155 260 46205
rect 1821 46155 1855 46221
rect 226 46121 297 46155
rect 226 45951 260 46001
rect 1821 45951 1855 46017
rect 226 45917 297 45951
rect 226 45747 260 45797
rect 1821 45747 1855 45813
rect 226 45713 297 45747
rect 226 45543 260 45593
rect 1821 45543 1855 45609
rect 226 45509 297 45543
rect 226 45339 260 45389
rect 1821 45339 1855 45405
rect 226 45305 297 45339
rect 226 45135 260 45185
rect 1821 45135 1855 45201
rect 226 45101 297 45135
rect 226 44931 260 44981
rect 1821 44931 1855 44997
rect 226 44897 297 44931
rect 226 44727 260 44777
rect 1821 44727 1855 44793
rect 226 44693 297 44727
rect 226 44523 260 44573
rect 1821 44523 1855 44589
rect 226 44489 297 44523
rect 226 44319 260 44369
rect 1821 44319 1855 44385
rect 226 44285 297 44319
rect 226 44115 260 44165
rect 1821 44115 1855 44181
rect 226 44081 297 44115
rect 226 43911 260 43961
rect 1821 43911 1855 43977
rect 226 43877 297 43911
rect 226 43707 260 43757
rect 1821 43707 1855 43773
rect 226 43673 297 43707
rect 226 43503 260 43553
rect 1821 43503 1855 43569
rect 226 43469 297 43503
rect 226 43299 260 43349
rect 1821 43299 1855 43365
rect 226 43265 297 43299
rect 226 43095 260 43145
rect 1821 43095 1855 43161
rect 226 43061 297 43095
rect 226 42891 260 42941
rect 1821 42891 1855 42957
rect 226 42857 297 42891
rect 226 42687 260 42737
rect 1821 42687 1855 42753
rect 226 42653 297 42687
rect 226 42483 260 42533
rect 1821 42483 1855 42549
rect 226 42449 297 42483
rect 226 42279 260 42329
rect 1821 42279 1855 42345
rect 226 42245 297 42279
rect 226 42075 260 42125
rect 1821 42075 1855 42141
rect 226 42041 297 42075
rect 226 41871 260 41921
rect 1821 41871 1855 41937
rect 226 41837 297 41871
rect 226 41667 260 41717
rect 1821 41667 1855 41733
rect 226 41633 297 41667
rect 226 41463 260 41513
rect 1821 41463 1855 41529
rect 226 41429 297 41463
rect 226 41259 260 41309
rect 1821 41259 1855 41325
rect 226 41225 297 41259
rect 226 41055 260 41105
rect 1821 41055 1855 41121
rect 226 41021 297 41055
rect 226 40851 260 40901
rect 1821 40851 1855 40917
rect 226 40817 297 40851
rect 226 40647 260 40697
rect 1821 40647 1855 40713
rect 226 40613 297 40647
rect 226 40443 260 40493
rect 1821 40443 1855 40509
rect 226 40409 297 40443
rect 226 40239 260 40289
rect 1821 40239 1855 40305
rect 226 40205 297 40239
rect 226 40035 260 40085
rect 1821 40035 1855 40101
rect 226 40001 297 40035
rect 226 39831 260 39881
rect 1821 39831 1855 39897
rect 226 39797 297 39831
rect 226 39627 260 39677
rect 1821 39627 1855 39693
rect 226 39593 297 39627
rect 226 39423 260 39473
rect 1821 39423 1855 39489
rect 226 39389 297 39423
rect 226 39219 260 39269
rect 1821 39219 1855 39285
rect 226 39185 297 39219
rect 226 39015 260 39065
rect 1821 39015 1855 39081
rect 226 38981 297 39015
rect 226 38811 260 38861
rect 1821 38811 1855 38877
rect 226 38777 297 38811
rect 226 38607 260 38657
rect 1821 38607 1855 38673
rect 226 38573 297 38607
rect 226 38403 260 38453
rect 1821 38403 1855 38469
rect 226 38369 297 38403
rect 226 38199 260 38249
rect 1821 38199 1855 38265
rect 226 38165 297 38199
rect 226 37995 260 38045
rect 1821 37995 1855 38061
rect 226 37961 297 37995
rect 226 37791 260 37841
rect 1821 37791 1855 37857
rect 226 37757 297 37791
rect 226 37587 260 37637
rect 1821 37587 1855 37653
rect 226 37553 297 37587
rect 226 37383 260 37433
rect 1821 37383 1855 37449
rect 226 37349 297 37383
rect 226 37179 260 37229
rect 1821 37179 1855 37245
rect 226 37145 297 37179
rect 226 36975 260 37025
rect 1821 36975 1855 37041
rect 226 36941 297 36975
rect 226 36771 260 36821
rect 1821 36771 1855 36837
rect 226 36737 297 36771
rect 226 36567 260 36617
rect 1821 36567 1855 36633
rect 226 36533 297 36567
rect 226 36363 260 36413
rect 1821 36363 1855 36429
rect 226 36329 297 36363
rect 226 36159 260 36209
rect 1821 36159 1855 36225
rect 226 36125 297 36159
rect 226 35955 260 36005
rect 1821 35955 1855 36021
rect 226 35921 297 35955
rect 226 35751 260 35801
rect 1821 35751 1855 35817
rect 226 35717 297 35751
rect 226 35547 260 35597
rect 1821 35547 1855 35613
rect 226 35513 297 35547
rect 226 35343 260 35393
rect 1821 35343 1855 35409
rect 226 35309 297 35343
rect 226 35139 260 35189
rect 1821 35139 1855 35205
rect 226 35105 297 35139
rect 226 34935 260 34985
rect 1821 34935 1855 35001
rect 226 34901 297 34935
rect 226 34731 260 34781
rect 1821 34731 1855 34797
rect 226 34697 297 34731
rect 226 34527 260 34577
rect 1821 34527 1855 34593
rect 226 34493 297 34527
rect 226 34323 260 34373
rect 1821 34323 1855 34389
rect 226 34289 297 34323
rect 226 34119 260 34169
rect 1821 34119 1855 34185
rect 226 34085 297 34119
rect 226 33915 260 33965
rect 1821 33915 1855 33981
rect 226 33881 297 33915
rect 226 33711 260 33761
rect 1821 33711 1855 33777
rect 226 33677 297 33711
rect 226 33507 260 33557
rect 1821 33507 1855 33573
rect 226 33473 297 33507
rect 226 33303 260 33353
rect 1821 33303 1855 33369
rect 226 33269 297 33303
rect 226 33099 260 33149
rect 1821 33099 1855 33165
rect 226 33065 297 33099
rect 226 32895 260 32945
rect 1821 32895 1855 32961
rect 226 32861 297 32895
rect 226 32691 260 32741
rect 1821 32691 1855 32757
rect 226 32657 297 32691
rect 226 32487 260 32537
rect 1821 32487 1855 32553
rect 226 32453 297 32487
rect 226 32283 260 32333
rect 1821 32283 1855 32349
rect 226 32249 297 32283
rect 226 32079 260 32129
rect 1821 32079 1855 32145
rect 226 32045 297 32079
rect 226 31875 260 31925
rect 1821 31875 1855 31941
rect 226 31841 297 31875
rect 226 31671 260 31721
rect 1821 31671 1855 31737
rect 226 31637 297 31671
rect 226 31467 260 31517
rect 1821 31467 1855 31533
rect 226 31433 297 31467
rect 226 31263 260 31313
rect 1821 31263 1855 31329
rect 226 31229 297 31263
rect 226 31059 260 31109
rect 1821 31059 1855 31125
rect 226 31025 297 31059
rect 226 30855 260 30905
rect 1821 30855 1855 30921
rect 226 30821 297 30855
rect 226 30651 260 30701
rect 1821 30651 1855 30717
rect 226 30617 297 30651
rect 226 30447 260 30497
rect 1821 30447 1855 30513
rect 226 30413 297 30447
rect 226 30243 260 30293
rect 1821 30243 1855 30309
rect 226 30209 297 30243
rect 226 30039 260 30089
rect 1821 30039 1855 30105
rect 226 30005 297 30039
rect 226 29835 260 29885
rect 1821 29835 1855 29901
rect 226 29801 297 29835
rect 226 29631 260 29681
rect 1821 29631 1855 29697
rect 226 29597 297 29631
rect 226 29427 260 29477
rect 1821 29427 1855 29493
rect 226 29393 297 29427
rect 226 29223 260 29273
rect 1821 29223 1855 29289
rect 226 29189 297 29223
rect 226 29019 260 29069
rect 1821 29019 1855 29085
rect 226 28985 297 29019
rect 226 28815 260 28865
rect 1821 28815 1855 28881
rect 226 28781 297 28815
rect 226 28611 260 28661
rect 1821 28611 1855 28677
rect 226 28577 297 28611
rect 226 28407 260 28457
rect 1821 28407 1855 28473
rect 226 28373 297 28407
rect 226 28203 260 28253
rect 1821 28203 1855 28269
rect 226 28169 297 28203
rect 226 27999 260 28049
rect 1821 27999 1855 28065
rect 226 27965 297 27999
rect 226 27795 260 27845
rect 1821 27795 1855 27861
rect 226 27761 297 27795
rect 226 27591 260 27641
rect 1821 27591 1855 27657
rect 226 27557 297 27591
rect 226 27387 260 27437
rect 1821 27387 1855 27453
rect 226 27353 297 27387
rect 226 27183 260 27233
rect 1821 27183 1855 27249
rect 226 27149 297 27183
rect 226 26979 260 27029
rect 1821 26979 1855 27045
rect 226 26945 297 26979
rect 226 26775 260 26825
rect 1821 26775 1855 26841
rect 226 26741 297 26775
rect 226 26571 260 26621
rect 1821 26571 1855 26637
rect 226 26537 297 26571
rect 226 26367 260 26417
rect 1821 26367 1855 26433
rect 226 26333 297 26367
rect 226 26163 260 26213
rect 1821 26163 1855 26229
rect 226 26129 297 26163
rect 226 25959 260 26009
rect 1821 25959 1855 26025
rect 226 25925 297 25959
rect 226 25755 260 25805
rect 1821 25755 1855 25821
rect 226 25721 297 25755
rect 226 25551 260 25601
rect 1821 25551 1855 25617
rect 226 25517 297 25551
rect 226 25347 260 25397
rect 1821 25347 1855 25413
rect 226 25313 297 25347
rect 226 25143 260 25193
rect 1821 25143 1855 25209
rect 226 25109 297 25143
rect 226 24939 260 24989
rect 1821 24939 1855 25005
rect 226 24905 297 24939
rect 226 24735 260 24785
rect 1821 24735 1855 24801
rect 226 24701 297 24735
rect 226 24531 260 24581
rect 1821 24531 1855 24597
rect 226 24497 297 24531
rect 226 24327 260 24377
rect 1821 24327 1855 24393
rect 226 24293 297 24327
rect 226 24123 260 24173
rect 1821 24123 1855 24189
rect 226 24089 297 24123
rect 226 23919 260 23969
rect 1821 23919 1855 23985
rect 226 23885 297 23919
rect 226 23715 260 23765
rect 1821 23715 1855 23781
rect 226 23681 297 23715
rect 226 23511 260 23561
rect 1821 23511 1855 23577
rect 226 23477 297 23511
rect 226 23307 260 23357
rect 1821 23307 1855 23373
rect 226 23273 297 23307
rect 226 23103 260 23153
rect 1821 23103 1855 23169
rect 226 23069 297 23103
rect 226 22899 260 22949
rect 1821 22899 1855 22965
rect 226 22865 297 22899
rect 226 22695 260 22745
rect 1821 22695 1855 22761
rect 226 22661 297 22695
rect 226 22491 260 22541
rect 1821 22491 1855 22557
rect 226 22457 297 22491
rect 226 22287 260 22337
rect 1821 22287 1855 22353
rect 226 22253 297 22287
rect 226 22083 260 22133
rect 1821 22083 1855 22149
rect 226 22049 297 22083
rect 226 21879 260 21929
rect 1821 21879 1855 21945
rect 226 21845 297 21879
rect 226 21675 260 21725
rect 1821 21675 1855 21741
rect 226 21641 297 21675
rect 226 21471 260 21521
rect 1821 21471 1855 21537
rect 226 21437 297 21471
rect 226 21267 260 21317
rect 1821 21267 1855 21333
rect 226 21233 297 21267
rect 226 21063 260 21113
rect 1821 21063 1855 21129
rect 226 21029 297 21063
rect 226 20859 260 20909
rect 1821 20859 1855 20925
rect 226 20825 297 20859
rect 226 20655 260 20705
rect 1821 20655 1855 20721
rect 226 20621 297 20655
rect 226 20451 260 20501
rect 1821 20451 1855 20517
rect 226 20417 297 20451
rect 226 20247 260 20297
rect 1821 20247 1855 20313
rect 226 20213 297 20247
rect 226 20043 260 20093
rect 1821 20043 1855 20109
rect 226 20009 297 20043
rect 226 19839 260 19889
rect 1821 19839 1855 19905
rect 226 19805 297 19839
rect 226 19635 260 19685
rect 1821 19635 1855 19701
rect 226 19601 297 19635
rect 226 19431 260 19481
rect 1821 19431 1855 19497
rect 226 19397 297 19431
rect 226 19227 260 19277
rect 1821 19227 1855 19293
rect 226 19193 297 19227
rect 226 19023 260 19073
rect 1821 19023 1855 19089
rect 226 18989 297 19023
rect 226 18819 260 18869
rect 1821 18819 1855 18885
rect 226 18785 297 18819
rect 226 18615 260 18665
rect 1821 18615 1855 18681
rect 226 18581 297 18615
rect 226 18411 260 18461
rect 1821 18411 1855 18477
rect 226 18377 297 18411
rect 226 18207 260 18257
rect 1821 18207 1855 18273
rect 226 18173 297 18207
rect 226 18003 260 18053
rect 1821 18003 1855 18069
rect 226 17969 297 18003
rect 226 17799 260 17849
rect 1821 17799 1855 17865
rect 226 17765 297 17799
rect 226 17595 260 17645
rect 1821 17595 1855 17661
rect 226 17561 297 17595
rect 226 17391 260 17441
rect 1821 17391 1855 17457
rect 226 17357 297 17391
rect 226 17187 260 17237
rect 1821 17187 1855 17253
rect 226 17153 297 17187
rect 226 16983 260 17033
rect 1821 16983 1855 17049
rect 226 16949 297 16983
rect 226 16779 260 16829
rect 1821 16779 1855 16845
rect 226 16745 297 16779
rect 226 16575 260 16625
rect 1821 16575 1855 16641
rect 226 16541 297 16575
rect 226 16371 260 16421
rect 1821 16371 1855 16437
rect 226 16337 297 16371
rect 226 16167 260 16217
rect 1821 16167 1855 16233
rect 226 16133 297 16167
rect 226 15963 260 16013
rect 1821 15963 1855 16029
rect 226 15929 297 15963
rect 226 15759 260 15809
rect 1821 15759 1855 15825
rect 226 15725 297 15759
rect 226 15555 260 15605
rect 1821 15555 1855 15621
rect 226 15521 297 15555
rect 226 15351 260 15401
rect 1821 15351 1855 15417
rect 226 15317 297 15351
rect 226 15147 260 15197
rect 1821 15147 1855 15213
rect 226 15113 297 15147
rect 226 14943 260 14993
rect 1821 14943 1855 15009
rect 226 14909 297 14943
rect 226 14739 260 14789
rect 1821 14739 1855 14805
rect 226 14705 297 14739
rect 226 14535 260 14585
rect 1821 14535 1855 14601
rect 226 14501 297 14535
rect 226 14331 260 14381
rect 1821 14331 1855 14397
rect 226 14297 297 14331
rect 226 14127 260 14177
rect 1821 14127 1855 14193
rect 226 14093 297 14127
rect 226 13923 260 13973
rect 1821 13923 1855 13989
rect 226 13889 297 13923
rect 226 13719 260 13769
rect 1821 13719 1855 13785
rect 226 13685 297 13719
rect 226 13515 260 13565
rect 1821 13515 1855 13581
rect 226 13481 297 13515
rect 226 13311 260 13361
rect 1821 13311 1855 13377
rect 226 13277 297 13311
rect 226 13107 260 13157
rect 1821 13107 1855 13173
rect 226 13073 297 13107
rect 226 12903 260 12953
rect 1821 12903 1855 12969
rect 226 12869 297 12903
rect 226 12699 260 12749
rect 1821 12699 1855 12765
rect 226 12665 297 12699
rect 226 12495 260 12545
rect 1821 12495 1855 12561
rect 226 12461 297 12495
rect 226 12291 260 12341
rect 1821 12291 1855 12357
rect 226 12257 297 12291
rect 226 12087 260 12137
rect 1821 12087 1855 12153
rect 226 12053 297 12087
rect 226 11883 260 11933
rect 1821 11883 1855 11949
rect 226 11849 297 11883
rect 226 11679 260 11729
rect 1821 11679 1855 11745
rect 226 11645 297 11679
rect 226 11475 260 11525
rect 1821 11475 1855 11541
rect 226 11441 297 11475
rect 226 11271 260 11321
rect 1821 11271 1855 11337
rect 226 11237 297 11271
rect 226 11067 260 11117
rect 1821 11067 1855 11133
rect 226 11033 297 11067
rect 226 10863 260 10913
rect 1821 10863 1855 10929
rect 226 10829 297 10863
rect 226 10659 260 10709
rect 1821 10659 1855 10725
rect 226 10625 297 10659
rect 226 10455 260 10505
rect 1821 10455 1855 10521
rect 226 10421 297 10455
rect 226 10251 260 10301
rect 1821 10251 1855 10317
rect 226 10217 297 10251
rect 226 10047 260 10097
rect 1821 10047 1855 10113
rect 226 10013 297 10047
rect 226 9843 260 9893
rect 1821 9843 1855 9909
rect 226 9809 297 9843
rect 226 9639 260 9689
rect 1821 9639 1855 9705
rect 226 9605 297 9639
rect 226 9435 260 9485
rect 1821 9435 1855 9501
rect 226 9401 297 9435
rect 226 9231 260 9281
rect 1821 9231 1855 9297
rect 226 9197 297 9231
rect 226 9027 260 9077
rect 1821 9027 1855 9093
rect 226 8993 297 9027
rect 226 8823 260 8873
rect 1821 8823 1855 8889
rect 226 8789 297 8823
rect 226 8619 260 8669
rect 1821 8619 1855 8685
rect 226 8585 297 8619
rect 226 8415 260 8465
rect 1821 8415 1855 8481
rect 226 8381 297 8415
rect 226 8211 260 8261
rect 1821 8211 1855 8277
rect 226 8177 297 8211
rect 226 8007 260 8057
rect 1821 8007 1855 8073
rect 226 7973 297 8007
rect 226 7803 260 7853
rect 1821 7803 1855 7869
rect 226 7769 297 7803
rect 226 7599 260 7649
rect 1821 7599 1855 7665
rect 226 7565 297 7599
rect 226 7395 260 7445
rect 1821 7395 1855 7461
rect 226 7361 297 7395
rect 226 7191 260 7241
rect 1821 7191 1855 7257
rect 226 7157 297 7191
rect 226 6987 260 7037
rect 1821 6987 1855 7053
rect 226 6953 297 6987
rect 226 6783 260 6833
rect 1821 6783 1855 6849
rect 226 6749 297 6783
rect 226 6579 260 6629
rect 1821 6579 1855 6645
rect 226 6545 297 6579
rect 226 6375 260 6425
rect 1821 6375 1855 6441
rect 226 6341 297 6375
rect 226 6171 260 6221
rect 1821 6171 1855 6237
rect 226 6137 297 6171
rect 226 5967 260 6017
rect 1821 5967 1855 6033
rect 226 5933 297 5967
rect 226 5763 260 5813
rect 1821 5763 1855 5829
rect 226 5729 297 5763
rect 226 5559 260 5609
rect 1821 5559 1855 5625
rect 226 5525 297 5559
rect 226 5355 260 5405
rect 1821 5355 1855 5421
rect 226 5321 297 5355
rect 226 5151 260 5201
rect 1821 5151 1855 5217
rect 226 5117 297 5151
rect 226 4947 260 4997
rect 1821 4947 1855 5013
rect 226 4913 297 4947
rect 226 4743 260 4793
rect 1821 4743 1855 4809
rect 226 4709 297 4743
rect 226 4539 260 4589
rect 1821 4539 1855 4605
rect 226 4505 297 4539
rect 226 4335 260 4385
rect 1821 4335 1855 4401
rect 226 4301 297 4335
rect 226 4131 260 4181
rect 1821 4131 1855 4197
rect 226 4097 297 4131
rect 226 3927 260 3977
rect 1821 3927 1855 3993
rect 226 3893 297 3927
rect 226 3723 260 3773
rect 1821 3723 1855 3789
rect 226 3689 297 3723
rect 226 3519 260 3569
rect 1821 3519 1855 3585
rect 226 3485 297 3519
rect 226 3315 260 3365
rect 1821 3315 1855 3381
rect 226 3281 297 3315
rect 226 3111 260 3161
rect 1821 3111 1855 3177
rect 226 3077 297 3111
rect 226 2907 260 2957
rect 1821 2907 1855 2973
rect 226 2873 297 2907
rect 226 2703 260 2753
rect 1821 2703 1855 2769
rect 226 2669 297 2703
rect 226 2499 260 2549
rect 1821 2499 1855 2565
rect 226 2465 297 2499
rect 226 2295 260 2345
rect 1821 2295 1855 2361
rect 226 2261 297 2295
rect 226 2091 260 2141
rect 1821 2091 1855 2157
rect 226 2057 297 2091
rect 226 1887 260 1937
rect 1821 1887 1855 1953
rect 226 1853 297 1887
rect 226 1683 260 1733
rect 1821 1683 1855 1749
rect 226 1649 297 1683
rect 226 1479 260 1529
rect 1821 1479 1855 1545
rect 226 1445 297 1479
rect 226 1275 260 1325
rect 1821 1275 1855 1341
rect 226 1241 297 1275
rect 226 1071 260 1121
rect 1821 1071 1855 1137
rect 226 1037 297 1071
rect 226 867 260 917
rect 1821 867 1855 933
rect 226 833 297 867
rect 226 663 260 713
rect 1821 663 1855 729
rect 226 629 297 663
rect 226 459 260 509
rect 1821 459 1855 525
rect 226 425 297 459
rect 226 255 260 305
rect 1821 255 1855 321
rect 226 221 297 255
rect 226 51 260 101
rect 1821 51 1855 117
rect 226 17 297 51
<< metal1 >>
rect 316 -14 344 52238
rect 1232 -14 1260 52238
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_0
timestamp 1581365163
transform 1 0 0 0 1 52020
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_1
timestamp 1581365163
transform 1 0 0 0 1 51816
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_2
timestamp 1581365163
transform 1 0 0 0 1 51612
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_3
timestamp 1581365163
transform 1 0 0 0 1 51408
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_4
timestamp 1581365163
transform 1 0 0 0 1 51204
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_5
timestamp 1581365163
transform 1 0 0 0 1 51000
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_6
timestamp 1581365163
transform 1 0 0 0 1 50796
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_7
timestamp 1581365163
transform 1 0 0 0 1 50592
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_8
timestamp 1581365163
transform 1 0 0 0 1 50388
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_9
timestamp 1581365163
transform 1 0 0 0 1 50184
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_10
timestamp 1581365163
transform 1 0 0 0 1 49980
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_11
timestamp 1581365163
transform 1 0 0 0 1 49776
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_12
timestamp 1581365163
transform 1 0 0 0 1 49572
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_13
timestamp 1581365163
transform 1 0 0 0 1 49368
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_14
timestamp 1581365163
transform 1 0 0 0 1 49164
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_15
timestamp 1581365163
transform 1 0 0 0 1 48960
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_16
timestamp 1581365163
transform 1 0 0 0 1 48756
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_17
timestamp 1581365163
transform 1 0 0 0 1 48552
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_18
timestamp 1581365163
transform 1 0 0 0 1 48348
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_19
timestamp 1581365163
transform 1 0 0 0 1 48144
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_20
timestamp 1581365163
transform 1 0 0 0 1 47940
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_21
timestamp 1581365163
transform 1 0 0 0 1 47736
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_22
timestamp 1581365163
transform 1 0 0 0 1 47532
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_23
timestamp 1581365163
transform 1 0 0 0 1 47328
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_24
timestamp 1581365163
transform 1 0 0 0 1 47124
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_25
timestamp 1581365163
transform 1 0 0 0 1 46920
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_26
timestamp 1581365163
transform 1 0 0 0 1 46716
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_27
timestamp 1581365163
transform 1 0 0 0 1 46512
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_28
timestamp 1581365163
transform 1 0 0 0 1 46308
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_29
timestamp 1581365163
transform 1 0 0 0 1 46104
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_30
timestamp 1581365163
transform 1 0 0 0 1 45900
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_31
timestamp 1581365163
transform 1 0 0 0 1 45696
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_32
timestamp 1581365163
transform 1 0 0 0 1 45492
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_33
timestamp 1581365163
transform 1 0 0 0 1 45288
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_34
timestamp 1581365163
transform 1 0 0 0 1 45084
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_35
timestamp 1581365163
transform 1 0 0 0 1 44880
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_36
timestamp 1581365163
transform 1 0 0 0 1 44676
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_37
timestamp 1581365163
transform 1 0 0 0 1 44472
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_38
timestamp 1581365163
transform 1 0 0 0 1 44268
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_39
timestamp 1581365163
transform 1 0 0 0 1 44064
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_40
timestamp 1581365163
transform 1 0 0 0 1 43860
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_41
timestamp 1581365163
transform 1 0 0 0 1 43656
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_42
timestamp 1581365163
transform 1 0 0 0 1 43452
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_43
timestamp 1581365163
transform 1 0 0 0 1 43248
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_44
timestamp 1581365163
transform 1 0 0 0 1 43044
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_45
timestamp 1581365163
transform 1 0 0 0 1 42840
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_46
timestamp 1581365163
transform 1 0 0 0 1 42636
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_47
timestamp 1581365163
transform 1 0 0 0 1 42432
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_48
timestamp 1581365163
transform 1 0 0 0 1 42228
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_49
timestamp 1581365163
transform 1 0 0 0 1 42024
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_50
timestamp 1581365163
transform 1 0 0 0 1 41820
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_51
timestamp 1581365163
transform 1 0 0 0 1 41616
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_52
timestamp 1581365163
transform 1 0 0 0 1 41412
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_53
timestamp 1581365163
transform 1 0 0 0 1 41208
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_54
timestamp 1581365163
transform 1 0 0 0 1 41004
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_55
timestamp 1581365163
transform 1 0 0 0 1 40800
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_56
timestamp 1581365163
transform 1 0 0 0 1 40596
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_57
timestamp 1581365163
transform 1 0 0 0 1 40392
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_58
timestamp 1581365163
transform 1 0 0 0 1 40188
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_59
timestamp 1581365163
transform 1 0 0 0 1 39984
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_60
timestamp 1581365163
transform 1 0 0 0 1 39780
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_61
timestamp 1581365163
transform 1 0 0 0 1 39576
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_62
timestamp 1581365163
transform 1 0 0 0 1 39372
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_63
timestamp 1581365163
transform 1 0 0 0 1 39168
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_64
timestamp 1581365163
transform 1 0 0 0 1 38964
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_65
timestamp 1581365163
transform 1 0 0 0 1 38760
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_66
timestamp 1581365163
transform 1 0 0 0 1 38556
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_67
timestamp 1581365163
transform 1 0 0 0 1 38352
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_68
timestamp 1581365163
transform 1 0 0 0 1 38148
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_69
timestamp 1581365163
transform 1 0 0 0 1 37944
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_70
timestamp 1581365163
transform 1 0 0 0 1 37740
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_71
timestamp 1581365163
transform 1 0 0 0 1 37536
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_72
timestamp 1581365163
transform 1 0 0 0 1 37332
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_73
timestamp 1581365163
transform 1 0 0 0 1 37128
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_74
timestamp 1581365163
transform 1 0 0 0 1 36924
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_75
timestamp 1581365163
transform 1 0 0 0 1 36720
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_76
timestamp 1581365163
transform 1 0 0 0 1 36516
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_77
timestamp 1581365163
transform 1 0 0 0 1 36312
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_78
timestamp 1581365163
transform 1 0 0 0 1 36108
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_79
timestamp 1581365163
transform 1 0 0 0 1 35904
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_80
timestamp 1581365163
transform 1 0 0 0 1 35700
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_81
timestamp 1581365163
transform 1 0 0 0 1 35496
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_82
timestamp 1581365163
transform 1 0 0 0 1 35292
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_83
timestamp 1581365163
transform 1 0 0 0 1 35088
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_84
timestamp 1581365163
transform 1 0 0 0 1 34884
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_85
timestamp 1581365163
transform 1 0 0 0 1 34680
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_86
timestamp 1581365163
transform 1 0 0 0 1 34476
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_87
timestamp 1581365163
transform 1 0 0 0 1 34272
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_88
timestamp 1581365163
transform 1 0 0 0 1 34068
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_89
timestamp 1581365163
transform 1 0 0 0 1 33864
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_90
timestamp 1581365163
transform 1 0 0 0 1 33660
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_91
timestamp 1581365163
transform 1 0 0 0 1 33456
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_92
timestamp 1581365163
transform 1 0 0 0 1 33252
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_93
timestamp 1581365163
transform 1 0 0 0 1 33048
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_94
timestamp 1581365163
transform 1 0 0 0 1 32844
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_95
timestamp 1581365163
transform 1 0 0 0 1 32640
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_96
timestamp 1581365163
transform 1 0 0 0 1 32436
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_97
timestamp 1581365163
transform 1 0 0 0 1 32232
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_98
timestamp 1581365163
transform 1 0 0 0 1 32028
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_99
timestamp 1581365163
transform 1 0 0 0 1 31824
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_100
timestamp 1581365163
transform 1 0 0 0 1 31620
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_101
timestamp 1581365163
transform 1 0 0 0 1 31416
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_102
timestamp 1581365163
transform 1 0 0 0 1 31212
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_103
timestamp 1581365163
transform 1 0 0 0 1 31008
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_104
timestamp 1581365163
transform 1 0 0 0 1 30804
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_105
timestamp 1581365163
transform 1 0 0 0 1 30600
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_106
timestamp 1581365163
transform 1 0 0 0 1 30396
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_107
timestamp 1581365163
transform 1 0 0 0 1 30192
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_108
timestamp 1581365163
transform 1 0 0 0 1 29988
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_109
timestamp 1581365163
transform 1 0 0 0 1 29784
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_110
timestamp 1581365163
transform 1 0 0 0 1 29580
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_111
timestamp 1581365163
transform 1 0 0 0 1 29376
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_112
timestamp 1581365163
transform 1 0 0 0 1 29172
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_113
timestamp 1581365163
transform 1 0 0 0 1 28968
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_114
timestamp 1581365163
transform 1 0 0 0 1 28764
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_115
timestamp 1581365163
transform 1 0 0 0 1 28560
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_116
timestamp 1581365163
transform 1 0 0 0 1 28356
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_117
timestamp 1581365163
transform 1 0 0 0 1 28152
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_118
timestamp 1581365163
transform 1 0 0 0 1 27948
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_119
timestamp 1581365163
transform 1 0 0 0 1 27744
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_120
timestamp 1581365163
transform 1 0 0 0 1 27540
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_121
timestamp 1581365163
transform 1 0 0 0 1 27336
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_122
timestamp 1581365163
transform 1 0 0 0 1 27132
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_123
timestamp 1581365163
transform 1 0 0 0 1 26928
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_124
timestamp 1581365163
transform 1 0 0 0 1 26724
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_125
timestamp 1581365163
transform 1 0 0 0 1 26520
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_126
timestamp 1581365163
transform 1 0 0 0 1 26316
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_127
timestamp 1581365163
transform 1 0 0 0 1 26112
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_128
timestamp 1581365163
transform 1 0 0 0 1 25908
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_129
timestamp 1581365163
transform 1 0 0 0 1 25704
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_130
timestamp 1581365163
transform 1 0 0 0 1 25500
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_131
timestamp 1581365163
transform 1 0 0 0 1 25296
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_132
timestamp 1581365163
transform 1 0 0 0 1 25092
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_133
timestamp 1581365163
transform 1 0 0 0 1 24888
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_134
timestamp 1581365163
transform 1 0 0 0 1 24684
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_135
timestamp 1581365163
transform 1 0 0 0 1 24480
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_136
timestamp 1581365163
transform 1 0 0 0 1 24276
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_137
timestamp 1581365163
transform 1 0 0 0 1 24072
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_138
timestamp 1581365163
transform 1 0 0 0 1 23868
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_139
timestamp 1581365163
transform 1 0 0 0 1 23664
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_140
timestamp 1581365163
transform 1 0 0 0 1 23460
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_141
timestamp 1581365163
transform 1 0 0 0 1 23256
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_142
timestamp 1581365163
transform 1 0 0 0 1 23052
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_143
timestamp 1581365163
transform 1 0 0 0 1 22848
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_144
timestamp 1581365163
transform 1 0 0 0 1 22644
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_145
timestamp 1581365163
transform 1 0 0 0 1 22440
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_146
timestamp 1581365163
transform 1 0 0 0 1 22236
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_147
timestamp 1581365163
transform 1 0 0 0 1 22032
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_148
timestamp 1581365163
transform 1 0 0 0 1 21828
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_149
timestamp 1581365163
transform 1 0 0 0 1 21624
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_150
timestamp 1581365163
transform 1 0 0 0 1 21420
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_151
timestamp 1581365163
transform 1 0 0 0 1 21216
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_152
timestamp 1581365163
transform 1 0 0 0 1 21012
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_153
timestamp 1581365163
transform 1 0 0 0 1 20808
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_154
timestamp 1581365163
transform 1 0 0 0 1 20604
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_155
timestamp 1581365163
transform 1 0 0 0 1 20400
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_156
timestamp 1581365163
transform 1 0 0 0 1 20196
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_157
timestamp 1581365163
transform 1 0 0 0 1 19992
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_158
timestamp 1581365163
transform 1 0 0 0 1 19788
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_159
timestamp 1581365163
transform 1 0 0 0 1 19584
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_160
timestamp 1581365163
transform 1 0 0 0 1 19380
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_161
timestamp 1581365163
transform 1 0 0 0 1 19176
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_162
timestamp 1581365163
transform 1 0 0 0 1 18972
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_163
timestamp 1581365163
transform 1 0 0 0 1 18768
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_164
timestamp 1581365163
transform 1 0 0 0 1 18564
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_165
timestamp 1581365163
transform 1 0 0 0 1 18360
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_166
timestamp 1581365163
transform 1 0 0 0 1 18156
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_167
timestamp 1581365163
transform 1 0 0 0 1 17952
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_168
timestamp 1581365163
transform 1 0 0 0 1 17748
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_169
timestamp 1581365163
transform 1 0 0 0 1 17544
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_170
timestamp 1581365163
transform 1 0 0 0 1 17340
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_171
timestamp 1581365163
transform 1 0 0 0 1 17136
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_172
timestamp 1581365163
transform 1 0 0 0 1 16932
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_173
timestamp 1581365163
transform 1 0 0 0 1 16728
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_174
timestamp 1581365163
transform 1 0 0 0 1 16524
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_175
timestamp 1581365163
transform 1 0 0 0 1 16320
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_176
timestamp 1581365163
transform 1 0 0 0 1 16116
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_177
timestamp 1581365163
transform 1 0 0 0 1 15912
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_178
timestamp 1581365163
transform 1 0 0 0 1 15708
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_179
timestamp 1581365163
transform 1 0 0 0 1 15504
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_180
timestamp 1581365163
transform 1 0 0 0 1 15300
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_181
timestamp 1581365163
transform 1 0 0 0 1 15096
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_182
timestamp 1581365163
transform 1 0 0 0 1 14892
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_183
timestamp 1581365163
transform 1 0 0 0 1 14688
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_184
timestamp 1581365163
transform 1 0 0 0 1 14484
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_185
timestamp 1581365163
transform 1 0 0 0 1 14280
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_186
timestamp 1581365163
transform 1 0 0 0 1 14076
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_187
timestamp 1581365163
transform 1 0 0 0 1 13872
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_188
timestamp 1581365163
transform 1 0 0 0 1 13668
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_189
timestamp 1581365163
transform 1 0 0 0 1 13464
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_190
timestamp 1581365163
transform 1 0 0 0 1 13260
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_191
timestamp 1581365163
transform 1 0 0 0 1 13056
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_192
timestamp 1581365163
transform 1 0 0 0 1 12852
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_193
timestamp 1581365163
transform 1 0 0 0 1 12648
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_194
timestamp 1581365163
transform 1 0 0 0 1 12444
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_195
timestamp 1581365163
transform 1 0 0 0 1 12240
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_196
timestamp 1581365163
transform 1 0 0 0 1 12036
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_197
timestamp 1581365163
transform 1 0 0 0 1 11832
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_198
timestamp 1581365163
transform 1 0 0 0 1 11628
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_199
timestamp 1581365163
transform 1 0 0 0 1 11424
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_200
timestamp 1581365163
transform 1 0 0 0 1 11220
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_201
timestamp 1581365163
transform 1 0 0 0 1 11016
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_202
timestamp 1581365163
transform 1 0 0 0 1 10812
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_203
timestamp 1581365163
transform 1 0 0 0 1 10608
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_204
timestamp 1581365163
transform 1 0 0 0 1 10404
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_205
timestamp 1581365163
transform 1 0 0 0 1 10200
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_206
timestamp 1581365163
transform 1 0 0 0 1 9996
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_207
timestamp 1581365163
transform 1 0 0 0 1 9792
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_208
timestamp 1581365163
transform 1 0 0 0 1 9588
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_209
timestamp 1581365163
transform 1 0 0 0 1 9384
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_210
timestamp 1581365163
transform 1 0 0 0 1 9180
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_211
timestamp 1581365163
transform 1 0 0 0 1 8976
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_212
timestamp 1581365163
transform 1 0 0 0 1 8772
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_213
timestamp 1581365163
transform 1 0 0 0 1 8568
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_214
timestamp 1581365163
transform 1 0 0 0 1 8364
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_215
timestamp 1581365163
transform 1 0 0 0 1 8160
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_216
timestamp 1581365163
transform 1 0 0 0 1 7956
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_217
timestamp 1581365163
transform 1 0 0 0 1 7752
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_218
timestamp 1581365163
transform 1 0 0 0 1 7548
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_219
timestamp 1581365163
transform 1 0 0 0 1 7344
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_220
timestamp 1581365163
transform 1 0 0 0 1 7140
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_221
timestamp 1581365163
transform 1 0 0 0 1 6936
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_222
timestamp 1581365163
transform 1 0 0 0 1 6732
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_223
timestamp 1581365163
transform 1 0 0 0 1 6528
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_224
timestamp 1581365163
transform 1 0 0 0 1 6324
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_225
timestamp 1581365163
transform 1 0 0 0 1 6120
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_226
timestamp 1581365163
transform 1 0 0 0 1 5916
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_227
timestamp 1581365163
transform 1 0 0 0 1 5712
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_228
timestamp 1581365163
transform 1 0 0 0 1 5508
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_229
timestamp 1581365163
transform 1 0 0 0 1 5304
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_230
timestamp 1581365163
transform 1 0 0 0 1 5100
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_231
timestamp 1581365163
transform 1 0 0 0 1 4896
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_232
timestamp 1581365163
transform 1 0 0 0 1 4692
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_233
timestamp 1581365163
transform 1 0 0 0 1 4488
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_234
timestamp 1581365163
transform 1 0 0 0 1 4284
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_235
timestamp 1581365163
transform 1 0 0 0 1 4080
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_236
timestamp 1581365163
transform 1 0 0 0 1 3876
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_237
timestamp 1581365163
transform 1 0 0 0 1 3672
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_238
timestamp 1581365163
transform 1 0 0 0 1 3468
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_239
timestamp 1581365163
transform 1 0 0 0 1 3264
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_240
timestamp 1581365163
transform 1 0 0 0 1 3060
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_241
timestamp 1581365163
transform 1 0 0 0 1 2856
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_242
timestamp 1581365163
transform 1 0 0 0 1 2652
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_243
timestamp 1581365163
transform 1 0 0 0 1 2448
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_244
timestamp 1581365163
transform 1 0 0 0 1 2244
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_245
timestamp 1581365163
transform 1 0 0 0 1 2040
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_246
timestamp 1581365163
transform 1 0 0 0 1 1836
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_247
timestamp 1581365163
transform 1 0 0 0 1 1632
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_248
timestamp 1581365163
transform 1 0 0 0 1 1428
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_249
timestamp 1581365163
transform 1 0 0 0 1 1224
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_250
timestamp 1581365163
transform 1 0 0 0 1 1020
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_251
timestamp 1581365163
transform 1 0 0 0 1 816
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_252
timestamp 1581365163
transform 1 0 0 0 1 612
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_253
timestamp 1581365163
transform 1 0 0 0 1 408
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_254
timestamp 1581365163
transform 1 0 0 0 1 204
box 136 -79 1879 299
use sky130_rom_krom_pinv_dec_3  sky130_rom_krom_pinv_dec_3_255
timestamp 1581365163
transform 1 0 0 0 1 0
box 136 -79 1879 299
<< labels >>
rlabel locali s 1838 52104 1838 52104 4 in_0
port 2 nsew
rlabel locali s 243 52104 243 52104 4 out_0
port 3 nsew
rlabel locali s 1838 51900 1838 51900 4 in_1
port 4 nsew
rlabel locali s 243 51900 243 51900 4 out_1
port 5 nsew
rlabel locali s 1838 51696 1838 51696 4 in_2
port 6 nsew
rlabel locali s 243 51696 243 51696 4 out_2
port 7 nsew
rlabel locali s 1838 51492 1838 51492 4 in_3
port 8 nsew
rlabel locali s 243 51492 243 51492 4 out_3
port 9 nsew
rlabel locali s 1838 51288 1838 51288 4 in_4
port 10 nsew
rlabel locali s 243 51288 243 51288 4 out_4
port 11 nsew
rlabel locali s 1838 51084 1838 51084 4 in_5
port 12 nsew
rlabel locali s 243 51084 243 51084 4 out_5
port 13 nsew
rlabel locali s 1838 50880 1838 50880 4 in_6
port 14 nsew
rlabel locali s 243 50880 243 50880 4 out_6
port 15 nsew
rlabel locali s 1838 50676 1838 50676 4 in_7
port 16 nsew
rlabel locali s 243 50676 243 50676 4 out_7
port 17 nsew
rlabel locali s 1838 50472 1838 50472 4 in_8
port 18 nsew
rlabel locali s 243 50472 243 50472 4 out_8
port 19 nsew
rlabel locali s 1838 50268 1838 50268 4 in_9
port 20 nsew
rlabel locali s 243 50268 243 50268 4 out_9
port 21 nsew
rlabel locali s 1838 50064 1838 50064 4 in_10
port 22 nsew
rlabel locali s 243 50064 243 50064 4 out_10
port 23 nsew
rlabel locali s 1838 49860 1838 49860 4 in_11
port 24 nsew
rlabel locali s 243 49860 243 49860 4 out_11
port 25 nsew
rlabel locali s 1838 49656 1838 49656 4 in_12
port 26 nsew
rlabel locali s 243 49656 243 49656 4 out_12
port 27 nsew
rlabel locali s 1838 49452 1838 49452 4 in_13
port 28 nsew
rlabel locali s 243 49452 243 49452 4 out_13
port 29 nsew
rlabel locali s 1838 49248 1838 49248 4 in_14
port 30 nsew
rlabel locali s 243 49248 243 49248 4 out_14
port 31 nsew
rlabel locali s 1838 49044 1838 49044 4 in_15
port 32 nsew
rlabel locali s 243 49044 243 49044 4 out_15
port 33 nsew
rlabel locali s 1838 48840 1838 48840 4 in_16
port 34 nsew
rlabel locali s 243 48840 243 48840 4 out_16
port 35 nsew
rlabel locali s 1838 48636 1838 48636 4 in_17
port 36 nsew
rlabel locali s 243 48636 243 48636 4 out_17
port 37 nsew
rlabel locali s 1838 48432 1838 48432 4 in_18
port 38 nsew
rlabel locali s 243 48432 243 48432 4 out_18
port 39 nsew
rlabel locali s 1838 48228 1838 48228 4 in_19
port 40 nsew
rlabel locali s 243 48228 243 48228 4 out_19
port 41 nsew
rlabel locali s 1838 48024 1838 48024 4 in_20
port 42 nsew
rlabel locali s 243 48024 243 48024 4 out_20
port 43 nsew
rlabel locali s 1838 47820 1838 47820 4 in_21
port 44 nsew
rlabel locali s 243 47820 243 47820 4 out_21
port 45 nsew
rlabel locali s 1838 47616 1838 47616 4 in_22
port 46 nsew
rlabel locali s 243 47616 243 47616 4 out_22
port 47 nsew
rlabel locali s 1838 47412 1838 47412 4 in_23
port 48 nsew
rlabel locali s 243 47412 243 47412 4 out_23
port 49 nsew
rlabel locali s 1838 47208 1838 47208 4 in_24
port 50 nsew
rlabel locali s 243 47208 243 47208 4 out_24
port 51 nsew
rlabel locali s 1838 47004 1838 47004 4 in_25
port 52 nsew
rlabel locali s 243 47004 243 47004 4 out_25
port 53 nsew
rlabel locali s 1838 46800 1838 46800 4 in_26
port 54 nsew
rlabel locali s 243 46800 243 46800 4 out_26
port 55 nsew
rlabel locali s 1838 46596 1838 46596 4 in_27
port 56 nsew
rlabel locali s 243 46596 243 46596 4 out_27
port 57 nsew
rlabel locali s 1838 46392 1838 46392 4 in_28
port 58 nsew
rlabel locali s 243 46392 243 46392 4 out_28
port 59 nsew
rlabel locali s 1838 46188 1838 46188 4 in_29
port 60 nsew
rlabel locali s 243 46188 243 46188 4 out_29
port 61 nsew
rlabel locali s 1838 45984 1838 45984 4 in_30
port 62 nsew
rlabel locali s 243 45984 243 45984 4 out_30
port 63 nsew
rlabel locali s 1838 45780 1838 45780 4 in_31
port 64 nsew
rlabel locali s 243 45780 243 45780 4 out_31
port 65 nsew
rlabel locali s 1838 45576 1838 45576 4 in_32
port 66 nsew
rlabel locali s 243 45576 243 45576 4 out_32
port 67 nsew
rlabel locali s 1838 45372 1838 45372 4 in_33
port 68 nsew
rlabel locali s 243 45372 243 45372 4 out_33
port 69 nsew
rlabel locali s 1838 45168 1838 45168 4 in_34
port 70 nsew
rlabel locali s 243 45168 243 45168 4 out_34
port 71 nsew
rlabel locali s 1838 44964 1838 44964 4 in_35
port 72 nsew
rlabel locali s 243 44964 243 44964 4 out_35
port 73 nsew
rlabel locali s 1838 44760 1838 44760 4 in_36
port 74 nsew
rlabel locali s 243 44760 243 44760 4 out_36
port 75 nsew
rlabel locali s 1838 44556 1838 44556 4 in_37
port 76 nsew
rlabel locali s 243 44556 243 44556 4 out_37
port 77 nsew
rlabel locali s 1838 44352 1838 44352 4 in_38
port 78 nsew
rlabel locali s 243 44352 243 44352 4 out_38
port 79 nsew
rlabel locali s 1838 44148 1838 44148 4 in_39
port 80 nsew
rlabel locali s 243 44148 243 44148 4 out_39
port 81 nsew
rlabel locali s 1838 43944 1838 43944 4 in_40
port 82 nsew
rlabel locali s 243 43944 243 43944 4 out_40
port 83 nsew
rlabel locali s 1838 43740 1838 43740 4 in_41
port 84 nsew
rlabel locali s 243 43740 243 43740 4 out_41
port 85 nsew
rlabel locali s 1838 43536 1838 43536 4 in_42
port 86 nsew
rlabel locali s 243 43536 243 43536 4 out_42
port 87 nsew
rlabel locali s 1838 43332 1838 43332 4 in_43
port 88 nsew
rlabel locali s 243 43332 243 43332 4 out_43
port 89 nsew
rlabel locali s 1838 43128 1838 43128 4 in_44
port 90 nsew
rlabel locali s 243 43128 243 43128 4 out_44
port 91 nsew
rlabel locali s 1838 42924 1838 42924 4 in_45
port 92 nsew
rlabel locali s 243 42924 243 42924 4 out_45
port 93 nsew
rlabel locali s 1838 42720 1838 42720 4 in_46
port 94 nsew
rlabel locali s 243 42720 243 42720 4 out_46
port 95 nsew
rlabel locali s 1838 42516 1838 42516 4 in_47
port 96 nsew
rlabel locali s 243 42516 243 42516 4 out_47
port 97 nsew
rlabel locali s 1838 42312 1838 42312 4 in_48
port 98 nsew
rlabel locali s 243 42312 243 42312 4 out_48
port 99 nsew
rlabel locali s 1838 42108 1838 42108 4 in_49
port 100 nsew
rlabel locali s 243 42108 243 42108 4 out_49
port 101 nsew
rlabel locali s 1838 41904 1838 41904 4 in_50
port 102 nsew
rlabel locali s 243 41904 243 41904 4 out_50
port 103 nsew
rlabel locali s 1838 41700 1838 41700 4 in_51
port 104 nsew
rlabel locali s 243 41700 243 41700 4 out_51
port 105 nsew
rlabel locali s 1838 41496 1838 41496 4 in_52
port 106 nsew
rlabel locali s 243 41496 243 41496 4 out_52
port 107 nsew
rlabel locali s 1838 41292 1838 41292 4 in_53
port 108 nsew
rlabel locali s 243 41292 243 41292 4 out_53
port 109 nsew
rlabel locali s 1838 41088 1838 41088 4 in_54
port 110 nsew
rlabel locali s 243 41088 243 41088 4 out_54
port 111 nsew
rlabel locali s 1838 40884 1838 40884 4 in_55
port 112 nsew
rlabel locali s 243 40884 243 40884 4 out_55
port 113 nsew
rlabel locali s 1838 40680 1838 40680 4 in_56
port 114 nsew
rlabel locali s 243 40680 243 40680 4 out_56
port 115 nsew
rlabel locali s 1838 40476 1838 40476 4 in_57
port 116 nsew
rlabel locali s 243 40476 243 40476 4 out_57
port 117 nsew
rlabel locali s 1838 40272 1838 40272 4 in_58
port 118 nsew
rlabel locali s 243 40272 243 40272 4 out_58
port 119 nsew
rlabel locali s 1838 40068 1838 40068 4 in_59
port 120 nsew
rlabel locali s 243 40068 243 40068 4 out_59
port 121 nsew
rlabel locali s 1838 39864 1838 39864 4 in_60
port 122 nsew
rlabel locali s 243 39864 243 39864 4 out_60
port 123 nsew
rlabel locali s 1838 39660 1838 39660 4 in_61
port 124 nsew
rlabel locali s 243 39660 243 39660 4 out_61
port 125 nsew
rlabel locali s 1838 39456 1838 39456 4 in_62
port 126 nsew
rlabel locali s 243 39456 243 39456 4 out_62
port 127 nsew
rlabel locali s 1838 39252 1838 39252 4 in_63
port 128 nsew
rlabel locali s 243 39252 243 39252 4 out_63
port 129 nsew
rlabel locali s 1838 39048 1838 39048 4 in_64
port 130 nsew
rlabel locali s 243 39048 243 39048 4 out_64
port 131 nsew
rlabel locali s 1838 38844 1838 38844 4 in_65
port 132 nsew
rlabel locali s 243 38844 243 38844 4 out_65
port 133 nsew
rlabel locali s 1838 38640 1838 38640 4 in_66
port 134 nsew
rlabel locali s 243 38640 243 38640 4 out_66
port 135 nsew
rlabel locali s 1838 38436 1838 38436 4 in_67
port 136 nsew
rlabel locali s 243 38436 243 38436 4 out_67
port 137 nsew
rlabel locali s 1838 38232 1838 38232 4 in_68
port 138 nsew
rlabel locali s 243 38232 243 38232 4 out_68
port 139 nsew
rlabel locali s 1838 38028 1838 38028 4 in_69
port 140 nsew
rlabel locali s 243 38028 243 38028 4 out_69
port 141 nsew
rlabel locali s 1838 37824 1838 37824 4 in_70
port 142 nsew
rlabel locali s 243 37824 243 37824 4 out_70
port 143 nsew
rlabel locali s 1838 37620 1838 37620 4 in_71
port 144 nsew
rlabel locali s 243 37620 243 37620 4 out_71
port 145 nsew
rlabel locali s 1838 37416 1838 37416 4 in_72
port 146 nsew
rlabel locali s 243 37416 243 37416 4 out_72
port 147 nsew
rlabel locali s 1838 37212 1838 37212 4 in_73
port 148 nsew
rlabel locali s 243 37212 243 37212 4 out_73
port 149 nsew
rlabel locali s 1838 37008 1838 37008 4 in_74
port 150 nsew
rlabel locali s 243 37008 243 37008 4 out_74
port 151 nsew
rlabel locali s 1838 36804 1838 36804 4 in_75
port 152 nsew
rlabel locali s 243 36804 243 36804 4 out_75
port 153 nsew
rlabel locali s 1838 36600 1838 36600 4 in_76
port 154 nsew
rlabel locali s 243 36600 243 36600 4 out_76
port 155 nsew
rlabel locali s 1838 36396 1838 36396 4 in_77
port 156 nsew
rlabel locali s 243 36396 243 36396 4 out_77
port 157 nsew
rlabel locali s 1838 36192 1838 36192 4 in_78
port 158 nsew
rlabel locali s 243 36192 243 36192 4 out_78
port 159 nsew
rlabel locali s 1838 35988 1838 35988 4 in_79
port 160 nsew
rlabel locali s 243 35988 243 35988 4 out_79
port 161 nsew
rlabel locali s 1838 35784 1838 35784 4 in_80
port 162 nsew
rlabel locali s 243 35784 243 35784 4 out_80
port 163 nsew
rlabel locali s 1838 35580 1838 35580 4 in_81
port 164 nsew
rlabel locali s 243 35580 243 35580 4 out_81
port 165 nsew
rlabel locali s 1838 35376 1838 35376 4 in_82
port 166 nsew
rlabel locali s 243 35376 243 35376 4 out_82
port 167 nsew
rlabel locali s 1838 35172 1838 35172 4 in_83
port 168 nsew
rlabel locali s 243 35172 243 35172 4 out_83
port 169 nsew
rlabel locali s 1838 34968 1838 34968 4 in_84
port 170 nsew
rlabel locali s 243 34968 243 34968 4 out_84
port 171 nsew
rlabel locali s 1838 34764 1838 34764 4 in_85
port 172 nsew
rlabel locali s 243 34764 243 34764 4 out_85
port 173 nsew
rlabel locali s 1838 34560 1838 34560 4 in_86
port 174 nsew
rlabel locali s 243 34560 243 34560 4 out_86
port 175 nsew
rlabel locali s 1838 34356 1838 34356 4 in_87
port 176 nsew
rlabel locali s 243 34356 243 34356 4 out_87
port 177 nsew
rlabel locali s 1838 34152 1838 34152 4 in_88
port 178 nsew
rlabel locali s 243 34152 243 34152 4 out_88
port 179 nsew
rlabel locali s 1838 33948 1838 33948 4 in_89
port 180 nsew
rlabel locali s 243 33948 243 33948 4 out_89
port 181 nsew
rlabel locali s 1838 33744 1838 33744 4 in_90
port 182 nsew
rlabel locali s 243 33744 243 33744 4 out_90
port 183 nsew
rlabel locali s 1838 33540 1838 33540 4 in_91
port 184 nsew
rlabel locali s 243 33540 243 33540 4 out_91
port 185 nsew
rlabel locali s 1838 33336 1838 33336 4 in_92
port 186 nsew
rlabel locali s 243 33336 243 33336 4 out_92
port 187 nsew
rlabel locali s 1838 33132 1838 33132 4 in_93
port 188 nsew
rlabel locali s 243 33132 243 33132 4 out_93
port 189 nsew
rlabel locali s 1838 32928 1838 32928 4 in_94
port 190 nsew
rlabel locali s 243 32928 243 32928 4 out_94
port 191 nsew
rlabel locali s 1838 32724 1838 32724 4 in_95
port 192 nsew
rlabel locali s 243 32724 243 32724 4 out_95
port 193 nsew
rlabel locali s 1838 32520 1838 32520 4 in_96
port 194 nsew
rlabel locali s 243 32520 243 32520 4 out_96
port 195 nsew
rlabel locali s 1838 32316 1838 32316 4 in_97
port 196 nsew
rlabel locali s 243 32316 243 32316 4 out_97
port 197 nsew
rlabel locali s 1838 32112 1838 32112 4 in_98
port 198 nsew
rlabel locali s 243 32112 243 32112 4 out_98
port 199 nsew
rlabel locali s 1838 31908 1838 31908 4 in_99
port 200 nsew
rlabel locali s 243 31908 243 31908 4 out_99
port 201 nsew
rlabel locali s 1838 31704 1838 31704 4 in_100
port 202 nsew
rlabel locali s 243 31704 243 31704 4 out_100
port 203 nsew
rlabel locali s 1838 31500 1838 31500 4 in_101
port 204 nsew
rlabel locali s 243 31500 243 31500 4 out_101
port 205 nsew
rlabel locali s 1838 31296 1838 31296 4 in_102
port 206 nsew
rlabel locali s 243 31296 243 31296 4 out_102
port 207 nsew
rlabel locali s 1838 31092 1838 31092 4 in_103
port 208 nsew
rlabel locali s 243 31092 243 31092 4 out_103
port 209 nsew
rlabel locali s 1838 30888 1838 30888 4 in_104
port 210 nsew
rlabel locali s 243 30888 243 30888 4 out_104
port 211 nsew
rlabel locali s 1838 30684 1838 30684 4 in_105
port 212 nsew
rlabel locali s 243 30684 243 30684 4 out_105
port 213 nsew
rlabel locali s 1838 30480 1838 30480 4 in_106
port 214 nsew
rlabel locali s 243 30480 243 30480 4 out_106
port 215 nsew
rlabel locali s 1838 30276 1838 30276 4 in_107
port 216 nsew
rlabel locali s 243 30276 243 30276 4 out_107
port 217 nsew
rlabel locali s 1838 30072 1838 30072 4 in_108
port 218 nsew
rlabel locali s 243 30072 243 30072 4 out_108
port 219 nsew
rlabel locali s 1838 29868 1838 29868 4 in_109
port 220 nsew
rlabel locali s 243 29868 243 29868 4 out_109
port 221 nsew
rlabel locali s 1838 29664 1838 29664 4 in_110
port 222 nsew
rlabel locali s 243 29664 243 29664 4 out_110
port 223 nsew
rlabel locali s 1838 29460 1838 29460 4 in_111
port 224 nsew
rlabel locali s 243 29460 243 29460 4 out_111
port 225 nsew
rlabel locali s 1838 29256 1838 29256 4 in_112
port 226 nsew
rlabel locali s 243 29256 243 29256 4 out_112
port 227 nsew
rlabel locali s 1838 29052 1838 29052 4 in_113
port 228 nsew
rlabel locali s 243 29052 243 29052 4 out_113
port 229 nsew
rlabel locali s 1838 28848 1838 28848 4 in_114
port 230 nsew
rlabel locali s 243 28848 243 28848 4 out_114
port 231 nsew
rlabel locali s 1838 28644 1838 28644 4 in_115
port 232 nsew
rlabel locali s 243 28644 243 28644 4 out_115
port 233 nsew
rlabel locali s 1838 28440 1838 28440 4 in_116
port 234 nsew
rlabel locali s 243 28440 243 28440 4 out_116
port 235 nsew
rlabel locali s 1838 28236 1838 28236 4 in_117
port 236 nsew
rlabel locali s 243 28236 243 28236 4 out_117
port 237 nsew
rlabel locali s 1838 28032 1838 28032 4 in_118
port 238 nsew
rlabel locali s 243 28032 243 28032 4 out_118
port 239 nsew
rlabel locali s 1838 27828 1838 27828 4 in_119
port 240 nsew
rlabel locali s 243 27828 243 27828 4 out_119
port 241 nsew
rlabel locali s 1838 27624 1838 27624 4 in_120
port 242 nsew
rlabel locali s 243 27624 243 27624 4 out_120
port 243 nsew
rlabel locali s 1838 27420 1838 27420 4 in_121
port 244 nsew
rlabel locali s 243 27420 243 27420 4 out_121
port 245 nsew
rlabel locali s 1838 27216 1838 27216 4 in_122
port 246 nsew
rlabel locali s 243 27216 243 27216 4 out_122
port 247 nsew
rlabel locali s 1838 27012 1838 27012 4 in_123
port 248 nsew
rlabel locali s 243 27012 243 27012 4 out_123
port 249 nsew
rlabel locali s 1838 26808 1838 26808 4 in_124
port 250 nsew
rlabel locali s 243 26808 243 26808 4 out_124
port 251 nsew
rlabel locali s 1838 26604 1838 26604 4 in_125
port 252 nsew
rlabel locali s 243 26604 243 26604 4 out_125
port 253 nsew
rlabel locali s 1838 26400 1838 26400 4 in_126
port 254 nsew
rlabel locali s 243 26400 243 26400 4 out_126
port 255 nsew
rlabel locali s 1838 26196 1838 26196 4 in_127
port 256 nsew
rlabel locali s 243 26196 243 26196 4 out_127
port 257 nsew
rlabel locali s 1838 25992 1838 25992 4 in_128
port 258 nsew
rlabel locali s 243 25992 243 25992 4 out_128
port 259 nsew
rlabel locali s 1838 25788 1838 25788 4 in_129
port 260 nsew
rlabel locali s 243 25788 243 25788 4 out_129
port 261 nsew
rlabel locali s 1838 25584 1838 25584 4 in_130
port 262 nsew
rlabel locali s 243 25584 243 25584 4 out_130
port 263 nsew
rlabel locali s 1838 25380 1838 25380 4 in_131
port 264 nsew
rlabel locali s 243 25380 243 25380 4 out_131
port 265 nsew
rlabel locali s 1838 25176 1838 25176 4 in_132
port 266 nsew
rlabel locali s 243 25176 243 25176 4 out_132
port 267 nsew
rlabel locali s 1838 24972 1838 24972 4 in_133
port 268 nsew
rlabel locali s 243 24972 243 24972 4 out_133
port 269 nsew
rlabel locali s 1838 24768 1838 24768 4 in_134
port 270 nsew
rlabel locali s 243 24768 243 24768 4 out_134
port 271 nsew
rlabel locali s 1838 24564 1838 24564 4 in_135
port 272 nsew
rlabel locali s 243 24564 243 24564 4 out_135
port 273 nsew
rlabel locali s 1838 24360 1838 24360 4 in_136
port 274 nsew
rlabel locali s 243 24360 243 24360 4 out_136
port 275 nsew
rlabel locali s 1838 24156 1838 24156 4 in_137
port 276 nsew
rlabel locali s 243 24156 243 24156 4 out_137
port 277 nsew
rlabel locali s 1838 23952 1838 23952 4 in_138
port 278 nsew
rlabel locali s 243 23952 243 23952 4 out_138
port 279 nsew
rlabel locali s 1838 23748 1838 23748 4 in_139
port 280 nsew
rlabel locali s 243 23748 243 23748 4 out_139
port 281 nsew
rlabel locali s 1838 23544 1838 23544 4 in_140
port 282 nsew
rlabel locali s 243 23544 243 23544 4 out_140
port 283 nsew
rlabel locali s 1838 23340 1838 23340 4 in_141
port 284 nsew
rlabel locali s 243 23340 243 23340 4 out_141
port 285 nsew
rlabel locali s 1838 23136 1838 23136 4 in_142
port 286 nsew
rlabel locali s 243 23136 243 23136 4 out_142
port 287 nsew
rlabel locali s 1838 22932 1838 22932 4 in_143
port 288 nsew
rlabel locali s 243 22932 243 22932 4 out_143
port 289 nsew
rlabel locali s 1838 22728 1838 22728 4 in_144
port 290 nsew
rlabel locali s 243 22728 243 22728 4 out_144
port 291 nsew
rlabel locali s 1838 22524 1838 22524 4 in_145
port 292 nsew
rlabel locali s 243 22524 243 22524 4 out_145
port 293 nsew
rlabel locali s 1838 22320 1838 22320 4 in_146
port 294 nsew
rlabel locali s 243 22320 243 22320 4 out_146
port 295 nsew
rlabel locali s 1838 22116 1838 22116 4 in_147
port 296 nsew
rlabel locali s 243 22116 243 22116 4 out_147
port 297 nsew
rlabel locali s 1838 21912 1838 21912 4 in_148
port 298 nsew
rlabel locali s 243 21912 243 21912 4 out_148
port 299 nsew
rlabel locali s 1838 21708 1838 21708 4 in_149
port 300 nsew
rlabel locali s 243 21708 243 21708 4 out_149
port 301 nsew
rlabel locali s 1838 21504 1838 21504 4 in_150
port 302 nsew
rlabel locali s 243 21504 243 21504 4 out_150
port 303 nsew
rlabel locali s 1838 21300 1838 21300 4 in_151
port 304 nsew
rlabel locali s 243 21300 243 21300 4 out_151
port 305 nsew
rlabel locali s 1838 21096 1838 21096 4 in_152
port 306 nsew
rlabel locali s 243 21096 243 21096 4 out_152
port 307 nsew
rlabel locali s 1838 20892 1838 20892 4 in_153
port 308 nsew
rlabel locali s 243 20892 243 20892 4 out_153
port 309 nsew
rlabel locali s 1838 20688 1838 20688 4 in_154
port 310 nsew
rlabel locali s 243 20688 243 20688 4 out_154
port 311 nsew
rlabel locali s 1838 20484 1838 20484 4 in_155
port 312 nsew
rlabel locali s 243 20484 243 20484 4 out_155
port 313 nsew
rlabel locali s 1838 20280 1838 20280 4 in_156
port 314 nsew
rlabel locali s 243 20280 243 20280 4 out_156
port 315 nsew
rlabel locali s 1838 20076 1838 20076 4 in_157
port 316 nsew
rlabel locali s 243 20076 243 20076 4 out_157
port 317 nsew
rlabel locali s 1838 19872 1838 19872 4 in_158
port 318 nsew
rlabel locali s 243 19872 243 19872 4 out_158
port 319 nsew
rlabel locali s 1838 19668 1838 19668 4 in_159
port 320 nsew
rlabel locali s 243 19668 243 19668 4 out_159
port 321 nsew
rlabel locali s 1838 19464 1838 19464 4 in_160
port 322 nsew
rlabel locali s 243 19464 243 19464 4 out_160
port 323 nsew
rlabel locali s 1838 19260 1838 19260 4 in_161
port 324 nsew
rlabel locali s 243 19260 243 19260 4 out_161
port 325 nsew
rlabel locali s 1838 19056 1838 19056 4 in_162
port 326 nsew
rlabel locali s 243 19056 243 19056 4 out_162
port 327 nsew
rlabel locali s 1838 18852 1838 18852 4 in_163
port 328 nsew
rlabel locali s 243 18852 243 18852 4 out_163
port 329 nsew
rlabel locali s 1838 18648 1838 18648 4 in_164
port 330 nsew
rlabel locali s 243 18648 243 18648 4 out_164
port 331 nsew
rlabel locali s 1838 18444 1838 18444 4 in_165
port 332 nsew
rlabel locali s 243 18444 243 18444 4 out_165
port 333 nsew
rlabel locali s 1838 18240 1838 18240 4 in_166
port 334 nsew
rlabel locali s 243 18240 243 18240 4 out_166
port 335 nsew
rlabel locali s 1838 18036 1838 18036 4 in_167
port 336 nsew
rlabel locali s 243 18036 243 18036 4 out_167
port 337 nsew
rlabel locali s 1838 17832 1838 17832 4 in_168
port 338 nsew
rlabel locali s 243 17832 243 17832 4 out_168
port 339 nsew
rlabel locali s 1838 17628 1838 17628 4 in_169
port 340 nsew
rlabel locali s 243 17628 243 17628 4 out_169
port 341 nsew
rlabel locali s 1838 17424 1838 17424 4 in_170
port 342 nsew
rlabel locali s 243 17424 243 17424 4 out_170
port 343 nsew
rlabel locali s 1838 17220 1838 17220 4 in_171
port 344 nsew
rlabel locali s 243 17220 243 17220 4 out_171
port 345 nsew
rlabel locali s 1838 17016 1838 17016 4 in_172
port 346 nsew
rlabel locali s 243 17016 243 17016 4 out_172
port 347 nsew
rlabel locali s 1838 16812 1838 16812 4 in_173
port 348 nsew
rlabel locali s 243 16812 243 16812 4 out_173
port 349 nsew
rlabel locali s 1838 16608 1838 16608 4 in_174
port 350 nsew
rlabel locali s 243 16608 243 16608 4 out_174
port 351 nsew
rlabel locali s 1838 16404 1838 16404 4 in_175
port 352 nsew
rlabel locali s 243 16404 243 16404 4 out_175
port 353 nsew
rlabel locali s 1838 16200 1838 16200 4 in_176
port 354 nsew
rlabel locali s 243 16200 243 16200 4 out_176
port 355 nsew
rlabel locali s 1838 15996 1838 15996 4 in_177
port 356 nsew
rlabel locali s 243 15996 243 15996 4 out_177
port 357 nsew
rlabel locali s 1838 15792 1838 15792 4 in_178
port 358 nsew
rlabel locali s 243 15792 243 15792 4 out_178
port 359 nsew
rlabel locali s 1838 15588 1838 15588 4 in_179
port 360 nsew
rlabel locali s 243 15588 243 15588 4 out_179
port 361 nsew
rlabel locali s 1838 15384 1838 15384 4 in_180
port 362 nsew
rlabel locali s 243 15384 243 15384 4 out_180
port 363 nsew
rlabel locali s 1838 15180 1838 15180 4 in_181
port 364 nsew
rlabel locali s 243 15180 243 15180 4 out_181
port 365 nsew
rlabel locali s 1838 14976 1838 14976 4 in_182
port 366 nsew
rlabel locali s 243 14976 243 14976 4 out_182
port 367 nsew
rlabel locali s 1838 14772 1838 14772 4 in_183
port 368 nsew
rlabel locali s 243 14772 243 14772 4 out_183
port 369 nsew
rlabel locali s 1838 14568 1838 14568 4 in_184
port 370 nsew
rlabel locali s 243 14568 243 14568 4 out_184
port 371 nsew
rlabel locali s 1838 14364 1838 14364 4 in_185
port 372 nsew
rlabel locali s 243 14364 243 14364 4 out_185
port 373 nsew
rlabel locali s 1838 14160 1838 14160 4 in_186
port 374 nsew
rlabel locali s 243 14160 243 14160 4 out_186
port 375 nsew
rlabel locali s 1838 13956 1838 13956 4 in_187
port 376 nsew
rlabel locali s 243 13956 243 13956 4 out_187
port 377 nsew
rlabel locali s 1838 13752 1838 13752 4 in_188
port 378 nsew
rlabel locali s 243 13752 243 13752 4 out_188
port 379 nsew
rlabel locali s 1838 13548 1838 13548 4 in_189
port 380 nsew
rlabel locali s 243 13548 243 13548 4 out_189
port 381 nsew
rlabel locali s 1838 13344 1838 13344 4 in_190
port 382 nsew
rlabel locali s 243 13344 243 13344 4 out_190
port 383 nsew
rlabel locali s 1838 13140 1838 13140 4 in_191
port 384 nsew
rlabel locali s 243 13140 243 13140 4 out_191
port 385 nsew
rlabel locali s 1838 12936 1838 12936 4 in_192
port 386 nsew
rlabel locali s 243 12936 243 12936 4 out_192
port 387 nsew
rlabel locali s 1838 12732 1838 12732 4 in_193
port 388 nsew
rlabel locali s 243 12732 243 12732 4 out_193
port 389 nsew
rlabel locali s 1838 12528 1838 12528 4 in_194
port 390 nsew
rlabel locali s 243 12528 243 12528 4 out_194
port 391 nsew
rlabel locali s 1838 12324 1838 12324 4 in_195
port 392 nsew
rlabel locali s 243 12324 243 12324 4 out_195
port 393 nsew
rlabel locali s 1838 12120 1838 12120 4 in_196
port 394 nsew
rlabel locali s 243 12120 243 12120 4 out_196
port 395 nsew
rlabel locali s 1838 11916 1838 11916 4 in_197
port 396 nsew
rlabel locali s 243 11916 243 11916 4 out_197
port 397 nsew
rlabel locali s 1838 11712 1838 11712 4 in_198
port 398 nsew
rlabel locali s 243 11712 243 11712 4 out_198
port 399 nsew
rlabel locali s 1838 11508 1838 11508 4 in_199
port 400 nsew
rlabel locali s 243 11508 243 11508 4 out_199
port 401 nsew
rlabel locali s 1838 11304 1838 11304 4 in_200
port 402 nsew
rlabel locali s 243 11304 243 11304 4 out_200
port 403 nsew
rlabel locali s 1838 11100 1838 11100 4 in_201
port 404 nsew
rlabel locali s 243 11100 243 11100 4 out_201
port 405 nsew
rlabel locali s 1838 10896 1838 10896 4 in_202
port 406 nsew
rlabel locali s 243 10896 243 10896 4 out_202
port 407 nsew
rlabel locali s 1838 10692 1838 10692 4 in_203
port 408 nsew
rlabel locali s 243 10692 243 10692 4 out_203
port 409 nsew
rlabel locali s 1838 10488 1838 10488 4 in_204
port 410 nsew
rlabel locali s 243 10488 243 10488 4 out_204
port 411 nsew
rlabel locali s 1838 10284 1838 10284 4 in_205
port 412 nsew
rlabel locali s 243 10284 243 10284 4 out_205
port 413 nsew
rlabel locali s 1838 10080 1838 10080 4 in_206
port 414 nsew
rlabel locali s 243 10080 243 10080 4 out_206
port 415 nsew
rlabel locali s 1838 9876 1838 9876 4 in_207
port 416 nsew
rlabel locali s 243 9876 243 9876 4 out_207
port 417 nsew
rlabel locali s 1838 9672 1838 9672 4 in_208
port 418 nsew
rlabel locali s 243 9672 243 9672 4 out_208
port 419 nsew
rlabel locali s 1838 9468 1838 9468 4 in_209
port 420 nsew
rlabel locali s 243 9468 243 9468 4 out_209
port 421 nsew
rlabel locali s 1838 9264 1838 9264 4 in_210
port 422 nsew
rlabel locali s 243 9264 243 9264 4 out_210
port 423 nsew
rlabel locali s 1838 9060 1838 9060 4 in_211
port 424 nsew
rlabel locali s 243 9060 243 9060 4 out_211
port 425 nsew
rlabel locali s 1838 8856 1838 8856 4 in_212
port 426 nsew
rlabel locali s 243 8856 243 8856 4 out_212
port 427 nsew
rlabel locali s 1838 8652 1838 8652 4 in_213
port 428 nsew
rlabel locali s 243 8652 243 8652 4 out_213
port 429 nsew
rlabel locali s 1838 8448 1838 8448 4 in_214
port 430 nsew
rlabel locali s 243 8448 243 8448 4 out_214
port 431 nsew
rlabel locali s 1838 8244 1838 8244 4 in_215
port 432 nsew
rlabel locali s 243 8244 243 8244 4 out_215
port 433 nsew
rlabel locali s 1838 8040 1838 8040 4 in_216
port 434 nsew
rlabel locali s 243 8040 243 8040 4 out_216
port 435 nsew
rlabel locali s 1838 7836 1838 7836 4 in_217
port 436 nsew
rlabel locali s 243 7836 243 7836 4 out_217
port 437 nsew
rlabel locali s 1838 7632 1838 7632 4 in_218
port 438 nsew
rlabel locali s 243 7632 243 7632 4 out_218
port 439 nsew
rlabel locali s 1838 7428 1838 7428 4 in_219
port 440 nsew
rlabel locali s 243 7428 243 7428 4 out_219
port 441 nsew
rlabel locali s 1838 7224 1838 7224 4 in_220
port 442 nsew
rlabel locali s 243 7224 243 7224 4 out_220
port 443 nsew
rlabel locali s 1838 7020 1838 7020 4 in_221
port 444 nsew
rlabel locali s 243 7020 243 7020 4 out_221
port 445 nsew
rlabel locali s 1838 6816 1838 6816 4 in_222
port 446 nsew
rlabel locali s 243 6816 243 6816 4 out_222
port 447 nsew
rlabel locali s 1838 6612 1838 6612 4 in_223
port 448 nsew
rlabel locali s 243 6612 243 6612 4 out_223
port 449 nsew
rlabel locali s 1838 6408 1838 6408 4 in_224
port 450 nsew
rlabel locali s 243 6408 243 6408 4 out_224
port 451 nsew
rlabel locali s 1838 6204 1838 6204 4 in_225
port 452 nsew
rlabel locali s 243 6204 243 6204 4 out_225
port 453 nsew
rlabel locali s 1838 6000 1838 6000 4 in_226
port 454 nsew
rlabel locali s 243 6000 243 6000 4 out_226
port 455 nsew
rlabel locali s 1838 5796 1838 5796 4 in_227
port 456 nsew
rlabel locali s 243 5796 243 5796 4 out_227
port 457 nsew
rlabel locali s 1838 5592 1838 5592 4 in_228
port 458 nsew
rlabel locali s 243 5592 243 5592 4 out_228
port 459 nsew
rlabel locali s 1838 5388 1838 5388 4 in_229
port 460 nsew
rlabel locali s 243 5388 243 5388 4 out_229
port 461 nsew
rlabel locali s 1838 5184 1838 5184 4 in_230
port 462 nsew
rlabel locali s 243 5184 243 5184 4 out_230
port 463 nsew
rlabel locali s 1838 4980 1838 4980 4 in_231
port 464 nsew
rlabel locali s 243 4980 243 4980 4 out_231
port 465 nsew
rlabel locali s 1838 4776 1838 4776 4 in_232
port 466 nsew
rlabel locali s 243 4776 243 4776 4 out_232
port 467 nsew
rlabel locali s 1838 4572 1838 4572 4 in_233
port 468 nsew
rlabel locali s 243 4572 243 4572 4 out_233
port 469 nsew
rlabel locali s 1838 4368 1838 4368 4 in_234
port 470 nsew
rlabel locali s 243 4368 243 4368 4 out_234
port 471 nsew
rlabel locali s 1838 4164 1838 4164 4 in_235
port 472 nsew
rlabel locali s 243 4164 243 4164 4 out_235
port 473 nsew
rlabel locali s 1838 3960 1838 3960 4 in_236
port 474 nsew
rlabel locali s 243 3960 243 3960 4 out_236
port 475 nsew
rlabel locali s 1838 3756 1838 3756 4 in_237
port 476 nsew
rlabel locali s 243 3756 243 3756 4 out_237
port 477 nsew
rlabel locali s 1838 3552 1838 3552 4 in_238
port 478 nsew
rlabel locali s 243 3552 243 3552 4 out_238
port 479 nsew
rlabel locali s 1838 3348 1838 3348 4 in_239
port 480 nsew
rlabel locali s 243 3348 243 3348 4 out_239
port 481 nsew
rlabel locali s 1838 3144 1838 3144 4 in_240
port 482 nsew
rlabel locali s 243 3144 243 3144 4 out_240
port 483 nsew
rlabel locali s 1838 2940 1838 2940 4 in_241
port 484 nsew
rlabel locali s 243 2940 243 2940 4 out_241
port 485 nsew
rlabel locali s 1838 2736 1838 2736 4 in_242
port 486 nsew
rlabel locali s 243 2736 243 2736 4 out_242
port 487 nsew
rlabel locali s 1838 2532 1838 2532 4 in_243
port 488 nsew
rlabel locali s 243 2532 243 2532 4 out_243
port 489 nsew
rlabel locali s 1838 2328 1838 2328 4 in_244
port 490 nsew
rlabel locali s 243 2328 243 2328 4 out_244
port 491 nsew
rlabel locali s 1838 2124 1838 2124 4 in_245
port 492 nsew
rlabel locali s 243 2124 243 2124 4 out_245
port 493 nsew
rlabel locali s 1838 1920 1838 1920 4 in_246
port 494 nsew
rlabel locali s 243 1920 243 1920 4 out_246
port 495 nsew
rlabel locali s 1838 1716 1838 1716 4 in_247
port 496 nsew
rlabel locali s 243 1716 243 1716 4 out_247
port 497 nsew
rlabel locali s 1838 1512 1838 1512 4 in_248
port 498 nsew
rlabel locali s 243 1512 243 1512 4 out_248
port 499 nsew
rlabel locali s 1838 1308 1838 1308 4 in_249
port 500 nsew
rlabel locali s 243 1308 243 1308 4 out_249
port 501 nsew
rlabel locali s 1838 1104 1838 1104 4 in_250
port 502 nsew
rlabel locali s 243 1104 243 1104 4 out_250
port 503 nsew
rlabel locali s 1838 900 1838 900 4 in_251
port 504 nsew
rlabel locali s 243 900 243 900 4 out_251
port 505 nsew
rlabel locali s 1838 696 1838 696 4 in_252
port 506 nsew
rlabel locali s 243 696 243 696 4 out_252
port 507 nsew
rlabel locali s 1838 492 1838 492 4 in_253
port 508 nsew
rlabel locali s 243 492 243 492 4 out_253
port 509 nsew
rlabel locali s 1838 288 1838 288 4 in_254
port 510 nsew
rlabel locali s 243 288 243 288 4 out_254
port 511 nsew
rlabel locali s 1838 84 1838 84 4 in_255
port 512 nsew
rlabel locali s 243 84 243 84 4 out_255
port 513 nsew
rlabel metal1 s 316 -14 344 14 4 gnd
port 515 nsew
rlabel metal1 s 316 52210 344 52238 4 gnd
port 515 nsew
rlabel metal1 s 1232 52210 1260 52238 4 vdd
port 517 nsew
rlabel metal1 s 1232 -14 1260 14 4 vdd
port 517 nsew
<< properties >>
string FIXED_BBOX 0 0 1782 52224
<< end >>
