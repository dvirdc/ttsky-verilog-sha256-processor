magic
tech sky130A
magscale 1 2
timestamp 1581320207
<< checkpaint >>
rect -1296 -1277 3892 3946
<< nwell >>
rect -36 1261 2632 2686
<< locali >>
rect 0 2611 2596 2645
rect 64 1244 98 1310
rect 1395 1298 1769 1332
rect 2087 1298 2121 1332
rect 196 1260 449 1294
rect 564 1260 817 1294
rect 919 1182 953 1277
rect 919 1148 1293 1182
rect 1395 1165 1429 1298
rect 0 -17 2596 17
use sky130_rom_krom_pinv  sky130_rom_krom_pinv_0
timestamp 1581320207
transform 1 0 368 0 1 0
box -36 -17 404 2686
use sky130_rom_krom_pinv  sky130_rom_krom_pinv_1
timestamp 1581320207
transform 1 0 0 0 1 0
box -36 -17 404 2686
use sky130_rom_krom_pinv_3  sky130_rom_krom_pinv_3_0
timestamp 1581320207
transform 1 0 736 0 1 0
box -36 -17 512 2686
use sky130_rom_krom_pinv_4  sky130_rom_krom_pinv_4_0
timestamp 1581320207
transform 1 0 1212 0 1 0
box -36 -17 512 2686
use sky130_rom_krom_pinv_5  sky130_rom_krom_pinv_5_0
timestamp 1581320207
transform 1 0 1688 0 1 0
box -36 -17 944 2686
<< labels >>
rlabel locali s 2104 1315 2104 1315 4 Z
port 1 nsew
rlabel locali s 81 1277 81 1277 4 A
port 2 nsew
rlabel locali s 1298 0 1298 0 4 gnd
port 3 nsew
rlabel locali s 1298 2628 1298 2628 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2596 2628
<< end >>
