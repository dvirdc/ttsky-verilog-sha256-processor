magic
tech sky130A
magscale 1 2
timestamp 1581449089
<< checkpaint >>
rect -1216 -1310 3060 11211
<< nwell >>
rect 1162 9498 1330 9666
rect 1162 9190 1330 9358
rect 1162 8882 1330 9050
rect 1162 8574 1330 8742
rect 1162 8266 1330 8434
rect 1162 7958 1330 8126
rect 1162 7650 1330 7818
rect 1162 7342 1330 7510
rect 1162 7034 1330 7202
rect 1162 6726 1330 6894
rect 1162 6418 1330 6586
rect 1162 6110 1330 6278
rect 1162 5802 1330 5970
rect 1162 5494 1330 5662
rect 1162 5186 1330 5354
rect 1162 4878 1330 5046
rect 1162 4570 1330 4738
rect 1162 4262 1330 4430
rect 1162 3954 1330 4122
rect 1162 3646 1330 3814
rect 1162 3338 1330 3506
rect 1162 3030 1330 3198
rect 1162 2722 1330 2890
rect 1162 2414 1330 2582
rect 1162 2106 1330 2274
rect 1162 1798 1330 1966
rect 1162 1490 1330 1658
rect 1162 1182 1330 1350
rect 1162 874 1330 1042
rect 1162 566 1330 734
rect 1162 258 1330 426
rect 1162 -50 1330 118
<< pwell >>
rect 263 9531 397 9633
rect 263 9223 397 9325
rect 263 8915 397 9017
rect 263 8607 397 8709
rect 263 8299 397 8401
rect 263 7991 397 8093
rect 263 7683 397 7785
rect 263 7375 397 7477
rect 263 7067 397 7169
rect 263 6759 397 6861
rect 263 6451 397 6553
rect 263 6143 397 6245
rect 263 5835 397 5937
rect 263 5527 397 5629
rect 263 5219 397 5321
rect 263 4911 397 5013
rect 263 4603 397 4705
rect 263 4295 397 4397
rect 263 3987 397 4089
rect 263 3679 397 3781
rect 263 3371 397 3473
rect 263 3063 397 3165
rect 263 2755 397 2857
rect 263 2447 397 2549
rect 263 2139 397 2241
rect 263 1831 397 1933
rect 263 1523 397 1625
rect 263 1215 397 1317
rect 263 907 397 1009
rect 263 599 397 701
rect 263 291 397 393
rect 263 -17 397 85
<< psubdiff >>
rect 289 9599 371 9607
rect 289 9565 313 9599
rect 347 9565 371 9599
rect 289 9557 371 9565
rect 289 9291 371 9299
rect 289 9257 313 9291
rect 347 9257 371 9291
rect 289 9249 371 9257
rect 289 8983 371 8991
rect 289 8949 313 8983
rect 347 8949 371 8983
rect 289 8941 371 8949
rect 289 8675 371 8683
rect 289 8641 313 8675
rect 347 8641 371 8675
rect 289 8633 371 8641
rect 289 8367 371 8375
rect 289 8333 313 8367
rect 347 8333 371 8367
rect 289 8325 371 8333
rect 289 8059 371 8067
rect 289 8025 313 8059
rect 347 8025 371 8059
rect 289 8017 371 8025
rect 289 7751 371 7759
rect 289 7717 313 7751
rect 347 7717 371 7751
rect 289 7709 371 7717
rect 289 7443 371 7451
rect 289 7409 313 7443
rect 347 7409 371 7443
rect 289 7401 371 7409
rect 289 7135 371 7143
rect 289 7101 313 7135
rect 347 7101 371 7135
rect 289 7093 371 7101
rect 289 6827 371 6835
rect 289 6793 313 6827
rect 347 6793 371 6827
rect 289 6785 371 6793
rect 289 6519 371 6527
rect 289 6485 313 6519
rect 347 6485 371 6519
rect 289 6477 371 6485
rect 289 6211 371 6219
rect 289 6177 313 6211
rect 347 6177 371 6211
rect 289 6169 371 6177
rect 289 5903 371 5911
rect 289 5869 313 5903
rect 347 5869 371 5903
rect 289 5861 371 5869
rect 289 5595 371 5603
rect 289 5561 313 5595
rect 347 5561 371 5595
rect 289 5553 371 5561
rect 289 5287 371 5295
rect 289 5253 313 5287
rect 347 5253 371 5287
rect 289 5245 371 5253
rect 289 4979 371 4987
rect 289 4945 313 4979
rect 347 4945 371 4979
rect 289 4937 371 4945
rect 289 4671 371 4679
rect 289 4637 313 4671
rect 347 4637 371 4671
rect 289 4629 371 4637
rect 289 4363 371 4371
rect 289 4329 313 4363
rect 347 4329 371 4363
rect 289 4321 371 4329
rect 289 4055 371 4063
rect 289 4021 313 4055
rect 347 4021 371 4055
rect 289 4013 371 4021
rect 289 3747 371 3755
rect 289 3713 313 3747
rect 347 3713 371 3747
rect 289 3705 371 3713
rect 289 3439 371 3447
rect 289 3405 313 3439
rect 347 3405 371 3439
rect 289 3397 371 3405
rect 289 3131 371 3139
rect 289 3097 313 3131
rect 347 3097 371 3131
rect 289 3089 371 3097
rect 289 2823 371 2831
rect 289 2789 313 2823
rect 347 2789 371 2823
rect 289 2781 371 2789
rect 289 2515 371 2523
rect 289 2481 313 2515
rect 347 2481 371 2515
rect 289 2473 371 2481
rect 289 2207 371 2215
rect 289 2173 313 2207
rect 347 2173 371 2207
rect 289 2165 371 2173
rect 289 1899 371 1907
rect 289 1865 313 1899
rect 347 1865 371 1899
rect 289 1857 371 1865
rect 289 1591 371 1599
rect 289 1557 313 1591
rect 347 1557 371 1591
rect 289 1549 371 1557
rect 289 1283 371 1291
rect 289 1249 313 1283
rect 347 1249 371 1283
rect 289 1241 371 1249
rect 289 975 371 983
rect 289 941 313 975
rect 347 941 371 975
rect 289 933 371 941
rect 289 667 371 675
rect 289 633 313 667
rect 347 633 371 667
rect 289 625 371 633
rect 289 359 371 367
rect 289 325 313 359
rect 347 325 371 359
rect 289 317 371 325
rect 289 51 371 59
rect 289 17 313 51
rect 347 17 371 51
rect 289 9 371 17
<< nsubdiff >>
rect 1205 9599 1287 9607
rect 1205 9565 1229 9599
rect 1263 9565 1287 9599
rect 1205 9557 1287 9565
rect 1205 9291 1287 9299
rect 1205 9257 1229 9291
rect 1263 9257 1287 9291
rect 1205 9249 1287 9257
rect 1205 8983 1287 8991
rect 1205 8949 1229 8983
rect 1263 8949 1287 8983
rect 1205 8941 1287 8949
rect 1205 8675 1287 8683
rect 1205 8641 1229 8675
rect 1263 8641 1287 8675
rect 1205 8633 1287 8641
rect 1205 8367 1287 8375
rect 1205 8333 1229 8367
rect 1263 8333 1287 8367
rect 1205 8325 1287 8333
rect 1205 8059 1287 8067
rect 1205 8025 1229 8059
rect 1263 8025 1287 8059
rect 1205 8017 1287 8025
rect 1205 7751 1287 7759
rect 1205 7717 1229 7751
rect 1263 7717 1287 7751
rect 1205 7709 1287 7717
rect 1205 7443 1287 7451
rect 1205 7409 1229 7443
rect 1263 7409 1287 7443
rect 1205 7401 1287 7409
rect 1205 7135 1287 7143
rect 1205 7101 1229 7135
rect 1263 7101 1287 7135
rect 1205 7093 1287 7101
rect 1205 6827 1287 6835
rect 1205 6793 1229 6827
rect 1263 6793 1287 6827
rect 1205 6785 1287 6793
rect 1205 6519 1287 6527
rect 1205 6485 1229 6519
rect 1263 6485 1287 6519
rect 1205 6477 1287 6485
rect 1205 6211 1287 6219
rect 1205 6177 1229 6211
rect 1263 6177 1287 6211
rect 1205 6169 1287 6177
rect 1205 5903 1287 5911
rect 1205 5869 1229 5903
rect 1263 5869 1287 5903
rect 1205 5861 1287 5869
rect 1205 5595 1287 5603
rect 1205 5561 1229 5595
rect 1263 5561 1287 5595
rect 1205 5553 1287 5561
rect 1205 5287 1287 5295
rect 1205 5253 1229 5287
rect 1263 5253 1287 5287
rect 1205 5245 1287 5253
rect 1205 4979 1287 4987
rect 1205 4945 1229 4979
rect 1263 4945 1287 4979
rect 1205 4937 1287 4945
rect 1205 4671 1287 4679
rect 1205 4637 1229 4671
rect 1263 4637 1287 4671
rect 1205 4629 1287 4637
rect 1205 4363 1287 4371
rect 1205 4329 1229 4363
rect 1263 4329 1287 4363
rect 1205 4321 1287 4329
rect 1205 4055 1287 4063
rect 1205 4021 1229 4055
rect 1263 4021 1287 4055
rect 1205 4013 1287 4021
rect 1205 3747 1287 3755
rect 1205 3713 1229 3747
rect 1263 3713 1287 3747
rect 1205 3705 1287 3713
rect 1205 3439 1287 3447
rect 1205 3405 1229 3439
rect 1263 3405 1287 3439
rect 1205 3397 1287 3405
rect 1205 3131 1287 3139
rect 1205 3097 1229 3131
rect 1263 3097 1287 3131
rect 1205 3089 1287 3097
rect 1205 2823 1287 2831
rect 1205 2789 1229 2823
rect 1263 2789 1287 2823
rect 1205 2781 1287 2789
rect 1205 2515 1287 2523
rect 1205 2481 1229 2515
rect 1263 2481 1287 2515
rect 1205 2473 1287 2481
rect 1205 2207 1287 2215
rect 1205 2173 1229 2207
rect 1263 2173 1287 2207
rect 1205 2165 1287 2173
rect 1205 1899 1287 1907
rect 1205 1865 1229 1899
rect 1263 1865 1287 1899
rect 1205 1857 1287 1865
rect 1205 1591 1287 1599
rect 1205 1557 1229 1591
rect 1263 1557 1287 1591
rect 1205 1549 1287 1557
rect 1205 1283 1287 1291
rect 1205 1249 1229 1283
rect 1263 1249 1287 1283
rect 1205 1241 1287 1249
rect 1205 975 1287 983
rect 1205 941 1229 975
rect 1263 941 1287 975
rect 1205 933 1287 941
rect 1205 667 1287 675
rect 1205 633 1229 667
rect 1263 633 1287 667
rect 1205 625 1287 633
rect 1205 359 1287 367
rect 1205 325 1229 359
rect 1263 325 1287 359
rect 1205 317 1287 325
rect 1205 51 1287 59
rect 1205 17 1229 51
rect 1263 17 1287 51
rect 1205 9 1287 17
<< psubdiffcont >>
rect 313 9565 347 9599
rect 313 9257 347 9291
rect 313 8949 347 8983
rect 313 8641 347 8675
rect 313 8333 347 8367
rect 313 8025 347 8059
rect 313 7717 347 7751
rect 313 7409 347 7443
rect 313 7101 347 7135
rect 313 6793 347 6827
rect 313 6485 347 6519
rect 313 6177 347 6211
rect 313 5869 347 5903
rect 313 5561 347 5595
rect 313 5253 347 5287
rect 313 4945 347 4979
rect 313 4637 347 4671
rect 313 4329 347 4363
rect 313 4021 347 4055
rect 313 3713 347 3747
rect 313 3405 347 3439
rect 313 3097 347 3131
rect 313 2789 347 2823
rect 313 2481 347 2515
rect 313 2173 347 2207
rect 313 1865 347 1899
rect 313 1557 347 1591
rect 313 1249 347 1283
rect 313 941 347 975
rect 313 633 347 667
rect 313 325 347 359
rect 313 17 347 51
<< nsubdiffcont >>
rect 1229 9565 1263 9599
rect 1229 9257 1263 9291
rect 1229 8949 1263 8983
rect 1229 8641 1263 8675
rect 1229 8333 1263 8367
rect 1229 8025 1263 8059
rect 1229 7717 1263 7751
rect 1229 7409 1263 7443
rect 1229 7101 1263 7135
rect 1229 6793 1263 6827
rect 1229 6485 1263 6519
rect 1229 6177 1263 6211
rect 1229 5869 1263 5903
rect 1229 5561 1263 5595
rect 1229 5253 1263 5287
rect 1229 4945 1263 4979
rect 1229 4637 1263 4671
rect 1229 4329 1263 4363
rect 1229 4021 1263 4055
rect 1229 3713 1263 3747
rect 1229 3405 1263 3439
rect 1229 3097 1263 3131
rect 1229 2789 1263 2823
rect 1229 2481 1263 2515
rect 1229 2173 1263 2207
rect 1229 1865 1263 1899
rect 1229 1557 1263 1591
rect 1229 1249 1263 1283
rect 1229 941 1263 975
rect 1229 633 1263 667
rect 1229 325 1263 359
rect 1229 17 1263 51
<< locali >>
rect 60 9703 94 9769
rect 1748 9686 1782 9753
rect 297 9565 313 9599
rect 347 9565 363 9599
rect 1213 9565 1229 9599
rect 1263 9565 1279 9599
rect 60 9395 94 9461
rect 1748 9378 1782 9445
rect 297 9257 313 9291
rect 347 9257 363 9291
rect 1213 9257 1229 9291
rect 1263 9257 1279 9291
rect 60 9087 94 9153
rect 1748 9070 1782 9137
rect 297 8949 313 8983
rect 347 8949 363 8983
rect 1213 8949 1229 8983
rect 1263 8949 1279 8983
rect 60 8779 94 8845
rect 1748 8762 1782 8829
rect 297 8641 313 8675
rect 347 8641 363 8675
rect 1213 8641 1229 8675
rect 1263 8641 1279 8675
rect 60 8471 94 8537
rect 1748 8454 1782 8521
rect 297 8333 313 8367
rect 347 8333 363 8367
rect 1213 8333 1229 8367
rect 1263 8333 1279 8367
rect 60 8163 94 8229
rect 1748 8146 1782 8213
rect 297 8025 313 8059
rect 347 8025 363 8059
rect 1213 8025 1229 8059
rect 1263 8025 1279 8059
rect 60 7855 94 7921
rect 1748 7838 1782 7905
rect 297 7717 313 7751
rect 347 7717 363 7751
rect 1213 7717 1229 7751
rect 1263 7717 1279 7751
rect 60 7547 94 7613
rect 1748 7530 1782 7597
rect 297 7409 313 7443
rect 347 7409 363 7443
rect 1213 7409 1229 7443
rect 1263 7409 1279 7443
rect 60 7239 94 7305
rect 1748 7222 1782 7289
rect 297 7101 313 7135
rect 347 7101 363 7135
rect 1213 7101 1229 7135
rect 1263 7101 1279 7135
rect 60 6931 94 6997
rect 1748 6914 1782 6981
rect 297 6793 313 6827
rect 347 6793 363 6827
rect 1213 6793 1229 6827
rect 1263 6793 1279 6827
rect 60 6623 94 6689
rect 1748 6606 1782 6673
rect 297 6485 313 6519
rect 347 6485 363 6519
rect 1213 6485 1229 6519
rect 1263 6485 1279 6519
rect 60 6315 94 6381
rect 1748 6298 1782 6365
rect 297 6177 313 6211
rect 347 6177 363 6211
rect 1213 6177 1229 6211
rect 1263 6177 1279 6211
rect 60 6007 94 6073
rect 1748 5990 1782 6057
rect 297 5869 313 5903
rect 347 5869 363 5903
rect 1213 5869 1229 5903
rect 1263 5869 1279 5903
rect 60 5699 94 5765
rect 1748 5682 1782 5749
rect 297 5561 313 5595
rect 347 5561 363 5595
rect 1213 5561 1229 5595
rect 1263 5561 1279 5595
rect 60 5391 94 5457
rect 1748 5374 1782 5441
rect 297 5253 313 5287
rect 347 5253 363 5287
rect 1213 5253 1229 5287
rect 1263 5253 1279 5287
rect 60 5083 94 5149
rect 1748 5066 1782 5133
rect 297 4945 313 4979
rect 347 4945 363 4979
rect 1213 4945 1229 4979
rect 1263 4945 1279 4979
rect 60 4775 94 4841
rect 1748 4758 1782 4825
rect 297 4637 313 4671
rect 347 4637 363 4671
rect 1213 4637 1229 4671
rect 1263 4637 1279 4671
rect 60 4467 94 4533
rect 1748 4450 1782 4517
rect 297 4329 313 4363
rect 347 4329 363 4363
rect 1213 4329 1229 4363
rect 1263 4329 1279 4363
rect 60 4159 94 4225
rect 1748 4142 1782 4209
rect 297 4021 313 4055
rect 347 4021 363 4055
rect 1213 4021 1229 4055
rect 1263 4021 1279 4055
rect 60 3851 94 3917
rect 1748 3834 1782 3901
rect 297 3713 313 3747
rect 347 3713 363 3747
rect 1213 3713 1229 3747
rect 1263 3713 1279 3747
rect 60 3543 94 3609
rect 1748 3526 1782 3593
rect 297 3405 313 3439
rect 347 3405 363 3439
rect 1213 3405 1229 3439
rect 1263 3405 1279 3439
rect 60 3235 94 3301
rect 1748 3218 1782 3285
rect 297 3097 313 3131
rect 347 3097 363 3131
rect 1213 3097 1229 3131
rect 1263 3097 1279 3131
rect 60 2927 94 2993
rect 1748 2910 1782 2977
rect 297 2789 313 2823
rect 347 2789 363 2823
rect 1213 2789 1229 2823
rect 1263 2789 1279 2823
rect 60 2619 94 2685
rect 1748 2602 1782 2669
rect 297 2481 313 2515
rect 347 2481 363 2515
rect 1213 2481 1229 2515
rect 1263 2481 1279 2515
rect 60 2311 94 2377
rect 1748 2294 1782 2361
rect 297 2173 313 2207
rect 347 2173 363 2207
rect 1213 2173 1229 2207
rect 1263 2173 1279 2207
rect 60 2003 94 2069
rect 1748 1986 1782 2053
rect 297 1865 313 1899
rect 347 1865 363 1899
rect 1213 1865 1229 1899
rect 1263 1865 1279 1899
rect 60 1695 94 1761
rect 1748 1678 1782 1745
rect 297 1557 313 1591
rect 347 1557 363 1591
rect 1213 1557 1229 1591
rect 1263 1557 1279 1591
rect 60 1387 94 1453
rect 1748 1370 1782 1437
rect 297 1249 313 1283
rect 347 1249 363 1283
rect 1213 1249 1229 1283
rect 1263 1249 1279 1283
rect 60 1079 94 1145
rect 1748 1062 1782 1129
rect 297 941 313 975
rect 347 941 363 975
rect 1213 941 1229 975
rect 1263 941 1279 975
rect 60 771 94 837
rect 1748 754 1782 821
rect 297 633 313 667
rect 347 633 363 667
rect 1213 633 1229 667
rect 1263 633 1279 667
rect 60 463 94 529
rect 1748 446 1782 513
rect 297 325 313 359
rect 347 325 363 359
rect 1213 325 1229 359
rect 1263 325 1279 359
rect 60 155 94 221
rect 1748 138 1782 205
rect 297 17 313 51
rect 347 17 363 51
rect 1213 17 1229 51
rect 1263 17 1279 51
<< viali >>
rect 313 9565 347 9599
rect 1229 9565 1263 9599
rect 313 9257 347 9291
rect 1229 9257 1263 9291
rect 313 8949 347 8983
rect 1229 8949 1263 8983
rect 313 8641 347 8675
rect 1229 8641 1263 8675
rect 313 8333 347 8367
rect 1229 8333 1263 8367
rect 313 8025 347 8059
rect 1229 8025 1263 8059
rect 313 7717 347 7751
rect 1229 7717 1263 7751
rect 313 7409 347 7443
rect 1229 7409 1263 7443
rect 313 7101 347 7135
rect 1229 7101 1263 7135
rect 313 6793 347 6827
rect 1229 6793 1263 6827
rect 313 6485 347 6519
rect 1229 6485 1263 6519
rect 313 6177 347 6211
rect 1229 6177 1263 6211
rect 313 5869 347 5903
rect 1229 5869 1263 5903
rect 313 5561 347 5595
rect 1229 5561 1263 5595
rect 313 5253 347 5287
rect 1229 5253 1263 5287
rect 313 4945 347 4979
rect 1229 4945 1263 4979
rect 313 4637 347 4671
rect 1229 4637 1263 4671
rect 313 4329 347 4363
rect 1229 4329 1263 4363
rect 313 4021 347 4055
rect 1229 4021 1263 4055
rect 313 3713 347 3747
rect 1229 3713 1263 3747
rect 313 3405 347 3439
rect 1229 3405 1263 3439
rect 313 3097 347 3131
rect 1229 3097 1263 3131
rect 313 2789 347 2823
rect 1229 2789 1263 2823
rect 313 2481 347 2515
rect 1229 2481 1263 2515
rect 313 2173 347 2207
rect 1229 2173 1263 2207
rect 313 1865 347 1899
rect 1229 1865 1263 1899
rect 313 1557 347 1591
rect 1229 1557 1263 1591
rect 313 1249 347 1283
rect 1229 1249 1263 1283
rect 313 941 347 975
rect 1229 941 1263 975
rect 313 633 347 667
rect 1229 633 1263 667
rect 313 325 347 359
rect 1229 325 1263 359
rect 313 17 347 51
rect 1229 17 1263 51
<< metal1 >>
rect 316 9611 344 9870
rect 1232 9611 1260 9870
rect 307 9599 353 9611
rect 307 9565 313 9599
rect 347 9565 353 9599
rect 307 9553 353 9565
rect 1223 9599 1269 9611
rect 1223 9565 1229 9599
rect 1263 9565 1269 9599
rect 1223 9553 1269 9565
rect 316 9303 344 9553
rect 1232 9303 1260 9553
rect 307 9291 353 9303
rect 307 9257 313 9291
rect 347 9257 353 9291
rect 307 9245 353 9257
rect 1223 9291 1269 9303
rect 1223 9257 1229 9291
rect 1263 9257 1269 9291
rect 1223 9245 1269 9257
rect 316 8995 344 9245
rect 1232 8995 1260 9245
rect 307 8983 353 8995
rect 307 8949 313 8983
rect 347 8949 353 8983
rect 307 8937 353 8949
rect 1223 8983 1269 8995
rect 1223 8949 1229 8983
rect 1263 8949 1269 8983
rect 1223 8937 1269 8949
rect 316 8687 344 8937
rect 1232 8687 1260 8937
rect 307 8675 353 8687
rect 307 8641 313 8675
rect 347 8641 353 8675
rect 307 8629 353 8641
rect 1223 8675 1269 8687
rect 1223 8641 1229 8675
rect 1263 8641 1269 8675
rect 1223 8629 1269 8641
rect 316 8379 344 8629
rect 1232 8379 1260 8629
rect 307 8367 353 8379
rect 307 8333 313 8367
rect 347 8333 353 8367
rect 307 8321 353 8333
rect 1223 8367 1269 8379
rect 1223 8333 1229 8367
rect 1263 8333 1269 8367
rect 1223 8321 1269 8333
rect 316 8071 344 8321
rect 1232 8071 1260 8321
rect 307 8059 353 8071
rect 307 8025 313 8059
rect 347 8025 353 8059
rect 307 8013 353 8025
rect 1223 8059 1269 8071
rect 1223 8025 1229 8059
rect 1263 8025 1269 8059
rect 1223 8013 1269 8025
rect 316 7763 344 8013
rect 1232 7763 1260 8013
rect 307 7751 353 7763
rect 307 7717 313 7751
rect 347 7717 353 7751
rect 307 7705 353 7717
rect 1223 7751 1269 7763
rect 1223 7717 1229 7751
rect 1263 7717 1269 7751
rect 1223 7705 1269 7717
rect 316 7455 344 7705
rect 1232 7455 1260 7705
rect 307 7443 353 7455
rect 307 7409 313 7443
rect 347 7409 353 7443
rect 307 7397 353 7409
rect 1223 7443 1269 7455
rect 1223 7409 1229 7443
rect 1263 7409 1269 7443
rect 1223 7397 1269 7409
rect 316 7147 344 7397
rect 1232 7147 1260 7397
rect 307 7135 353 7147
rect 307 7101 313 7135
rect 347 7101 353 7135
rect 307 7089 353 7101
rect 1223 7135 1269 7147
rect 1223 7101 1229 7135
rect 1263 7101 1269 7135
rect 1223 7089 1269 7101
rect 316 6839 344 7089
rect 1232 6839 1260 7089
rect 307 6827 353 6839
rect 307 6793 313 6827
rect 347 6793 353 6827
rect 307 6781 353 6793
rect 1223 6827 1269 6839
rect 1223 6793 1229 6827
rect 1263 6793 1269 6827
rect 1223 6781 1269 6793
rect 316 6531 344 6781
rect 1232 6531 1260 6781
rect 307 6519 353 6531
rect 307 6485 313 6519
rect 347 6485 353 6519
rect 307 6473 353 6485
rect 1223 6519 1269 6531
rect 1223 6485 1229 6519
rect 1263 6485 1269 6519
rect 1223 6473 1269 6485
rect 316 6223 344 6473
rect 1232 6223 1260 6473
rect 307 6211 353 6223
rect 307 6177 313 6211
rect 347 6177 353 6211
rect 307 6165 353 6177
rect 1223 6211 1269 6223
rect 1223 6177 1229 6211
rect 1263 6177 1269 6211
rect 1223 6165 1269 6177
rect 316 5915 344 6165
rect 1232 5915 1260 6165
rect 307 5903 353 5915
rect 307 5869 313 5903
rect 347 5869 353 5903
rect 307 5857 353 5869
rect 1223 5903 1269 5915
rect 1223 5869 1229 5903
rect 1263 5869 1269 5903
rect 1223 5857 1269 5869
rect 316 5607 344 5857
rect 1232 5607 1260 5857
rect 307 5595 353 5607
rect 307 5561 313 5595
rect 347 5561 353 5595
rect 307 5549 353 5561
rect 1223 5595 1269 5607
rect 1223 5561 1229 5595
rect 1263 5561 1269 5595
rect 1223 5549 1269 5561
rect 316 5299 344 5549
rect 1232 5299 1260 5549
rect 307 5287 353 5299
rect 307 5253 313 5287
rect 347 5253 353 5287
rect 307 5241 353 5253
rect 1223 5287 1269 5299
rect 1223 5253 1229 5287
rect 1263 5253 1269 5287
rect 1223 5241 1269 5253
rect 316 4991 344 5241
rect 1232 4991 1260 5241
rect 307 4979 353 4991
rect 307 4945 313 4979
rect 347 4945 353 4979
rect 307 4933 353 4945
rect 1223 4979 1269 4991
rect 1223 4945 1229 4979
rect 1263 4945 1269 4979
rect 1223 4933 1269 4945
rect 316 4683 344 4933
rect 1232 4683 1260 4933
rect 307 4671 353 4683
rect 307 4637 313 4671
rect 347 4637 353 4671
rect 307 4625 353 4637
rect 1223 4671 1269 4683
rect 1223 4637 1229 4671
rect 1263 4637 1269 4671
rect 1223 4625 1269 4637
rect 316 4375 344 4625
rect 1232 4375 1260 4625
rect 307 4363 353 4375
rect 307 4329 313 4363
rect 347 4329 353 4363
rect 307 4317 353 4329
rect 1223 4363 1269 4375
rect 1223 4329 1229 4363
rect 1263 4329 1269 4363
rect 1223 4317 1269 4329
rect 316 4067 344 4317
rect 1232 4067 1260 4317
rect 307 4055 353 4067
rect 307 4021 313 4055
rect 347 4021 353 4055
rect 307 4009 353 4021
rect 1223 4055 1269 4067
rect 1223 4021 1229 4055
rect 1263 4021 1269 4055
rect 1223 4009 1269 4021
rect 316 3759 344 4009
rect 1232 3759 1260 4009
rect 307 3747 353 3759
rect 307 3713 313 3747
rect 347 3713 353 3747
rect 307 3701 353 3713
rect 1223 3747 1269 3759
rect 1223 3713 1229 3747
rect 1263 3713 1269 3747
rect 1223 3701 1269 3713
rect 316 3451 344 3701
rect 1232 3451 1260 3701
rect 307 3439 353 3451
rect 307 3405 313 3439
rect 347 3405 353 3439
rect 307 3393 353 3405
rect 1223 3439 1269 3451
rect 1223 3405 1229 3439
rect 1263 3405 1269 3439
rect 1223 3393 1269 3405
rect 316 3143 344 3393
rect 1232 3143 1260 3393
rect 307 3131 353 3143
rect 307 3097 313 3131
rect 347 3097 353 3131
rect 307 3085 353 3097
rect 1223 3131 1269 3143
rect 1223 3097 1229 3131
rect 1263 3097 1269 3131
rect 1223 3085 1269 3097
rect 316 2835 344 3085
rect 1232 2835 1260 3085
rect 307 2823 353 2835
rect 307 2789 313 2823
rect 347 2789 353 2823
rect 307 2777 353 2789
rect 1223 2823 1269 2835
rect 1223 2789 1229 2823
rect 1263 2789 1269 2823
rect 1223 2777 1269 2789
rect 316 2527 344 2777
rect 1232 2527 1260 2777
rect 307 2515 353 2527
rect 307 2481 313 2515
rect 347 2481 353 2515
rect 307 2469 353 2481
rect 1223 2515 1269 2527
rect 1223 2481 1229 2515
rect 1263 2481 1269 2515
rect 1223 2469 1269 2481
rect 316 2219 344 2469
rect 1232 2219 1260 2469
rect 307 2207 353 2219
rect 307 2173 313 2207
rect 347 2173 353 2207
rect 307 2161 353 2173
rect 1223 2207 1269 2219
rect 1223 2173 1229 2207
rect 1263 2173 1269 2207
rect 1223 2161 1269 2173
rect 316 1911 344 2161
rect 1232 1911 1260 2161
rect 307 1899 353 1911
rect 307 1865 313 1899
rect 347 1865 353 1899
rect 307 1853 353 1865
rect 1223 1899 1269 1911
rect 1223 1865 1229 1899
rect 1263 1865 1269 1899
rect 1223 1853 1269 1865
rect 316 1603 344 1853
rect 1232 1603 1260 1853
rect 307 1591 353 1603
rect 307 1557 313 1591
rect 347 1557 353 1591
rect 307 1545 353 1557
rect 1223 1591 1269 1603
rect 1223 1557 1229 1591
rect 1263 1557 1269 1591
rect 1223 1545 1269 1557
rect 316 1295 344 1545
rect 1232 1295 1260 1545
rect 307 1283 353 1295
rect 307 1249 313 1283
rect 347 1249 353 1283
rect 307 1237 353 1249
rect 1223 1283 1269 1295
rect 1223 1249 1229 1283
rect 1263 1249 1269 1283
rect 1223 1237 1269 1249
rect 316 987 344 1237
rect 1232 987 1260 1237
rect 307 975 353 987
rect 307 941 313 975
rect 347 941 353 975
rect 307 929 353 941
rect 1223 975 1269 987
rect 1223 941 1229 975
rect 1263 941 1269 975
rect 1223 929 1269 941
rect 316 679 344 929
rect 1232 679 1260 929
rect 307 667 353 679
rect 307 633 313 667
rect 347 633 353 667
rect 307 621 353 633
rect 1223 667 1269 679
rect 1223 633 1229 667
rect 1263 633 1269 667
rect 1223 621 1269 633
rect 316 371 344 621
rect 1232 371 1260 621
rect 307 359 353 371
rect 307 325 313 359
rect 347 325 353 359
rect 307 313 353 325
rect 1223 359 1269 371
rect 1223 325 1229 359
rect 1263 325 1269 359
rect 1223 313 1269 325
rect 316 63 344 313
rect 1232 63 1260 313
rect 307 51 353 63
rect 307 17 313 51
rect 347 17 353 51
rect 307 5 353 17
rect 1223 51 1269 63
rect 1223 17 1229 51
rect 1263 17 1269 51
rect 1223 5 1269 17
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_0
timestamp 1581449089
transform 1 0 0 0 1 9652
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_1
timestamp 1581449089
transform 1 0 0 0 1 9344
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_2
timestamp 1581449089
transform 1 0 0 0 1 9036
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_3
timestamp 1581449089
transform 1 0 0 0 1 8728
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_4
timestamp 1581449089
transform 1 0 0 0 1 8420
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_5
timestamp 1581449089
transform 1 0 0 0 1 8112
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_6
timestamp 1581449089
transform 1 0 0 0 1 7804
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_7
timestamp 1581449089
transform 1 0 0 0 1 7496
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_8
timestamp 1581449089
transform 1 0 0 0 1 7188
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_9
timestamp 1581449089
transform 1 0 0 0 1 6880
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_10
timestamp 1581449089
transform 1 0 0 0 1 6572
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_11
timestamp 1581449089
transform 1 0 0 0 1 6264
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_12
timestamp 1581449089
transform 1 0 0 0 1 5956
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_13
timestamp 1581449089
transform 1 0 0 0 1 5648
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_14
timestamp 1581449089
transform 1 0 0 0 1 5340
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_15
timestamp 1581449089
transform 1 0 0 0 1 5032
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_16
timestamp 1581449089
transform 1 0 0 0 1 4724
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_17
timestamp 1581449089
transform 1 0 0 0 1 4416
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_18
timestamp 1581449089
transform 1 0 0 0 1 4108
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_19
timestamp 1581449089
transform 1 0 0 0 1 3800
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_20
timestamp 1581449089
transform 1 0 0 0 1 3492
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_21
timestamp 1581449089
transform 1 0 0 0 1 3184
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_22
timestamp 1581449089
transform 1 0 0 0 1 2876
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_23
timestamp 1581449089
transform 1 0 0 0 1 2568
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_24
timestamp 1581449089
transform 1 0 0 0 1 2260
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_25
timestamp 1581449089
transform 1 0 0 0 1 1952
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_26
timestamp 1581449089
transform 1 0 0 0 1 1644
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_27
timestamp 1581449089
transform 1 0 0 0 1 1336
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_28
timestamp 1581449089
transform 1 0 0 0 1 1028
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_29
timestamp 1581449089
transform 1 0 0 0 1 720
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_30
timestamp 1581449089
transform 1 0 0 0 1 412
box 44 -50 1800 299
use sky130_rom_krom_pinv_dec_4  sky130_rom_krom_pinv_dec_4_31
timestamp 1581449089
transform 1 0 0 0 1 104
box 44 -50 1800 299
<< labels >>
rlabel locali s 77 188 77 188 4 in_0
port 2 nsew
rlabel locali s 1765 188 1765 188 4 out_0
port 3 nsew
rlabel locali s 77 496 77 496 4 in_1
port 4 nsew
rlabel locali s 1765 496 1765 496 4 out_1
port 5 nsew
rlabel locali s 77 804 77 804 4 in_2
port 6 nsew
rlabel locali s 1765 804 1765 804 4 out_2
port 7 nsew
rlabel locali s 77 1112 77 1112 4 in_3
port 8 nsew
rlabel locali s 1765 1112 1765 1112 4 out_3
port 9 nsew
rlabel locali s 77 1420 77 1420 4 in_4
port 10 nsew
rlabel locali s 1765 1420 1765 1420 4 out_4
port 11 nsew
rlabel locali s 77 1728 77 1728 4 in_5
port 12 nsew
rlabel locali s 1765 1728 1765 1728 4 out_5
port 13 nsew
rlabel locali s 77 2036 77 2036 4 in_6
port 14 nsew
rlabel locali s 1765 2036 1765 2036 4 out_6
port 15 nsew
rlabel locali s 77 2344 77 2344 4 in_7
port 16 nsew
rlabel locali s 1765 2344 1765 2344 4 out_7
port 17 nsew
rlabel locali s 77 2652 77 2652 4 in_8
port 18 nsew
rlabel locali s 1765 2652 1765 2652 4 out_8
port 19 nsew
rlabel locali s 77 2960 77 2960 4 in_9
port 20 nsew
rlabel locali s 1765 2960 1765 2960 4 out_9
port 21 nsew
rlabel locali s 77 3268 77 3268 4 in_10
port 22 nsew
rlabel locali s 1765 3268 1765 3268 4 out_10
port 23 nsew
rlabel locali s 77 3576 77 3576 4 in_11
port 24 nsew
rlabel locali s 1765 3576 1765 3576 4 out_11
port 25 nsew
rlabel locali s 77 3884 77 3884 4 in_12
port 26 nsew
rlabel locali s 1765 3884 1765 3884 4 out_12
port 27 nsew
rlabel locali s 77 4192 77 4192 4 in_13
port 28 nsew
rlabel locali s 1765 4192 1765 4192 4 out_13
port 29 nsew
rlabel locali s 77 4500 77 4500 4 in_14
port 30 nsew
rlabel locali s 1765 4500 1765 4500 4 out_14
port 31 nsew
rlabel locali s 77 4808 77 4808 4 in_15
port 32 nsew
rlabel locali s 1765 4808 1765 4808 4 out_15
port 33 nsew
rlabel locali s 77 5116 77 5116 4 in_16
port 34 nsew
rlabel locali s 1765 5116 1765 5116 4 out_16
port 35 nsew
rlabel locali s 77 5424 77 5424 4 in_17
port 36 nsew
rlabel locali s 1765 5424 1765 5424 4 out_17
port 37 nsew
rlabel locali s 77 5732 77 5732 4 in_18
port 38 nsew
rlabel locali s 1765 5732 1765 5732 4 out_18
port 39 nsew
rlabel locali s 77 6040 77 6040 4 in_19
port 40 nsew
rlabel locali s 1765 6040 1765 6040 4 out_19
port 41 nsew
rlabel locali s 77 6348 77 6348 4 in_20
port 42 nsew
rlabel locali s 1765 6348 1765 6348 4 out_20
port 43 nsew
rlabel locali s 77 6656 77 6656 4 in_21
port 44 nsew
rlabel locali s 1765 6656 1765 6656 4 out_21
port 45 nsew
rlabel locali s 77 6964 77 6964 4 in_22
port 46 nsew
rlabel locali s 1765 6964 1765 6964 4 out_22
port 47 nsew
rlabel locali s 77 7272 77 7272 4 in_23
port 48 nsew
rlabel locali s 1765 7272 1765 7272 4 out_23
port 49 nsew
rlabel locali s 77 7580 77 7580 4 in_24
port 50 nsew
rlabel locali s 1765 7580 1765 7580 4 out_24
port 51 nsew
rlabel locali s 77 7888 77 7888 4 in_25
port 52 nsew
rlabel locali s 1765 7888 1765 7888 4 out_25
port 53 nsew
rlabel locali s 77 8196 77 8196 4 in_26
port 54 nsew
rlabel locali s 1765 8196 1765 8196 4 out_26
port 55 nsew
rlabel locali s 77 8504 77 8504 4 in_27
port 56 nsew
rlabel locali s 1765 8504 1765 8504 4 out_27
port 57 nsew
rlabel locali s 77 8812 77 8812 4 in_28
port 58 nsew
rlabel locali s 1765 8812 1765 8812 4 out_28
port 59 nsew
rlabel locali s 77 9120 77 9120 4 in_29
port 60 nsew
rlabel locali s 1765 9120 1765 9120 4 out_29
port 61 nsew
rlabel locali s 77 9428 77 9428 4 in_30
port 62 nsew
rlabel locali s 1765 9428 1765 9428 4 out_30
port 63 nsew
rlabel locali s 77 9736 77 9736 4 in_31
port 64 nsew
rlabel locali s 1765 9736 1765 9736 4 out_31
port 65 nsew
rlabel metal1 s 316 9842 344 9870 4 gnd
port 67 nsew
rlabel metal1 s 316 6 344 34 4 gnd
port 67 nsew
rlabel metal1 s 1232 6 1260 34 4 vdd
port 69 nsew
rlabel metal1 s 1232 9842 1260 9870 4 vdd
port 69 nsew
<< properties >>
string FIXED_BBOX 1162 -50 1330 0
<< end >>
