* NGSPICE file created from sky130_rom_krom.ext - technology: sky130A

.subckt sky130_rom_krom_rom_base_one_cell G D S gnd
X0 D G S gnd sky130_fd_pr__nfet_01v8 ad=0.108p pd=1.32u as=0.108p ps=1.32u w=0.36u l=0.15u
.ends

.subckt sky130_rom_krom_rom_base_zero_cell G S gnd
X0 S G S gnd sky130_fd_pr__nfet_01v8 ad=0.216p pd=2.64u as=0p ps=0u w=0.36u l=0.15u
.ends

.subckt sky130_rom_krom_precharge_cell D G vdd
X0 D G vdd vdd sky130_fd_pr__pfet_01v8 ad=0.126p pd=1.44u as=0.126p ps=1.44u w=0.42u l=0.15u
.ends

.subckt sky130_rom_krom_rom_precharge_array_0 pre_bl0_out pre_bl2_out pre_bl3_out
+ pre_bl6_out pre_bl4_out vdd pre_bl7_out gate pre_bl5_out pre_bl1_out
Xsky130_rom_krom_precharge_cell_2 pre_bl5_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_3 pre_bl4_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_4 pre_bl3_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_5 pre_bl2_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_6 pre_bl1_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_7 pre_bl0_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_0 pre_bl7_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_1 pre_bl6_out gate vdd sky130_rom_krom_precharge_cell
.ends

.subckt sky130_rom_krom_rom_row_decode_array bl_0_0 bl_0_1 bl_0_2 bl_0_3 bl_0_4 bl_0_5
+ bl_0_6 bl_0_7 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 gnd wl_0_0 vdd precharge
Xsky130_rom_krom_rom_base_one_cell_30 wl_0_0 sky130_rom_krom_rom_base_one_cell_30/D
+ bl_0_1 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_20 wl_0_2 sky130_rom_krom_rom_base_one_cell_9/S
+ sky130_rom_krom_rom_base_one_cell_26/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_31 wl_0_0 sky130_rom_krom_rom_base_one_cell_31/D
+ bl_0_0 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_10 wl_0_5 sky130_rom_krom_rom_base_one_cell_4/S
+ sky130_rom_krom_rom_base_zero_cell_6/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_21 wl_0_2 sky130_rom_krom_rom_base_zero_cell_9/S
+ sky130_rom_krom_rom_base_one_cell_27/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_11 wl_0_5 sky130_rom_krom_rom_base_one_cell_6/S
+ sky130_rom_krom_rom_base_zero_cell_7/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_22 wl_0_2 sky130_rom_krom_rom_base_zero_cell_7/S
+ sky130_rom_krom_rom_base_one_cell_30/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_0 precharge gnd sky130_rom_krom_rom_base_one_cell_8/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_12 wl_0_4 sky130_rom_krom_rom_base_one_cell_1/S
+ sky130_rom_krom_rom_base_one_cell_17/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_23 wl_0_2 sky130_rom_krom_rom_base_one_cell_23/D
+ sky130_rom_krom_rom_base_one_cell_31/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1 precharge gnd sky130_rom_krom_rom_base_one_cell_1/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_13 wl_0_4 sky130_rom_krom_rom_base_one_cell_3/S
+ sky130_rom_krom_rom_base_zero_cell_9/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_24 wl_0_1 sky130_rom_krom_rom_base_one_cell_24/D
+ bl_0_7 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_2 precharge gnd sky130_rom_krom_rom_base_one_cell_9/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_0 wl_0_5 sky130_rom_krom_rom_base_one_cell_1/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_14 wl_0_4 sky130_rom_krom_rom_base_one_cell_5/S
+ sky130_rom_krom_rom_base_one_cell_19/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_25 wl_0_1 sky130_rom_krom_rom_base_one_cell_25/D
+ bl_0_6 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_3 precharge gnd sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1 wl_0_5 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_2 wl_0_5 sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_15 wl_0_4 sky130_rom_krom_rom_base_one_cell_7/S
+ sky130_rom_krom_rom_base_one_cell_23/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_26 wl_0_1 sky130_rom_krom_rom_base_one_cell_26/D
+ bl_0_5 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_precharge_array_0_0 bl_0_0 bl_0_2 bl_0_3 bl_0_6 bl_0_4 vdd bl_0_7
+ precharge bl_0_5 bl_0_1 sky130_rom_krom_rom_precharge_array_0
Xsky130_rom_krom_rom_base_one_cell_4 precharge gnd sky130_rom_krom_rom_base_one_cell_4/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_3 wl_0_5 sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_16 wl_0_3 sky130_rom_krom_rom_base_one_cell_8/S
+ sky130_rom_krom_rom_base_one_cell_24/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_17 wl_0_3 sky130_rom_krom_rom_base_one_cell_17/D
+ sky130_rom_krom_rom_base_one_cell_25/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_28 wl_0_0 sky130_rom_krom_rom_base_one_cell_28/D
+ bl_0_3 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_27 wl_0_1 sky130_rom_krom_rom_base_one_cell_27/D
+ bl_0_4 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_5 precharge gnd sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_4 wl_0_4 sky130_rom_krom_rom_base_one_cell_8/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_18 wl_0_3 sky130_rom_krom_rom_base_zero_cell_6/S
+ sky130_rom_krom_rom_base_one_cell_28/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_29 wl_0_0 sky130_rom_krom_rom_base_one_cell_29/D
+ bl_0_2 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_7 precharge gnd sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_6 precharge gnd sky130_rom_krom_rom_base_one_cell_6/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_5 wl_0_4 sky130_rom_krom_rom_base_one_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_19 wl_0_3 sky130_rom_krom_rom_base_one_cell_19/D
+ sky130_rom_krom_rom_base_one_cell_29/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_8 wl_0_5 sky130_rom_krom_rom_base_one_cell_8/D
+ sky130_rom_krom_rom_base_one_cell_8/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_6 wl_0_4 sky130_rom_krom_rom_base_zero_cell_6/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_9 wl_0_5 sky130_rom_krom_rom_base_one_cell_9/D
+ sky130_rom_krom_rom_base_one_cell_9/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_7 wl_0_4 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_20 wl_0_0 bl_0_7 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_8 wl_0_3 sky130_rom_krom_rom_base_one_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_10 wl_0_3 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_21 wl_0_0 bl_0_6 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_9 wl_0_3 sky130_rom_krom_rom_base_zero_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_11 wl_0_3 sky130_rom_krom_rom_base_one_cell_23/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_22 wl_0_0 bl_0_5 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_12 wl_0_2 sky130_rom_krom_rom_base_one_cell_24/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_23 wl_0_0 bl_0_4 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_13 wl_0_2 sky130_rom_krom_rom_base_one_cell_25/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_14 wl_0_2 sky130_rom_krom_rom_base_one_cell_28/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_15 wl_0_2 sky130_rom_krom_rom_base_one_cell_29/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_16 wl_0_1 sky130_rom_krom_rom_base_one_cell_28/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_17 wl_0_1 sky130_rom_krom_rom_base_one_cell_29/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_18 wl_0_1 sky130_rom_krom_rom_base_one_cell_30/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_19 wl_0_1 sky130_rom_krom_rom_base_one_cell_31/D
+ gnd sky130_rom_krom_rom_base_zero_cell
.ends

.subckt sky130_rom_krom_inv_array_mod A Z vdd gnd w_504_0#
X0 vdd A Z w_504_0# sky130_fd_pr__pfet_01v8 ad=0.9p pd=6.6u as=0.9p ps=6.6u w=3u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.222p pd=2.08u as=0.222p ps=2.08u w=0.74u l=0.15u
.ends

.subckt sky130_fd_bd_sram__openram_sp_nand2_dec A B Z vdd gnd
X0 vdd B Z vdd sky130_fd_pr__pfet_01v8 ad=0.336p pd=2.84u as=0.6776p ps=5.69u w=1.12u l=0.15u
X1 a_174_144# B gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1554p pd=1.9u as=0.222p ps=2.08u w=0.74u l=0.15u
X2 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12u l=0.15u
X3 Z A a_174_144# gnd sky130_fd_pr__nfet_01v8 ad=0.2701p pd=2.21u as=0p ps=0u w=0.74u l=0.15u
.ends

.subckt sky130_rom_krom_rom_address_control_buf A_in A_out Abar_out clk vdd_uq0 vdd_uq1
+ vdd gnd
Xsky130_rom_krom_inv_array_mod_0 A_in sky130_rom_krom_inv_array_mod_0/Z vdd_uq1 gnd
+ vdd_uq1 sky130_rom_krom_inv_array_mod
Xsky130_fd_bd_sram__openram_sp_nand2_dec_0 clk A_out Abar_out vdd gnd sky130_fd_bd_sram__openram_sp_nand2_dec
Xsky130_fd_bd_sram__openram_sp_nand2_dec_1 clk sky130_rom_krom_inv_array_mod_0/Z A_out
+ vdd_uq0 gnd sky130_fd_bd_sram__openram_sp_nand2_dec
.ends

.subckt sky130_rom_krom_rom_address_control_array A0_in A1_in A2_in A0_out A1_out
+ A2_out Abar0_out Abar1_out clk vdd gnd vdd_uq0 vdd_uq1 Abar2_out
Xsky130_rom_krom_rom_address_control_buf_0 A2_in A2_out Abar2_out clk vdd vdd_uq0
+ vdd_uq1 gnd sky130_rom_krom_rom_address_control_buf
Xsky130_rom_krom_rom_address_control_buf_2 A0_in A0_out Abar0_out clk vdd vdd_uq0
+ vdd_uq1 gnd sky130_rom_krom_rom_address_control_buf
Xsky130_rom_krom_rom_address_control_buf_1 A1_in A1_out Abar1_out clk vdd vdd_uq0
+ vdd_uq1 gnd sky130_rom_krom_rom_address_control_buf
.ends

.subckt sky130_rom_krom_pinv_dec_1 A Z vdd w_1756_n45# gnd
X0 vdd A Z w_1756_n45# sky130_fd_pr__pfet_01v8 ad=2.1p pd=14.6u as=2.1p ps=14.6u w=7u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=2.1p pd=14.6u as=2.1p ps=14.6u w=7u l=0.15u
.ends

.subckt sky130_rom_krom_pinv_dec_0 A Z vdd gnd w_956_n45#
X0 vdd A Z w_956_n45# sky130_fd_pr__pfet_01v8 ad=2.1p pd=14.6u as=2.1p ps=14.6u w=7u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.9p pd=6.6u as=0.9p ps=6.6u w=3u l=0.15u
.ends

.subckt sky130_rom_krom_pbuf_dec Z vdd vdd_uq0 gnd A sky130_rom_krom_pinv_dec_0_0/w_956_n45#
+ sky130_rom_krom_pinv_dec_1_0/w_1756_n45#
Xsky130_rom_krom_pinv_dec_1_0 sky130_rom_krom_pinv_dec_1_0/A Z vdd_uq0 sky130_rom_krom_pinv_dec_1_0/w_1756_n45#
+ gnd sky130_rom_krom_pinv_dec_1
Xsky130_rom_krom_pinv_dec_0_0 A sky130_rom_krom_pinv_dec_1_0/A vdd gnd sky130_rom_krom_pinv_dec_0_0/w_956_n45#
+ sky130_rom_krom_pinv_dec_0
.ends

.subckt sky130_rom_krom_rom_row_decode_wordline_buffer in_0 in_1 in_2 in_3 in_4 in_6
+ in_7 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd_uq0 in_5 vdd gnd
Xsky130_rom_krom_pbuf_dec_0 out_7 vdd vdd_uq0 gnd in_7 vdd vdd_uq0 sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_1 out_6 vdd vdd_uq0 gnd in_6 vdd vdd_uq0 sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_2 out_5 vdd vdd_uq0 gnd in_5 vdd vdd_uq0 sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_3 out_4 vdd vdd_uq0 gnd in_4 vdd vdd_uq0 sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_5 out_2 vdd vdd_uq0 gnd in_2 vdd vdd_uq0 sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_4 out_3 vdd vdd_uq0 gnd in_3 vdd vdd_uq0 sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_6 out_1 vdd vdd_uq0 gnd in_1 vdd vdd_uq0 sky130_rom_krom_pbuf_dec
Xsky130_rom_krom_pbuf_dec_7 out_0 vdd vdd_uq0 gnd in_0 vdd vdd_uq0 sky130_rom_krom_pbuf_dec
.ends

.subckt sky130_rom_krom_rom_row_decode A0 A1 A2 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6
+ wl_7 clk vdd_uq0 vdd_uq2 vdd_uq5 vdd_uq6 vdd vdd_uq1 precharge gnd
Xsky130_rom_krom_rom_row_decode_array_0 sky130_rom_krom_rom_row_decode_array_0/bl_0_0
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_1 sky130_rom_krom_rom_row_decode_array_0/bl_0_2
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_3 sky130_rom_krom_rom_row_decode_array_0/bl_0_4
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_5 sky130_rom_krom_rom_row_decode_array_0/bl_0_6
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_7 sky130_rom_krom_rom_row_decode_array_0/wl_0_1
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_2 sky130_rom_krom_rom_row_decode_array_0/wl_0_3
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_4 sky130_rom_krom_rom_row_decode_array_0/wl_0_5
+ gnd sky130_rom_krom_rom_row_decode_array_0/wl_0_0 vdd_uq0 precharge sky130_rom_krom_rom_row_decode_array
Xsky130_rom_krom_rom_address_control_array_0 A0 A1 A2 sky130_rom_krom_rom_row_decode_array_0/wl_0_5
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_3 sky130_rom_krom_rom_row_decode_array_0/wl_0_1
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_4 sky130_rom_krom_rom_row_decode_array_0/wl_0_2
+ clk vdd_uq1 gnd vdd vdd_uq2 sky130_rom_krom_rom_row_decode_array_0/wl_0_0 sky130_rom_krom_rom_address_control_array
Xsky130_rom_krom_rom_row_decode_wordline_buffer_0 sky130_rom_krom_rom_row_decode_array_0/bl_0_0
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_1 sky130_rom_krom_rom_row_decode_array_0/bl_0_2
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_3 sky130_rom_krom_rom_row_decode_array_0/bl_0_4
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_6 sky130_rom_krom_rom_row_decode_array_0/bl_0_7
+ wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 vdd_uq5 sky130_rom_krom_rom_row_decode_array_0/bl_0_5
+ vdd_uq6 gnd sky130_rom_krom_rom_row_decode_wordline_buffer
.ends

.subckt sky130_rom_krom_pinv_dec_4 A Z vdd gnd w_692_n45#
X0 vdd A Z w_692_n45# sky130_fd_pr__pfet_01v8 ad=1.5p pd=10.6u as=1.5p ps=10.6u w=5u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.504p pd=3.96u as=0.504p ps=3.96u w=1.68u l=0.15u
.ends

.subckt sky130_rom_krom_rom_output_buffer in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7
+ in_8 in_9 in_10 in_11 in_12 in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21
+ in_22 in_23 in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 out_0 out_1 out_2 out_3
+ out_4 out_5 out_6 out_7 out_8 out_9 out_10 out_11 out_12 out_13 out_14 out_15 out_16
+ out_17 out_18 out_19 out_20 out_21 out_22 out_23 out_24 out_25 out_26 out_27 out_28
+ out_29 out_30 out_31 gnd vdd
Xsky130_rom_krom_pinv_dec_4_20 in_11 out_11 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_31 in_0 out_0 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_10 in_21 out_21 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_21 in_10 out_10 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_11 in_20 out_20 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_12 in_19 out_19 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_22 in_9 out_9 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_23 in_8 out_8 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_13 in_18 out_18 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_24 in_7 out_7 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_14 in_17 out_17 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_25 in_6 out_6 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_15 in_16 out_16 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_26 in_5 out_5 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_16 in_15 out_15 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_27 in_4 out_4 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_17 in_14 out_14 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_28 in_3 out_3 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_18 in_13 out_13 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_29 in_2 out_2 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_19 in_12 out_12 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_0 in_31 out_31 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_1 in_30 out_30 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_2 in_29 out_29 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_3 in_28 out_28 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_4 in_27 out_27 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_5 in_26 out_26 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_6 in_25 out_25 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_7 in_24 out_24 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_8 in_23 out_23 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_9 in_22 out_22 vdd gnd vdd sky130_rom_krom_pinv_dec_4
Xsky130_rom_krom_pinv_dec_4_30 in_1 out_1 vdd gnd vdd sky130_rom_krom_pinv_dec_4
.ends

.subckt sky130_rom_krom_pinv_0 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.2886p pd=2.26u as=0.444p ps=4.16u w=0.74u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0.74u l=0.15u
X2 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0.756p pd=6.24u as=0.4914p ps=3.3u w=1.26u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26u l=0.15u
.ends

.subckt sky130_rom_krom_pinv_1 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=2.07p pd=13.38u as=2.07p ps=13.38u w=3u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X2 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=2.07p pd=13.38u as=2.07p ps=13.38u w=3u l=0.15u
X4 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X5 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
.ends

.subckt sky130_rom_krom_pinv A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.108p pd=1.32u as=0.108p ps=1.32u w=0.36u l=0.15u
X1 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.336p pd=2.84u as=0.336p ps=2.84u w=1.12u l=0.15u
.ends

.subckt sky130_rom_krom_rom_clock_driver A Z vdd gnd
Xsky130_rom_krom_pinv_0_0 sky130_rom_krom_pinv_0/Z sky130_rom_krom_pinv_1_0/A vdd
+ gnd sky130_rom_krom_pinv_0
Xsky130_rom_krom_pinv_1_0 sky130_rom_krom_pinv_1_0/A Z vdd gnd sky130_rom_krom_pinv_1
Xsky130_rom_krom_pinv_0 sky130_rom_krom_pinv_1/Z sky130_rom_krom_pinv_0/Z vdd gnd
+ sky130_rom_krom_pinv
Xsky130_rom_krom_pinv_1 A sky130_rom_krom_pinv_1/Z vdd gnd sky130_rom_krom_pinv
.ends

.subckt sky130_rom_krom_rom_control_nand A B Z vdd gnd w_n36_1262#
X0 a_144_51# A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.259p pd=2.18u as=0.222p ps=2.08u w=0.74u l=0.15u
X1 vdd B Z w_n36_1262# sky130_fd_pr__pfet_01v8 ad=0.672p pd=5.68u as=0.392p ps=2.94u w=1.12u l=0.15u
X2 Z A vdd w_n36_1262# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12u l=0.15u
X3 Z B a_144_51# gnd sky130_fd_pr__nfet_01v8 ad=0.222p pd=2.08u as=0p ps=0u w=0.74u l=0.15u
.ends

.subckt sky130_rom_krom_pinv_4 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=4.41p pd=26.94u as=4.41p ps=26.94u w=3u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X2 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X3 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=7.35p pd=42.94u as=7.35p ps=42.94u w=5u l=0.15u
X4 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X5 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X6 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X7 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X8 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X9 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X10 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X11 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X12 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X13 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
.ends

.subckt sky130_rom_krom_pinv_2 A Z vdd gnd
X0 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=1.2p pd=9.2u as=0.78p ps=4.78u w=2u l=0.15u
X1 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.4914p pd=3.3u as=0.756p ps=6.24u w=1.26u l=0.15u
X3 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26u l=0.15u
.ends

.subckt sky130_rom_krom_pinv_5 A Z vdd gnd
X0 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=19.5p pd=107.8u as=20.55p ps=118.22u w=5u l=0.15u
X1 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X2 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=20.55p pd=118.22u as=19.5p ps=107.8u w=5u l=0.15u
X3 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X4 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X5 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X6 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X7 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X8 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X9 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X10 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X11 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X12 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X13 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X14 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X15 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X16 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X17 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X18 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X19 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X20 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X21 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X22 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X23 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X24 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X25 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X26 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X27 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X28 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X29 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X30 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X31 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X32 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X33 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X34 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X35 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X36 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X37 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X38 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
X39 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5u l=0.15u
.ends

.subckt sky130_rom_krom_pinv_3 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=1.56p pd=9.56u as=1.98p ps=13.98u w=2u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=2.97p pd=19.98u as=2.34p ps=13.56u w=3u l=0.15u
X4 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X5 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X6 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X7 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
.ends

.subckt sky130_rom_krom_rom_precharge_driver A Z vdd gnd
Xsky130_rom_krom_pinv_4_0 sky130_rom_krom_pinv_4_0/A sky130_rom_krom_pinv_5_0/A vdd
+ gnd sky130_rom_krom_pinv_4
Xsky130_rom_krom_pinv_2_0 sky130_rom_krom_pinv_0/Z sky130_rom_krom_pinv_3_0/A vdd
+ gnd sky130_rom_krom_pinv_2
Xsky130_rom_krom_pinv_5_0 sky130_rom_krom_pinv_5_0/A Z vdd gnd sky130_rom_krom_pinv_5
Xsky130_rom_krom_pinv_3_0 sky130_rom_krom_pinv_3_0/A sky130_rom_krom_pinv_4_0/A vdd
+ gnd sky130_rom_krom_pinv_3
Xsky130_rom_krom_pinv_0 sky130_rom_krom_pinv_1/Z sky130_rom_krom_pinv_0/Z vdd gnd
+ sky130_rom_krom_pinv
Xsky130_rom_krom_pinv_1 sky130_rom_krom_pinv_2/Z sky130_rom_krom_pinv_1/Z vdd gnd
+ sky130_rom_krom_pinv
Xsky130_rom_krom_pinv_2 A sky130_rom_krom_pinv_2/Z vdd gnd sky130_rom_krom_pinv
.ends

.subckt sky130_rom_krom_rom_control_logic clk_in CS prechrg clk_out vdd gnd
Xsky130_rom_krom_rom_clock_driver_0 clk_in clk_out vdd gnd sky130_rom_krom_rom_clock_driver
Xsky130_rom_krom_rom_control_nand_0 CS clk_out sky130_rom_krom_rom_control_nand_0/Z
+ vdd gnd vdd sky130_rom_krom_rom_control_nand
Xsky130_rom_krom_rom_precharge_driver_0 sky130_rom_krom_rom_control_nand_0/Z prechrg
+ vdd gnd sky130_rom_krom_rom_precharge_driver
.ends

.subckt sky130_rom_krom_rom_column_mux bl bl_out sel gnd
X0 bl_out sel bl gnd sky130_fd_pr__nfet_01v8 ad=0.864p pd=6.36u as=0.864p ps=6.36u w=2.88u l=0.15u
.ends

.subckt sky130_rom_krom_rom_column_mux_array bl_0 bl_1 bl_3 bl_4 bl_6 bl_8 bl_9 bl_11
+ bl_15 bl_16 bl_17 bl_18 bl_19 bl_26 bl_27 bl_28 bl_29 bl_30 bl_37 bl_38 bl_39 bl_41
+ bl_48 bl_49 bl_59 bl_71 bl_74 bl_76 bl_79 bl_82 bl_85 bl_87 bl_90 bl_93 bl_98 bl_100
+ bl_101 bl_102 bl_104 bl_105 bl_106 bl_107 bl_109 bl_110 bl_112 bl_113 bl_115 bl_117
+ bl_118 bl_120 bl_121 bl_123 bl_124 bl_126 bl_128 bl_129 bl_130 bl_131 bl_132 bl_134
+ bl_135 bl_136 bl_137 bl_139 bl_140 bl_141 bl_142 bl_143 bl_145 bl_147 bl_148 bl_150
+ bl_151 bl_153 bl_154 bl_157 bl_158 bl_160 bl_161 bl_163 bl_164 bl_166 bl_168 bl_169
+ bl_170 bl_171 bl_172 bl_174 bl_175 bl_176 bl_177 bl_179 bl_182 bl_183 bl_184 bl_185
+ bl_187 bl_188 bl_189 bl_192 bl_193 bl_194 bl_195 bl_196 bl_197 bl_198 bl_199 bl_200
+ bl_203 bl_208 bl_211 bl_214 bl_216 bl_219 bl_222 bl_225 bl_227 bl_230 bl_233 bl_238
+ bl_241 bl_244 bl_248 bl_251 bl_254 sel_4 sel_5 bl_out_0 bl_out_1 bl_out_2 bl_out_3
+ bl_out_4 bl_out_5 bl_out_6 bl_out_7 bl_out_8 bl_out_9 bl_out_10 bl_out_11 bl_out_12
+ bl_out_13 bl_out_14 bl_out_15 bl_out_16 bl_out_17 bl_out_18 bl_out_19 bl_out_20
+ bl_out_21 bl_out_22 bl_out_23 bl_out_24 bl_out_25 bl_out_26 bl_out_27 bl_out_28
+ bl_out_29 bl_out_30 bl_out_31 bl_14 bl_22 bl_25 bl_33 bl_46 bl_44 bl_52 bl_55 bl_58
+ bl_66 bl_61 bl_69 bl_64 bl_190 bl_77 bl_72 bl_80 bl_206 bl_75 bl_201 bl_88 bl_83
+ bl_209 bl_204 bl_96 bl_91 bl_217 bl_212 bl_99 bl_94 bl_220 bl_215 bl_12 bl_246 bl_228
+ bl_223 bl_20 bl_236 bl_231 bl_249 bl_23 bl_239 bl_36 bl_252 bl_234 bl_31 bl_242
+ bl_255 bl_34 bl_245 bl_47 bl_42 bl_50 bl_45 bl_53 bl_56 bl_180 bl_67 bl_62 bl_70
+ bl_65 bl_191 bl_78 bl_73 bl_86 bl_81 bl_207 bl_202 bl_89 bl_84 bl_210 bl_7 bl_205
+ bl_97 bl_92 bl_2 bl_218 bl_213 bl_10 bl_95 bl_5 bl_226 bl_221 bl_108 bl_103 bl_13
+ bl_229 bl_247 bl_224 bl_116 bl_111 bl_21 bl_237 bl_250 bl_232 bl_119 bl_114 bl_24
+ bl_240 bl_235 bl_127 bl_253 bl_32 bl_122 bl_243 bl_40 bl_125 bl_35 bl_138 bl_133
+ bl_43 bl_146 bl_51 bl_149 bl_144 bl_54 bl_152 bl_156 bl_155 bl_159 bl_167 bl_162
+ sel_0 sel_7 sel_6 bl_57 bl_165 sel_1 bl_178 bl_173 gnd bl_60 bl_186 bl_181 bl_68
+ sel_3 bl_63 sel_2
Xsky130_rom_krom_rom_column_mux_110 bl_145 bl_out_18 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_121 bl_134 bl_out_16 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_132 bl_123 bl_out_15 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_143 bl_112 bl_out_14 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_154 bl_101 bl_out_12 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_198 bl_57 bl_out_7 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_187 bl_68 bl_out_8 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_176 bl_79 bl_out_9 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_165 bl_90 bl_out_11 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_100 bl_155 bl_out_19 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_111 bl_144 bl_out_18 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_122 bl_133 bl_out_16 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_133 bl_122 bl_out_15 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_144 bl_111 bl_out_13 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_155 bl_100 bl_out_12 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_199 bl_56 bl_out_7 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_188 bl_67 bl_out_8 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_177 bl_78 bl_out_9 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_166 bl_89 bl_out_11 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_101 bl_154 bl_out_19 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_112 bl_143 bl_out_17 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_123 bl_132 bl_out_16 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_134 bl_121 bl_out_15 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_145 bl_110 bl_out_13 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_156 bl_99 bl_out_12 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_189 bl_66 bl_out_8 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_178 bl_77 bl_out_9 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_167 bl_88 bl_out_11 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_102 bl_153 bl_out_19 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_113 bl_142 bl_out_17 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_124 bl_131 bl_out_16 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_135 bl_120 bl_out_15 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_146 bl_109 bl_out_13 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_157 bl_98 bl_out_12 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_179 bl_76 bl_out_9 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_168 bl_87 bl_out_10 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_103 bl_152 bl_out_19 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_114 bl_141 bl_out_17 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_125 bl_130 bl_out_16 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_136 bl_119 bl_out_14 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_147 bl_108 bl_out_13 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_158 bl_97 bl_out_12 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_169 bl_86 bl_out_10 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_104 bl_151 bl_out_18 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_115 bl_140 bl_out_17 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_126 bl_129 bl_out_16 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_137 bl_118 bl_out_14 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_148 bl_107 bl_out_13 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_159 bl_96 bl_out_12 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_90 bl_165 bl_out_20 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_105 bl_150 bl_out_18 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_116 bl_139 bl_out_17 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_127 bl_128 bl_out_16 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_138 bl_117 bl_out_14 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_149 bl_106 bl_out_13 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_80 bl_175 bl_out_21 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_91 bl_164 bl_out_20 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_106 bl_149 bl_out_18 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_117 bl_138 bl_out_17 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_128 bl_127 bl_out_15 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_139 bl_116 bl_out_14 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_70 bl_185 bl_out_23 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_81 bl_174 bl_out_21 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_92 bl_163 bl_out_20 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_107 bl_148 bl_out_18 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_118 bl_137 bl_out_17 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_129 bl_126 bl_out_15 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_60 bl_195 bl_out_24 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_71 bl_184 bl_out_23 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_82 bl_173 bl_out_21 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_93 bl_162 bl_out_20 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_108 bl_147 bl_out_18 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_119 bl_136 bl_out_17 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_50 bl_205 bl_out_25 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_61 bl_194 bl_out_24 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_72 bl_183 bl_out_22 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_83 bl_172 bl_out_21 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_94 bl_161 bl_out_20 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_109 bl_146 bl_out_18 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_40 bl_215 bl_out_26 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_51 bl_204 bl_out_25 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_62 bl_193 bl_out_24 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_73 bl_182 bl_out_22 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_84 bl_171 bl_out_21 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_95 bl_160 bl_out_20 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_30 bl_225 bl_out_28 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_41 bl_214 bl_out_26 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_52 bl_203 bl_out_25 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_63 bl_192 bl_out_24 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_74 bl_181 bl_out_22 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_85 bl_170 bl_out_21 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_96 bl_159 bl_out_19 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_250 bl_5 bl_out_0 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_20 bl_235 bl_out_29 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_31 bl_224 bl_out_28 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_42 bl_213 bl_out_26 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_53 bl_202 bl_out_25 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_64 bl_191 bl_out_23 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_75 bl_180 bl_out_22 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_86 bl_169 bl_out_21 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_97 bl_158 bl_out_19 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_251 bl_4 bl_out_0 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_240 bl_15 bl_out_1 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_10 bl_245 bl_out_30 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_21 bl_234 bl_out_29 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_32 bl_223 bl_out_27 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_43 bl_212 bl_out_26 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_54 bl_201 bl_out_25 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_65 bl_190 bl_out_23 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_76 bl_179 bl_out_22 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_87 bl_168 bl_out_21 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_98 bl_157 bl_out_19 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_252 bl_3 bl_out_0 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_241 bl_14 bl_out_1 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_230 bl_25 bl_out_3 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_11 bl_244 bl_out_30 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_22 bl_233 bl_out_29 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_33 bl_222 bl_out_27 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_44 bl_211 bl_out_26 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_55 bl_200 bl_out_25 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_66 bl_189 bl_out_23 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_77 bl_178 bl_out_22 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_88 bl_167 bl_out_20 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_99 bl_156 bl_out_19 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_253 bl_2 bl_out_0 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_242 bl_13 bl_out_1 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_231 bl_24 bl_out_3 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_220 bl_35 bl_out_4 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_12 bl_243 bl_out_30 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_23 bl_232 bl_out_29 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_34 bl_221 bl_out_27 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_45 bl_210 bl_out_26 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_56 bl_199 bl_out_24 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_67 bl_188 bl_out_23 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_78 bl_177 bl_out_22 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_89 bl_166 bl_out_20 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_254 bl_1 bl_out_0 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_243 bl_12 bl_out_1 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_232 bl_23 bl_out_2 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_221 bl_34 bl_out_4 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_210 bl_45 bl_out_5 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_13 bl_242 bl_out_30 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_24 bl_231 bl_out_28 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_35 bl_220 bl_out_27 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_46 bl_209 bl_out_26 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_57 bl_198 bl_out_24 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_68 bl_187 bl_out_23 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_79 bl_176 bl_out_22 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_255 bl_0 bl_out_0 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_244 bl_11 bl_out_1 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_233 bl_22 bl_out_2 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_222 bl_33 bl_out_4 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_211 bl_44 bl_out_5 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_200 bl_55 bl_out_6 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_14 bl_241 bl_out_30 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_25 bl_230 bl_out_28 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_36 bl_219 bl_out_27 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_47 bl_208 bl_out_26 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_58 bl_197 bl_out_24 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_69 bl_186 bl_out_23 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_245 bl_10 bl_out_1 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_234 bl_21 bl_out_2 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_223 bl_32 bl_out_4 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_212 bl_43 bl_out_5 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_201 bl_54 bl_out_6 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_15 bl_240 bl_out_30 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_26 bl_229 bl_out_28 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_37 bl_218 bl_out_27 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_48 bl_207 bl_out_25 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_59 bl_196 bl_out_24 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_246 bl_9 bl_out_1 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_235 bl_20 bl_out_2 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_224 bl_31 bl_out_3 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_213 bl_42 bl_out_5 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_202 bl_53 bl_out_6 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_16 bl_239 bl_out_29 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_27 bl_228 bl_out_28 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_38 bl_217 bl_out_27 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_49 bl_206 bl_out_25 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_17 bl_238 bl_out_29 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_28 bl_227 bl_out_28 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_39 bl_216 bl_out_27 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_247 bl_8 bl_out_1 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_236 bl_19 bl_out_2 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_225 bl_30 bl_out_3 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_214 bl_41 bl_out_5 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_203 bl_52 bl_out_6 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_248 bl_7 bl_out_0 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_237 bl_18 bl_out_2 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_226 bl_29 bl_out_3 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_215 bl_40 bl_out_5 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_204 bl_51 bl_out_6 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_18 bl_237 bl_out_29 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_29 bl_226 bl_out_28 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_249 bl_6 bl_out_0 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_238 bl_17 bl_out_2 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_227 bl_28 bl_out_3 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_216 bl_39 bl_out_4 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_205 bl_50 bl_out_6 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_19 bl_236 bl_out_29 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_239 bl_16 bl_out_2 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_228 bl_27 bl_out_3 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_217 bl_38 bl_out_4 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_206 bl_49 bl_out_6 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_229 bl_26 bl_out_3 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_218 bl_37 bl_out_4 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_207 bl_48 bl_out_6 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_219 bl_36 bl_out_4 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_208 bl_47 bl_out_5 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_0 bl_255 bl_out_31 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_209 bl_46 bl_out_5 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_1 bl_254 bl_out_31 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_2 bl_253 bl_out_31 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_190 bl_65 bl_out_8 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_3 bl_252 bl_out_31 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_191 bl_64 bl_out_8 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_180 bl_75 bl_out_9 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_4 bl_251 bl_out_31 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_192 bl_63 bl_out_7 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_181 bl_74 bl_out_9 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_170 bl_85 bl_out_10 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_5 bl_250 bl_out_31 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_193 bl_62 bl_out_7 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_182 bl_73 bl_out_9 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_171 bl_84 bl_out_10 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_160 bl_95 bl_out_11 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_6 bl_249 bl_out_31 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_150 bl_105 bl_out_13 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_194 bl_61 bl_out_7 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_183 bl_72 bl_out_9 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_172 bl_83 bl_out_10 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_161 bl_94 bl_out_11 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_7 bl_248 bl_out_31 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_140 bl_115 bl_out_14 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_151 bl_104 bl_out_13 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_195 bl_60 bl_out_7 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_184 bl_71 bl_out_8 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_173 bl_82 bl_out_10 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_162 bl_93 bl_out_11 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_8 bl_247 bl_out_30 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_130 bl_125 bl_out_15 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_141 bl_114 bl_out_14 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_152 bl_103 bl_out_12 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_196 bl_59 bl_out_7 sel_3 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_185 bl_70 bl_out_8 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_174 bl_81 bl_out_10 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_163 bl_92 bl_out_11 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_9 bl_246 bl_out_30 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_120 bl_135 bl_out_16 sel_7 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_131 bl_124 bl_out_15 sel_4 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_142 bl_113 bl_out_14 sel_1 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_153 bl_102 bl_out_12 sel_6 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_197 bl_58 bl_out_7 sel_2 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_186 bl_69 bl_out_8 sel_5 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_175 bl_80 bl_out_10 sel_0 gnd sky130_rom_krom_rom_column_mux
Xsky130_rom_krom_rom_column_mux_164 bl_91 bl_out_11 sel_3 gnd sky130_rom_krom_rom_column_mux
.ends

.subckt sky130_rom_krom_rom_precharge_array pre_bl0_out pre_bl1_out pre_bl3_out pre_bl6_out
+ pre_bl8_out pre_bl9_out pre_bl10_out pre_bl13_out pre_bl15_out pre_bl16_out pre_bl22_out
+ pre_bl24_out pre_bl26_out pre_bl29_out pre_bl31_out pre_bl33_out pre_bl34_out pre_bl36_out
+ pre_bl38_out pre_bl40_out pre_bl43_out pre_bl44_out pre_bl46_out pre_bl47_out pre_bl52_out
+ pre_bl53_out pre_bl54_out pre_bl56_out pre_bl58_out pre_bl59_out pre_bl60_out pre_bl61_out
+ pre_bl62_out pre_bl65_out pre_bl68_out pre_bl70_out pre_bl71_out pre_bl74_out pre_bl77_out
+ pre_bl79_out pre_bl80_out pre_bl81_out pre_bl83_out pre_bl86_out pre_bl88_out pre_bl89_out
+ pre_bl90_out pre_bl91_out pre_bl95_out pre_bl97_out pre_bl98_out pre_bl102_out pre_bl104_out
+ pre_bl106_out pre_bl109_out pre_bl111_out pre_bl113_out pre_bl114_out pre_bl116_out
+ pre_bl118_out pre_bl120_out pre_bl123_out pre_bl124_out pre_bl127_out pre_bl132_out
+ pre_bl133_out pre_bl134_out pre_bl139_out pre_bl141_out pre_bl142_out pre_bl143_out
+ pre_bl144_out pre_bl145_out pre_bl148_out pre_bl150_out pre_bl151_out pre_bl153_out
+ pre_bl156_out pre_bl157_out pre_bl160_out pre_bl162_out pre_bl163_out pre_bl165_out
+ pre_bl166_out pre_bl167_out pre_bl172_out pre_bl174_out pre_bl175_out pre_bl177_out
+ pre_bl181_out pre_bl183_out pre_bl184_out pre_bl185_out pre_bl186_out pre_bl190_out
+ pre_bl192_out pre_bl193_out pre_bl195_out pre_bl196_out pre_bl202_out pre_bl204_out
+ pre_bl206_out pre_bl209_out pre_bl211_out pre_bl213_out pre_bl214_out pre_bl215_out
+ pre_bl218_out pre_bl220_out pre_bl222_out pre_bl223_out pre_bl224_out pre_bl227_out
+ pre_bl229_out pre_bl232_out pre_bl233_out pre_bl234_out pre_bl239_out pre_bl241_out
+ pre_bl242_out pre_bl243_out pre_bl245_out pre_bl248_out pre_bl250_out pre_bl251_out
+ pre_bl252_out pre_bl254_out gate pre_bl197_out pre_bl158_out pre_bl188_out pre_bl146_out
+ pre_bl72_out pre_bl216_out pre_bl179_out pre_bl45_out pre_bl125_out pre_bl27_out
+ pre_bl107_out pre_bl155_out pre_bl20_out pre_bl137_out pre_bl100_out pre_bl50_out
+ pre_bl63_out pre_bl130_out pre_bl93_out pre_bl225_out pre_bl207_out pre_bl170_out
+ pre_bl237_out pre_bl200_out pre_bl246_out pre_bl18_out pre_bl230_out pre_bl48_out
+ pre_bl11_out pre_bl128_out pre_bl41_out pre_bl4_out pre_bl121_out pre_bl168_out
+ pre_bl84_out pre_bl66_out pre_bl198_out pre_bl161_out pre_bl255_out pre_bl96_out
+ pre_bl228_out pre_bl191_out pre_bl126_out pre_bl39_out pre_bl221_out pre_bl2_out
+ pre_bl119_out pre_bl82_out pre_bl32_out pre_bl149_out pre_bl112_out pre_bl244_out
+ pre_bl75_out pre_bl159_out pre_bl25_out pre_bl253_out pre_bl226_out pre_bl57_out
+ pre_bl189_out pre_bl105_out pre_bl7_out pre_bl55_out pre_bl87_out pre_bl37_out pre_bl135_out
+ pre_bl219_out pre_bl182_out pre_bl117_out pre_bl212_out pre_bl30_out pre_bl147_out
+ pre_bl110_out pre_bl73_out pre_bl205_out pre_bl23_out pre_bl140_out pre_bl187_out
+ pre_bl103_out pre_bl235_out pre_bl217_out pre_bl180_out pre_bl78_out pre_bl210_out
+ pre_bl28_out pre_bl173_out pre_bl108_out pre_bl240_out pre_bl203_out pre_bl249_out
+ pre_bl21_out pre_bl138_out pre_bl101_out pre_bl51_out pre_bl64_out pre_bl14_out
+ pre_bl131_out pre_bl178_out pre_bl94_out pre_bl76_out pre_bl208_out pre_bl171_out
+ pre_bl238_out pre_bl154_out pre_bl69_out pre_bl19_out pre_bl201_out pre_bl247_out
+ pre_bl136_out pre_bl164_out pre_bl99_out pre_bl231_out pre_bl49_out pre_bl194_out
+ pre_bl12_out pre_bl129_out pre_bl176_out pre_bl92_out pre_bl42_out pre_bl5_out pre_bl122_out
+ pre_bl85_out pre_bl169_out pre_bl35_out pre_bl236_out pre_bl152_out pre_bl67_out
+ vdd pre_bl199_out pre_bl115_out pre_bl17_out
Xsky130_rom_krom_precharge_cell_2 pre_bl253_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_209 pre_bl46_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_90 pre_bl165_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_3 pre_bl252_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_80 pre_bl175_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_91 pre_bl164_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_190 pre_bl65_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_4 pre_bl251_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_70 pre_bl185_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_81 pre_bl174_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_92 pre_bl163_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_191 pre_bl64_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_180 pre_bl75_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_5 pre_bl250_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_60 pre_bl195_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_71 pre_bl184_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_82 pre_bl173_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_93 pre_bl162_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_6 pre_bl249_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_170 pre_bl85_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_192 pre_bl63_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_181 pre_bl74_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_50 pre_bl205_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_61 pre_bl194_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_72 pre_bl183_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_83 pre_bl172_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_94 pre_bl161_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_160 pre_bl95_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_193 pre_bl62_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_182 pre_bl73_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_171 pre_bl84_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_7 pre_bl248_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_40 pre_bl215_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_51 pre_bl204_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_62 pre_bl193_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_73 pre_bl182_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_84 pre_bl171_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_95 pre_bl160_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_8 pre_bl247_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_150 pre_bl105_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_161 pre_bl94_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_194 pre_bl61_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_183 pre_bl72_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_172 pre_bl83_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_30 pre_bl225_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_41 pre_bl214_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_52 pre_bl203_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_63 pre_bl192_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_74 pre_bl181_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_85 pre_bl170_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_96 pre_bl159_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_140 pre_bl115_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_151 pre_bl104_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_162 pre_bl93_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_195 pre_bl60_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_184 pre_bl71_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_173 pre_bl82_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_9 pre_bl246_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_20 pre_bl235_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_31 pre_bl224_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_42 pre_bl213_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_53 pre_bl202_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_64 pre_bl191_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_75 pre_bl180_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_86 pre_bl169_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_97 pre_bl158_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_130 pre_bl125_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_141 pre_bl114_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_152 pre_bl103_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_163 pre_bl92_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_196 pre_bl59_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_185 pre_bl70_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_174 pre_bl81_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_10 pre_bl245_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_21 pre_bl234_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_32 pre_bl223_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_43 pre_bl212_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_54 pre_bl201_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_65 pre_bl190_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_76 pre_bl179_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_87 pre_bl168_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_98 pre_bl157_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_120 pre_bl135_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_131 pre_bl124_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_142 pre_bl113_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_153 pre_bl102_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_164 pre_bl91_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_197 pre_bl58_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_186 pre_bl69_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_175 pre_bl80_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_11 pre_bl244_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_22 pre_bl233_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_33 pre_bl222_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_44 pre_bl211_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_55 pre_bl200_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_66 pre_bl189_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_77 pre_bl178_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_88 pre_bl167_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_99 pre_bl156_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_110 pre_bl145_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_121 pre_bl134_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_132 pre_bl123_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_143 pre_bl112_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_154 pre_bl101_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_165 pre_bl90_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_198 pre_bl57_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_187 pre_bl68_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_176 pre_bl79_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_12 pre_bl243_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_23 pre_bl232_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_34 pre_bl221_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_45 pre_bl210_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_56 pre_bl199_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_67 pre_bl188_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_78 pre_bl177_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_89 pre_bl166_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_100 pre_bl155_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_111 pre_bl144_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_122 pre_bl133_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_133 pre_bl122_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_144 pre_bl111_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_155 pre_bl100_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_166 pre_bl89_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_199 pre_bl56_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_188 pre_bl67_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_177 pre_bl78_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_13 pre_bl242_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_24 pre_bl231_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_35 pre_bl220_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_46 pre_bl209_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_57 pre_bl198_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_68 pre_bl187_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_79 pre_bl176_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_101 pre_bl154_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_112 pre_bl143_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_123 pre_bl132_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_134 pre_bl121_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_145 pre_bl110_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_156 pre_bl99_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_167 pre_bl88_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_189 pre_bl66_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_178 pre_bl77_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_14 pre_bl241_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_25 pre_bl230_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_36 pre_bl219_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_47 pre_bl208_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_58 pre_bl197_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_69 pre_bl186_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_102 pre_bl153_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_113 pre_bl142_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_124 pre_bl131_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_135 pre_bl120_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_146 pre_bl109_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_157 pre_bl98_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_168 pre_bl87_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_179 pre_bl76_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_15 pre_bl240_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_26 pre_bl229_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_37 pre_bl218_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_48 pre_bl207_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_59 pre_bl196_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_103 pre_bl152_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_114 pre_bl141_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_125 pre_bl130_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_136 pre_bl119_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_147 pre_bl108_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_158 pre_bl97_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_169 pre_bl86_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_16 pre_bl239_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_27 pre_bl228_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_38 pre_bl217_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_49 pre_bl206_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_104 pre_bl151_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_115 pre_bl140_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_126 pre_bl129_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_137 pre_bl118_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_148 pre_bl107_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_159 pre_bl96_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_17 pre_bl238_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_28 pre_bl227_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_39 pre_bl216_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_105 pre_bl150_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_116 pre_bl139_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_127 pre_bl128_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_138 pre_bl117_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_149 pre_bl106_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_18 pre_bl237_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_29 pre_bl226_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_106 pre_bl149_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_117 pre_bl138_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_128 pre_bl127_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_139 pre_bl116_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_19 pre_bl236_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_107 pre_bl148_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_118 pre_bl137_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_129 pre_bl126_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_108 pre_bl147_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_119 pre_bl136_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_109 pre_bl146_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_250 pre_bl5_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_251 pre_bl4_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_240 pre_bl15_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_252 pre_bl3_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_241 pre_bl14_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_230 pre_bl25_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_253 pre_bl2_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_242 pre_bl13_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_231 pre_bl24_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_220 pre_bl35_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_254 pre_bl1_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_243 pre_bl12_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_232 pre_bl23_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_221 pre_bl34_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_210 pre_bl45_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_255 pre_bl0_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_244 pre_bl11_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_233 pre_bl22_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_222 pre_bl33_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_211 pre_bl44_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_200 pre_bl55_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_245 pre_bl10_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_234 pre_bl21_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_223 pre_bl32_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_212 pre_bl43_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_201 pre_bl54_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_246 pre_bl9_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_235 pre_bl20_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_224 pre_bl31_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_213 pre_bl42_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_202 pre_bl53_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_247 pre_bl8_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_236 pre_bl19_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_225 pre_bl30_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_214 pre_bl41_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_203 pre_bl52_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_248 pre_bl7_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_237 pre_bl18_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_226 pre_bl29_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_215 pre_bl40_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_204 pre_bl51_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_249 pre_bl6_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_238 pre_bl17_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_227 pre_bl28_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_216 pre_bl39_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_205 pre_bl50_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_239 pre_bl16_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_228 pre_bl27_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_217 pre_bl38_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_206 pre_bl49_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_0 pre_bl255_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_229 pre_bl26_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_218 pre_bl37_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_207 pre_bl48_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_1 pre_bl254_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_219 pre_bl36_out gate vdd sky130_rom_krom_precharge_cell
Xsky130_rom_krom_precharge_cell_208 pre_bl47_out gate vdd sky130_rom_krom_precharge_cell
.ends

.subckt sky130_rom_krom_rom_base_array bl_0_0 bl_0_1 bl_0_2 bl_0_3 bl_0_4 bl_0_5 bl_0_6
+ bl_0_7 bl_0_8 bl_0_9 bl_0_10 bl_0_11 bl_0_12 bl_0_13 bl_0_14 bl_0_16 bl_0_17 bl_0_18
+ bl_0_19 bl_0_20 bl_0_21 bl_0_22 bl_0_23 bl_0_24 bl_0_25 bl_0_26 bl_0_27 bl_0_28
+ bl_0_29 bl_0_30 bl_0_31 bl_0_32 bl_0_33 bl_0_34 bl_0_35 bl_0_36 bl_0_37 bl_0_38
+ bl_0_39 bl_0_40 bl_0_41 bl_0_42 bl_0_43 bl_0_44 bl_0_45 bl_0_46 bl_0_47 bl_0_48
+ bl_0_49 bl_0_50 bl_0_51 bl_0_52 bl_0_53 bl_0_54 bl_0_55 bl_0_56 bl_0_57 bl_0_58
+ bl_0_59 bl_0_60 bl_0_61 bl_0_62 bl_0_63 bl_0_64 bl_0_65 bl_0_66 bl_0_67 bl_0_68
+ bl_0_69 bl_0_70 bl_0_71 bl_0_72 bl_0_73 bl_0_74 bl_0_75 bl_0_76 bl_0_77 bl_0_78
+ bl_0_79 bl_0_80 bl_0_81 bl_0_82 bl_0_83 bl_0_84 bl_0_85 bl_0_86 bl_0_87 bl_0_88
+ bl_0_89 bl_0_90 bl_0_91 bl_0_92 bl_0_93 bl_0_94 bl_0_95 bl_0_96 bl_0_97 bl_0_98
+ bl_0_99 bl_0_100 bl_0_101 bl_0_102 bl_0_103 bl_0_104 bl_0_105 bl_0_106 bl_0_107
+ bl_0_108 bl_0_109 bl_0_110 bl_0_111 bl_0_112 bl_0_113 bl_0_114 bl_0_115 bl_0_116
+ bl_0_117 bl_0_118 bl_0_119 bl_0_120 bl_0_121 bl_0_122 bl_0_123 bl_0_124 bl_0_125
+ bl_0_126 bl_0_127 bl_0_128 bl_0_129 bl_0_130 bl_0_131 bl_0_132 bl_0_133 bl_0_134
+ bl_0_135 bl_0_136 bl_0_137 bl_0_138 bl_0_139 bl_0_140 bl_0_141 bl_0_142 bl_0_143
+ bl_0_144 bl_0_145 bl_0_146 bl_0_147 bl_0_148 bl_0_149 bl_0_150 bl_0_151 bl_0_152
+ bl_0_153 bl_0_154 bl_0_155 bl_0_156 bl_0_157 bl_0_158 bl_0_159 bl_0_160 bl_0_161
+ bl_0_162 bl_0_163 bl_0_164 bl_0_165 bl_0_166 bl_0_167 bl_0_168 bl_0_169 bl_0_170
+ bl_0_171 bl_0_172 bl_0_173 bl_0_174 bl_0_175 bl_0_176 bl_0_177 bl_0_178 bl_0_179
+ bl_0_180 bl_0_181 bl_0_182 bl_0_183 bl_0_184 bl_0_185 bl_0_186 bl_0_187 bl_0_188
+ bl_0_189 bl_0_190 bl_0_191 bl_0_192 bl_0_193 bl_0_194 bl_0_195 bl_0_196 bl_0_197
+ bl_0_198 bl_0_199 bl_0_200 bl_0_201 bl_0_202 bl_0_203 bl_0_204 bl_0_205 bl_0_206
+ bl_0_207 bl_0_208 bl_0_209 bl_0_210 bl_0_211 bl_0_212 bl_0_213 bl_0_214 bl_0_215
+ bl_0_216 bl_0_217 bl_0_218 bl_0_219 bl_0_220 bl_0_221 bl_0_222 bl_0_223 bl_0_224
+ bl_0_225 bl_0_226 bl_0_227 bl_0_228 bl_0_229 bl_0_230 bl_0_231 bl_0_232 bl_0_233
+ bl_0_234 bl_0_235 bl_0_236 bl_0_237 bl_0_238 bl_0_239 bl_0_240 bl_0_241 bl_0_242
+ bl_0_243 bl_0_244 bl_0_245 bl_0_246 bl_0_247 bl_0_248 bl_0_249 bl_0_250 bl_0_251
+ bl_0_252 bl_0_253 bl_0_254 bl_0_255 wl_0_1 wl_0_2 wl_0_4 wl_0_5 wl_0_6 wl_0_7 gnd
+ gnd_uq0 bl_0_15 wl_0_0 precharge wl_0_3 vdd
Xsky130_rom_krom_rom_base_one_cell_998 wl_0_1 sky130_rom_krom_rom_base_one_cell_998/D
+ sky130_rom_krom_rom_base_one_cell_998/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_987 wl_0_2 sky130_rom_krom_rom_base_one_cell_987/D
+ sky130_rom_krom_rom_base_one_cell_987/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_976 wl_0_2 sky130_rom_krom_rom_base_one_cell_976/D
+ bl_0_34 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_965 wl_0_2 sky130_rom_krom_rom_base_one_cell_965/D
+ sky130_rom_krom_rom_base_one_cell_965/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_954 wl_0_2 sky130_rom_krom_rom_base_one_cell_954/D
+ sky130_rom_krom_rom_base_one_cell_954/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_943 wl_0_2 sky130_rom_krom_rom_base_one_cell_943/D
+ bl_0_88 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_932 wl_0_2 sky130_rom_krom_rom_base_one_cell_932/D
+ sky130_rom_krom_rom_base_one_cell_932/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_921 wl_0_2 sky130_rom_krom_rom_base_one_cell_921/D
+ sky130_rom_krom_rom_base_one_cell_921/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_910 wl_0_2 sky130_rom_krom_rom_base_one_cell_910/D
+ sky130_rom_krom_rom_base_one_cell_910/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_206 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_99/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_217 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_369/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_228 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_502/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_239 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_379/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_260 wl_0_5 sky130_rom_krom_rom_base_one_cell_629/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_271 wl_0_5 sky130_rom_krom_rom_base_one_cell_24/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_282 wl_0_5 sky130_rom_krom_rom_base_one_cell_646/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_293 wl_0_5 sky130_rom_krom_rom_base_one_cell_61/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1085 wl_0_1 sky130_rom_krom_rom_base_one_cell_704/S
+ bl_0_82 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1096 wl_0_1 sky130_rom_krom_rom_base_one_cell_837/S
+ sky130_rom_krom_rom_base_one_cell_1224/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1074 wl_0_1 sky130_rom_krom_rom_base_one_cell_934/S
+ sky130_rom_krom_rom_base_one_cell_1197/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1063 wl_0_1 sky130_rom_krom_rom_base_one_cell_928/S
+ bl_0_120 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1052 wl_0_1 sky130_rom_krom_rom_base_one_cell_445/S
+ sky130_rom_krom_rom_base_one_cell_1175/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1041 wl_0_1 sky130_rom_krom_rom_base_one_cell_437/S
+ bl_0_161 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1030 wl_0_1 sky130_rom_krom_rom_base_one_cell_900/S
+ sky130_rom_krom_rom_base_one_cell_1154/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_50 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_50/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_61 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_61/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_72 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_72/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_83 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_83/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_94 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_94/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_740 wl_0_4 sky130_rom_krom_rom_base_one_cell_740/D
+ sky130_rom_krom_rom_base_one_cell_740/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_795 wl_0_3 sky130_rom_krom_rom_base_zero_cell_47/S
+ bl_0_152 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_784 wl_0_3 sky130_rom_krom_rom_base_one_cell_784/D
+ sky130_rom_krom_rom_base_one_cell_784/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_773 wl_0_3 sky130_rom_krom_rom_base_one_cell_773/D
+ sky130_rom_krom_rom_base_one_cell_894/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_762 wl_0_3 sky130_rom_krom_rom_base_one_cell_762/D
+ sky130_rom_krom_rom_base_one_cell_884/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_751 wl_0_3 sky130_rom_krom_rom_base_one_cell_751/D
+ bl_0_240 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1051 wl_0_0 bl_0_5 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1040 wl_0_0 bl_0_32 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_570 wl_0_5 sky130_rom_krom_rom_base_zero_cell_64/S
+ sky130_rom_krom_rom_base_one_cell_813/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_581 wl_0_5 sky130_rom_krom_rom_base_zero_cell_73/S
+ sky130_rom_krom_rom_base_one_cell_696/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_592 wl_0_5 sky130_rom_krom_rom_base_one_cell_592/D
+ sky130_rom_krom_rom_base_one_cell_952/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_804 wl_0_1 bl_0_248 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_859 wl_0_1 bl_0_129 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_848 wl_0_1 bl_0_150 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_837 wl_0_1 sky130_rom_krom_rom_base_one_cell_664/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_826 wl_0_1 bl_0_200 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_815 wl_0_1 bl_0_227 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_656 wl_0_3 sky130_rom_krom_rom_base_one_cell_979/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_645 wl_0_3 sky130_rom_krom_rom_base_one_cell_964/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_634 wl_0_3 sky130_rom_krom_rom_base_one_cell_956/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_623 wl_0_3 sky130_rom_krom_rom_base_zero_cell_75/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_612 wl_0_3 sky130_rom_krom_rom_base_one_cell_932/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_601 wl_0_3 sky130_rom_krom_rom_base_one_cell_563/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_689 wl_0_2 bl_0_219 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_678 wl_0_2 sky130_rom_krom_rom_base_one_cell_995/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_667 wl_0_3 bl_0_10 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1201 wl_0_0 sky130_rom_krom_rom_base_one_cell_1201/D
+ bl_0_94 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1245 wl_0_0 sky130_rom_krom_rom_base_one_cell_1245/D
+ bl_0_7 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1234 wl_0_0 sky130_rom_krom_rom_base_one_cell_851/S
+ bl_0_26 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1223 wl_0_0 sky130_rom_krom_rom_base_one_cell_962/S
+ bl_0_55 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1212 wl_0_0 sky130_rom_krom_rom_base_one_cell_952/S
+ bl_0_74 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_497 wl_0_4 bl_0_73 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_486 wl_0_4 sky130_rom_krom_rom_base_one_cell_820/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_475 wl_0_4 sky130_rom_krom_rom_base_one_cell_809/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_464 wl_0_4 sky130_rom_krom_rom_base_one_cell_804/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_453 wl_0_4 sky130_rom_krom_rom_base_zero_cell_47/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_442 wl_0_4 sky130_rom_krom_rom_base_one_cell_905/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_431 wl_0_4 sky130_rom_krom_rom_base_one_cell_62/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_420 wl_0_4 sky130_rom_krom_rom_base_one_cell_528/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_922 wl_0_2 sky130_rom_krom_rom_base_one_cell_922/D
+ sky130_rom_krom_rom_base_one_cell_922/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_911 wl_0_2 sky130_rom_krom_rom_base_one_cell_911/D
+ sky130_rom_krom_rom_base_one_cell_911/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_900 wl_0_2 sky130_rom_krom_rom_base_one_cell_900/D
+ sky130_rom_krom_rom_base_one_cell_900/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_999 wl_0_1 sky130_rom_krom_rom_base_one_cell_999/D
+ sky130_rom_krom_rom_base_one_cell_999/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_988 wl_0_2 sky130_rom_krom_rom_base_one_cell_988/D
+ sky130_rom_krom_rom_base_one_cell_988/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_977 wl_0_2 sky130_rom_krom_rom_base_one_cell_977/D
+ bl_0_33 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_966 wl_0_2 sky130_rom_krom_rom_base_one_cell_966/D
+ bl_0_47 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_955 wl_0_2 sky130_rom_krom_rom_base_one_cell_955/D
+ sky130_rom_krom_rom_base_one_cell_955/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_944 wl_0_2 sky130_rom_krom_rom_base_one_cell_944/D
+ bl_0_87 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_933 wl_0_2 sky130_rom_krom_rom_base_one_cell_933/D
+ sky130_rom_krom_rom_base_one_cell_933/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_207 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_601/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1053 wl_0_1 sky130_rom_krom_rom_base_one_cell_679/S
+ sky130_rom_krom_rom_base_one_cell_1176/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1042 wl_0_1 sky130_rom_krom_rom_base_one_cell_912/S
+ sky130_rom_krom_rom_base_one_cell_1168/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1031 wl_0_1 sky130_rom_krom_rom_base_one_cell_901/S
+ bl_0_185 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1020 wl_0_1 sky130_rom_krom_rom_base_one_cell_888/S
+ bl_0_203 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_218 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_496/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_229 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_851/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_250 wl_0_6 sky130_rom_krom_rom_base_one_cell_619/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_261 wl_0_5 sky130_rom_krom_rom_base_one_cell_630/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_272 wl_0_5 sky130_rom_krom_rom_base_one_cell_637/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_283 wl_0_5 sky130_rom_krom_rom_base_one_cell_762/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_294 wl_0_5 sky130_rom_krom_rom_base_one_cell_62/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1086 wl_0_1 sky130_rom_krom_rom_base_one_cell_829/S
+ bl_0_78 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1097 wl_0_1 sky130_rom_krom_rom_base_one_cell_838/S
+ bl_0_52 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1075 wl_0_1 sky130_rom_krom_rom_base_one_cell_818/S
+ sky130_rom_krom_rom_base_one_cell_1198/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1064 wl_0_1 sky130_rom_krom_rom_base_one_cell_684/S
+ bl_0_119 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_40 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_40/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_51 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_51/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_62 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_62/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_73 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_73/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_84 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_84/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_95 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_95/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_763 wl_0_3 sky130_rom_krom_rom_base_one_cell_763/D
+ bl_0_209 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_752 wl_0_3 sky130_rom_krom_rom_base_one_cell_752/D
+ sky130_rom_krom_rom_base_one_cell_999/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_741 wl_0_3 sky130_rom_krom_rom_base_one_cell_741/D
+ sky130_rom_krom_rom_base_one_cell_741/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_730 wl_0_4 sky130_rom_krom_rom_base_one_cell_730/D
+ sky130_rom_krom_rom_base_one_cell_850/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_796 wl_0_3 sky130_rom_krom_rom_base_one_cell_796/D
+ sky130_rom_krom_rom_base_one_cell_796/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_785 wl_0_3 sky130_rom_krom_rom_base_one_cell_785/D
+ sky130_rom_krom_rom_base_one_cell_785/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_774 wl_0_3 sky130_rom_krom_rom_base_one_cell_774/D
+ sky130_rom_krom_rom_base_one_cell_895/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1030 wl_0_0 bl_0_47 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1052 wl_0_0 bl_0_4 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1041 wl_0_0 bl_0_31 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_560 wl_0_5 sky130_rom_krom_rom_base_zero_cell_53/S
+ sky130_rom_krom_rom_base_one_cell_920/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_571 wl_0_5 sky130_rom_krom_rom_base_one_cell_571/D
+ sky130_rom_krom_rom_base_one_cell_688/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_593 wl_0_5 sky130_rom_krom_rom_base_one_cell_593/D
+ sky130_rom_krom_rom_base_one_cell_833/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_582 wl_0_5 sky130_rom_krom_rom_base_one_cell_582/D
+ sky130_rom_krom_rom_base_one_cell_820/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_838 wl_0_1 bl_0_173 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_827 wl_0_1 sky130_rom_krom_rom_base_one_cell_891/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_816 wl_0_1 bl_0_225 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_805 wl_0_1 bl_0_247 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_390 wl_0_6 sky130_rom_krom_rom_base_one_cell_390/D
+ sky130_rom_krom_rom_base_one_cell_512/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_849 wl_0_1 bl_0_148 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_679 wl_0_2 sky130_rom_krom_rom_base_one_cell_997/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_668 wl_0_3 sky130_rom_krom_rom_base_one_cell_988/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_657 wl_0_3 sky130_rom_krom_rom_base_one_cell_609/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_646 wl_0_3 sky130_rom_krom_rom_base_one_cell_965/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_635 wl_0_3 sky130_rom_krom_rom_base_one_cell_957/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_624 wl_0_3 sky130_rom_krom_rom_base_one_cell_945/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_613 wl_0_3 bl_0_106 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_602 wl_0_3 sky130_rom_krom_rom_base_one_cell_327/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1202 wl_0_0 sky130_rom_krom_rom_base_one_cell_1202/D
+ bl_0_93 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1235 wl_0_0 sky130_rom_krom_rom_base_one_cell_1235/D
+ bl_0_25 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1224 wl_0_0 sky130_rom_krom_rom_base_one_cell_1224/D
+ bl_0_54 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1213 wl_0_0 sky130_rom_krom_rom_base_one_cell_1213/D
+ bl_0_69 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1246 wl_0_0 sky130_rom_krom_rom_base_one_cell_1246/D
+ bl_0_6 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_498 wl_0_4 bl_0_72 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_487 wl_0_4 sky130_rom_krom_rom_base_one_cell_940/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_476 wl_0_4 bl_0_115 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_465 wl_0_4 sky130_rom_krom_rom_base_one_cell_561/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_454 wl_0_4 sky130_rom_krom_rom_base_one_cell_797/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_443 wl_0_4 sky130_rom_krom_rom_base_one_cell_789/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_432 wl_0_4 sky130_rom_krom_rom_base_one_cell_775/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_421 wl_0_4 bl_0_208 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_410 wl_0_4 sky130_rom_krom_rom_base_one_cell_755/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_956 wl_0_2 sky130_rom_krom_rom_base_one_cell_956/D
+ sky130_rom_krom_rom_base_one_cell_956/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_945 wl_0_2 sky130_rom_krom_rom_base_one_cell_945/D
+ sky130_rom_krom_rom_base_one_cell_945/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_934 wl_0_2 sky130_rom_krom_rom_base_one_cell_934/D
+ sky130_rom_krom_rom_base_one_cell_934/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_923 wl_0_2 sky130_rom_krom_rom_base_one_cell_923/D
+ sky130_rom_krom_rom_base_one_cell_923/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_912 wl_0_2 sky130_rom_krom_rom_base_one_cell_912/D
+ sky130_rom_krom_rom_base_one_cell_912/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_901 wl_0_2 sky130_rom_krom_rom_base_one_cell_901/D
+ sky130_rom_krom_rom_base_one_cell_901/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_989 wl_0_2 sky130_rom_krom_rom_base_one_cell_989/D
+ sky130_rom_krom_rom_base_one_cell_989/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_978 wl_0_2 sky130_rom_krom_rom_base_one_cell_978/D
+ bl_0_31 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_967 wl_0_2 sky130_rom_krom_rom_base_one_cell_967/D
+ bl_0_46 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_208 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_363/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_219 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_497/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1076 wl_0_1 sky130_rom_krom_rom_base_one_cell_692/S
+ bl_0_101 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1065 wl_0_1 sky130_rom_krom_rom_base_one_cell_812/S
+ bl_0_117 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1054 wl_0_1 sky130_rom_krom_rom_base_one_cell_801/S
+ sky130_rom_krom_rom_base_one_cell_1177/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1043 wl_0_1 sky130_rom_krom_rom_base_one_cell_309/S
+ sky130_rom_krom_rom_base_one_cell_1169/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1032 wl_0_1 sky130_rom_krom_rom_base_one_cell_782/S
+ sky130_rom_krom_rom_base_one_cell_1157/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1021 wl_0_1 sky130_rom_krom_rom_base_one_cell_892/S
+ sky130_rom_krom_rom_base_one_cell_1146/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1010 wl_0_1 sky130_rom_krom_rom_base_one_cell_644/S
+ bl_0_218 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_240 wl_0_6 sky130_rom_krom_rom_base_one_cell_731/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_251 wl_0_6 sky130_rom_krom_rom_base_one_cell_620/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_262 wl_0_5 sky130_rom_krom_rom_base_one_cell_749/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_273 wl_0_5 sky130_rom_krom_rom_base_one_cell_638/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_284 wl_0_5 sky130_rom_krom_rom_base_one_cell_649/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_295 wl_0_5 sky130_rom_krom_rom_base_one_cell_775/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1087 wl_0_1 sky130_rom_krom_rom_base_one_cell_950/S
+ sky130_rom_krom_rom_base_one_cell_1210/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1098 wl_0_1 sky130_rom_krom_rom_base_one_cell_965/S
+ bl_0_49 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_30 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_30/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_41 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_41/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_52 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_52/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_63 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_63/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_74 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_74/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_85 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_85/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_96 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_96/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_797 wl_0_3 sky130_rom_krom_rom_base_one_cell_797/D
+ sky130_rom_krom_rom_base_one_cell_914/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_786 wl_0_3 sky130_rom_krom_rom_base_one_cell_786/D
+ sky130_rom_krom_rom_base_one_cell_903/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_775 wl_0_3 sky130_rom_krom_rom_base_one_cell_775/D
+ sky130_rom_krom_rom_base_one_cell_775/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_764 wl_0_3 sky130_rom_krom_rom_base_one_cell_764/D
+ sky130_rom_krom_rom_base_one_cell_885/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_753 wl_0_3 sky130_rom_krom_rom_base_one_cell_753/D
+ sky130_rom_krom_rom_base_one_cell_753/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_742 wl_0_3 sky130_rom_krom_rom_base_one_cell_742/D
+ sky130_rom_krom_rom_base_one_cell_992/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_731 wl_0_4 sky130_rom_krom_rom_base_one_cell_731/D
+ bl_0_21 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_720 wl_0_4 sky130_rom_krom_rom_base_one_cell_720/D
+ sky130_rom_krom_rom_base_one_cell_720/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1053 wl_0_0 bl_0_1 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1042 wl_0_0 bl_0_27 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1031 wl_0_0 bl_0_46 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1020 wl_0_0 bl_0_70 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_550 wl_0_5 sky130_rom_krom_rom_base_one_cell_550/D
+ sky130_rom_krom_rom_base_one_cell_794/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_561 wl_0_5 sky130_rom_krom_rom_base_one_cell_561/D
+ sky130_rom_krom_rom_base_one_cell_561/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_572 wl_0_5 sky130_rom_krom_rom_base_one_cell_572/D
+ sky130_rom_krom_rom_base_one_cell_689/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_594 wl_0_5 sky130_rom_krom_rom_base_one_cell_594/D
+ sky130_rom_krom_rom_base_one_cell_834/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_583 wl_0_5 sky130_rom_krom_rom_base_one_cell_583/D
+ sky130_rom_krom_rom_base_one_cell_941/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_839 wl_0_1 sky130_rom_krom_rom_base_one_cell_907/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_828 wl_0_1 bl_0_196 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_817 wl_0_1 bl_0_222 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_806 wl_0_1 sky130_rom_krom_rom_base_one_cell_868/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_380 wl_0_7 sky130_rom_krom_rom_base_one_cell_380/D
+ sky130_rom_krom_rom_base_one_cell_509/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_391 wl_0_6 sky130_rom_krom_rom_base_one_cell_3/S
+ sky130_rom_krom_rom_base_one_cell_513/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_669 wl_0_3 sky130_rom_krom_rom_base_one_cell_989/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_658 wl_0_3 sky130_rom_krom_rom_base_one_cell_503/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_647 wl_0_3 sky130_rom_krom_rom_base_one_cell_720/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_636 wl_0_3 sky130_rom_krom_rom_base_one_cell_958/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_625 wl_0_3 sky130_rom_krom_rom_base_one_cell_703/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_614 wl_0_3 sky130_rom_krom_rom_base_one_cell_933/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_603 wl_0_3 sky130_rom_krom_rom_base_zero_cell_59/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1203 wl_0_0 sky130_rom_krom_rom_base_one_cell_1203/D
+ bl_0_92 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1247 wl_0_0 sky130_rom_krom_rom_base_one_cell_860/S
+ bl_0_3 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1236 wl_0_0 sky130_rom_krom_rom_base_one_cell_980/S
+ bl_0_23 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1225 wl_0_0 sky130_rom_krom_rom_base_one_cell_720/S
+ bl_0_48 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1214 wl_0_0 sky130_rom_krom_rom_base_one_cell_480/S
+ bl_0_67 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_411 wl_0_4 sky130_rom_krom_rom_base_one_cell_24/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_400 wl_0_4 sky130_rom_krom_rom_base_one_cell_744/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_499 wl_0_4 sky130_rom_krom_rom_base_zero_cell_85/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_488 wl_0_4 sky130_rom_krom_rom_base_one_cell_941/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_477 wl_0_4 sky130_rom_krom_rom_base_one_cell_813/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_466 wl_0_4 sky130_rom_krom_rom_base_one_cell_923/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_455 wl_0_4 sky130_rom_krom_rom_base_one_cell_441/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_444 wl_0_4 sky130_rom_krom_rom_base_one_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_433 wl_0_4 sky130_rom_krom_rom_base_one_cell_66/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_422 wl_0_4 sky130_rom_krom_rom_base_one_cell_764/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_979 wl_0_2 sky130_rom_krom_rom_base_one_cell_979/D
+ sky130_rom_krom_rom_base_one_cell_979/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_968 wl_0_2 sky130_rom_krom_rom_base_one_cell_968/D
+ bl_0_44 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_957 wl_0_2 sky130_rom_krom_rom_base_one_cell_957/D
+ sky130_rom_krom_rom_base_one_cell_957/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_946 wl_0_2 sky130_rom_krom_rom_base_one_cell_946/D
+ sky130_rom_krom_rom_base_one_cell_946/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_935 wl_0_2 sky130_rom_krom_rom_base_one_cell_935/D
+ sky130_rom_krom_rom_base_one_cell_935/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_924 wl_0_2 sky130_rom_krom_rom_base_one_cell_924/D
+ sky130_rom_krom_rom_base_one_cell_924/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_913 wl_0_2 sky130_rom_krom_rom_base_one_cell_913/D
+ sky130_rom_krom_rom_base_one_cell_913/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_902 wl_0_2 sky130_rom_krom_rom_base_one_cell_902/D
+ sky130_rom_krom_rom_base_one_cell_902/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_209 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_364/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_230 wl_0_6 sky130_rom_krom_rom_base_one_cell_840/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_241 wl_0_6 sky130_rom_krom_rom_base_one_cell_611/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_252 wl_0_6 sky130_rom_krom_rom_base_one_cell_621/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_263 wl_0_5 sky130_rom_krom_rom_base_zero_cell_6/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1088 wl_0_1 sky130_rom_krom_rom_base_one_cell_953/S
+ bl_0_71 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1099 wl_0_1 sky130_rom_krom_rom_base_one_cell_969/S
+ bl_0_43 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1077 wl_0_1 sky130_rom_krom_rom_base_one_cell_935/S
+ bl_0_100 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1066 wl_0_1 sky130_rom_krom_rom_base_one_cell_687/S
+ sky130_rom_krom_rom_base_one_cell_1189/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1055 wl_0_1 sky130_rom_krom_rom_base_one_cell_918/S
+ sky130_rom_krom_rom_base_one_cell_1179/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1044 wl_0_1 sky130_rom_krom_rom_base_one_cell_793/S
+ sky130_rom_krom_rom_base_one_cell_1170/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1033 wl_0_1 sky130_rom_krom_rom_base_one_cell_903/S
+ bl_0_177 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1022 wl_0_1 sky130_rom_krom_rom_base_one_cell_893/S
+ sky130_rom_krom_rom_base_one_cell_1147/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1011 wl_0_1 sky130_rom_krom_rom_base_one_cell_760/S
+ sky130_rom_krom_rom_base_one_cell_1137/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1000 wl_0_1 sky130_rom_krom_rom_base_one_cell_871/S
+ sky130_rom_krom_rom_base_one_cell_1127/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_20 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_20/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_31 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_31/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_274 wl_0_5 sky130_rom_krom_rom_base_one_cell_880/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_285 wl_0_5 sky130_rom_krom_rom_base_one_cell_765/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_296 wl_0_5 sky130_rom_krom_rom_base_one_cell_66/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_42 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_42/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_53 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_53/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_64 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_64/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_75 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_75/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_86 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_86/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_97 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_97/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_798 wl_0_3 sky130_rom_krom_rom_base_one_cell_798/D
+ sky130_rom_krom_rom_base_one_cell_916/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_787 wl_0_3 sky130_rom_krom_rom_base_one_cell_787/D
+ sky130_rom_krom_rom_base_one_cell_787/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_776 wl_0_3 sky130_rom_krom_rom_base_one_cell_776/D
+ sky130_rom_krom_rom_base_one_cell_898/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_765 wl_0_3 sky130_rom_krom_rom_base_one_cell_765/D
+ sky130_rom_krom_rom_base_one_cell_886/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_754 wl_0_3 sky130_rom_krom_rom_base_one_cell_754/D
+ sky130_rom_krom_rom_base_one_cell_873/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_743 wl_0_3 sky130_rom_krom_rom_base_one_cell_743/D
+ sky130_rom_krom_rom_base_one_cell_743/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_732 wl_0_4 sky130_rom_krom_rom_base_one_cell_732/D
+ sky130_rom_krom_rom_base_one_cell_981/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_721 wl_0_4 sky130_rom_krom_rom_base_one_cell_721/D
+ sky130_rom_krom_rom_base_one_cell_842/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_710 wl_0_4 sky130_rom_krom_rom_base_one_cell_710/D
+ sky130_rom_krom_rom_base_one_cell_958/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1010 wl_0_0 bl_0_87 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1054 wl_0_0 bl_0_0 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1043 wl_0_0 bl_0_24 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1032 wl_0_0 bl_0_45 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1021 wl_0_0 bl_0_68 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_540 wl_0_5 sky130_rom_krom_rom_base_one_cell_540/D
+ sky130_rom_krom_rom_base_one_cell_661/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_551 wl_0_5 sky130_rom_krom_rom_base_one_cell_551/D
+ sky130_rom_krom_rom_base_one_cell_674/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_562 wl_0_5 sky130_rom_krom_rom_base_zero_cell_56/S
+ sky130_rom_krom_rom_base_one_cell_924/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_573 wl_0_5 sky130_rom_krom_rom_base_one_cell_573/D
+ sky130_rom_krom_rom_base_one_cell_573/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_595 wl_0_5 sky130_rom_krom_rom_base_one_cell_595/D
+ sky130_rom_krom_rom_base_one_cell_710/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_584 wl_0_5 sky130_rom_krom_rom_base_one_cell_584/D
+ sky130_rom_krom_rom_base_one_cell_584/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_370 wl_0_7 sky130_rom_krom_rom_base_one_cell_370/D
+ sky130_rom_krom_rom_base_one_cell_845/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_381 wl_0_7 sky130_rom_krom_rom_base_one_cell_381/D
+ sky130_rom_krom_rom_base_one_cell_988/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_829 wl_0_1 sky130_rom_krom_rom_base_one_cell_896/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_818 wl_0_1 bl_0_219 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_807 wl_0_1 bl_0_241 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_392 wl_0_6 sky130_rom_krom_rom_base_one_cell_4/S
+ sky130_rom_krom_rom_base_one_cell_514/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_604 wl_0_3 sky130_rom_krom_rom_base_one_cell_928/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_659 wl_0_3 sky130_rom_krom_rom_base_one_cell_980/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_648 wl_0_3 sky130_rom_krom_rom_base_one_cell_970/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_637 wl_0_3 sky130_rom_krom_rom_base_zero_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_626 wl_0_3 sky130_rom_krom_rom_base_one_cell_704/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_615 wl_0_3 sky130_rom_krom_rom_base_one_cell_692/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1204 wl_0_0 sky130_rom_krom_rom_base_one_cell_821/S
+ bl_0_91 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1248 wl_0_0 sky130_rom_krom_rom_base_one_cell_861/S
+ bl_0_2 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1237 wl_0_0 sky130_rom_krom_rom_base_one_cell_1237/D
+ bl_0_20 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1226 wl_0_0 sky130_rom_krom_rom_base_one_cell_1226/D
+ bl_0_42 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1215 wl_0_0 sky130_rom_krom_rom_base_one_cell_956/S
+ bl_0_66 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_445 wl_0_4 sky130_rom_krom_rom_base_one_cell_791/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_434 wl_0_4 sky130_rom_krom_rom_base_one_cell_781/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_423 wl_0_4 sky130_rom_krom_rom_base_one_cell_765/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_412 wl_0_4 sky130_rom_krom_rom_base_one_cell_879/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_401 wl_0_4 sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_489 wl_0_4 sky130_rom_krom_rom_base_one_cell_584/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_478 wl_0_4 sky130_rom_krom_rom_base_one_cell_457/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_467 wl_0_4 sky130_rom_krom_rom_base_one_cell_924/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_456 wl_0_4 sky130_rom_krom_rom_base_one_cell_798/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_990 wl_0_0 bl_0_129 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_969 wl_0_2 sky130_rom_krom_rom_base_one_cell_969/D
+ sky130_rom_krom_rom_base_one_cell_969/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_958 wl_0_2 sky130_rom_krom_rom_base_one_cell_958/D
+ sky130_rom_krom_rom_base_one_cell_958/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_947 wl_0_2 sky130_rom_krom_rom_base_one_cell_947/D
+ sky130_rom_krom_rom_base_one_cell_947/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_936 wl_0_2 sky130_rom_krom_rom_base_one_cell_936/D
+ sky130_rom_krom_rom_base_one_cell_936/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_925 wl_0_2 sky130_rom_krom_rom_base_one_cell_925/D
+ sky130_rom_krom_rom_base_one_cell_925/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_914 wl_0_2 sky130_rom_krom_rom_base_one_cell_914/D
+ bl_0_150 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_903 wl_0_2 sky130_rom_krom_rom_base_one_cell_903/D
+ sky130_rom_krom_rom_base_one_cell_903/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1001 wl_0_1 sky130_rom_krom_rom_base_one_cell_753/S
+ bl_0_237 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_220 wl_0_6 sky130_rom_krom_rom_base_one_cell_956/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_231 wl_0_6 sky130_rom_krom_rom_base_one_cell_602/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_242 wl_0_6 sky130_rom_krom_rom_base_one_cell_612/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_253 wl_0_6 sky130_rom_krom_rom_base_one_cell_622/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_264 wl_0_5 sky130_rom_krom_rom_base_one_cell_751/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_275 wl_0_5 sky130_rom_krom_rom_base_one_cell_639/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_286 wl_0_5 sky130_rom_krom_rom_base_one_cell_766/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_297 wl_0_5 sky130_rom_krom_rom_base_one_cell_657/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1089 wl_0_1 sky130_rom_krom_rom_base_one_cell_954/S
+ bl_0_70 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1078 wl_0_1 sky130_rom_krom_rom_base_one_cell_936/S
+ bl_0_99 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1067 wl_0_1 sky130_rom_krom_rom_base_one_cell_929/S
+ sky130_rom_krom_rom_base_one_cell_1190/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1056 wl_0_1 sky130_rom_krom_rom_base_one_cell_920/S
+ bl_0_135 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1045 wl_0_1 sky130_rom_krom_rom_base_one_cell_673/S
+ bl_0_156 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1034 wl_0_1 sky130_rom_krom_rom_base_one_cell_663/S
+ sky130_rom_krom_rom_base_one_cell_1161/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1023 wl_0_1 sky130_rom_krom_rom_base_one_cell_894/S
+ sky130_rom_krom_rom_base_one_cell_1148/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1012 wl_0_1 sky130_rom_krom_rom_base_one_cell_761/S
+ bl_0_215 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_10 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_10/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_21 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_21/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_32 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_32/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_43 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_43/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_54 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_54/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_65 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_65/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_76 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_76/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_87 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_87/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_98 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_98/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_711 wl_0_4 sky130_rom_krom_rom_base_one_cell_711/D
+ sky130_rom_krom_rom_base_one_cell_711/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_700 wl_0_4 sky130_rom_krom_rom_base_one_cell_700/D
+ sky130_rom_krom_rom_base_one_cell_823/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_799 wl_0_3 sky130_rom_krom_rom_base_one_cell_799/D
+ sky130_rom_krom_rom_base_one_cell_799/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_788 wl_0_3 sky130_rom_krom_rom_base_one_cell_788/D
+ sky130_rom_krom_rom_base_one_cell_906/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_777 wl_0_3 sky130_rom_krom_rom_base_one_cell_66/S
+ sky130_rom_krom_rom_base_one_cell_777/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_766 wl_0_3 sky130_rom_krom_rom_base_one_cell_766/D
+ sky130_rom_krom_rom_base_one_cell_766/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_755 wl_0_3 sky130_rom_krom_rom_base_one_cell_755/D
+ sky130_rom_krom_rom_base_one_cell_875/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_744 wl_0_3 sky130_rom_krom_rom_base_one_cell_744/D
+ sky130_rom_krom_rom_base_one_cell_864/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_733 wl_0_4 sky130_rom_krom_rom_base_one_cell_733/D
+ sky130_rom_krom_rom_base_one_cell_855/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_722 wl_0_4 sky130_rom_krom_rom_base_one_cell_722/D
+ sky130_rom_krom_rom_base_one_cell_843/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1000 wl_0_0 bl_0_109 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1011 wl_0_0 bl_0_84 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1044 wl_0_0 bl_0_22 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1033 wl_0_0 bl_0_44 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1022 wl_0_0 bl_0_65 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_530 wl_0_5 sky130_rom_krom_rom_base_one_cell_530/D
+ bl_0_208 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_541 wl_0_5 sky130_rom_krom_rom_base_one_cell_541/D
+ sky130_rom_krom_rom_base_one_cell_785/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_552 wl_0_5 sky130_rom_krom_rom_base_one_cell_552/D
+ sky130_rom_krom_rom_base_one_cell_797/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_563 wl_0_5 sky130_rom_krom_rom_base_one_cell_563/D
+ sky130_rom_krom_rom_base_one_cell_563/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_574 wl_0_5 sky130_rom_krom_rom_base_one_cell_574/D
+ sky130_rom_krom_rom_base_one_cell_932/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_596 wl_0_5 sky130_rom_krom_rom_base_one_cell_596/D
+ sky130_rom_krom_rom_base_one_cell_712/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_585 wl_0_5 sky130_rom_krom_rom_base_one_cell_585/D
+ sky130_rom_krom_rom_base_one_cell_699/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_360 wl_0_7 sky130_rom_krom_rom_base_one_cell_360/D
+ sky130_rom_krom_rom_base_one_cell_481/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_371 wl_0_7 sky130_rom_krom_rom_base_one_cell_371/D
+ sky130_rom_krom_rom_base_one_cell_498/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_382 wl_0_7 sky130_rom_krom_rom_base_one_cell_382/D
+ sky130_rom_krom_rom_base_one_cell_989/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_393 wl_0_6 sky130_rom_krom_rom_base_one_cell_393/D
+ sky130_rom_krom_rom_base_one_cell_747/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_819 wl_0_1 sky130_rom_krom_rom_base_one_cell_645/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_808 wl_0_1 bl_0_240 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_627 wl_0_3 sky130_rom_krom_rom_base_one_cell_949/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_616 wl_0_3 sky130_rom_krom_rom_base_one_cell_935/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_605 wl_0_3 sky130_rom_krom_rom_base_one_cell_684/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_190 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_359/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_649 wl_0_3 sky130_rom_krom_rom_base_one_cell_971/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_638 wl_0_3 sky130_rom_krom_rom_base_one_cell_711/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1205 wl_0_0 sky130_rom_krom_rom_base_one_cell_942/S
+ bl_0_89 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1238 wl_0_0 sky130_rom_krom_rom_base_one_cell_982/S
+ bl_0_19 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1227 wl_0_0 sky130_rom_krom_rom_base_one_cell_494/S
+ bl_0_39 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1216 wl_0_0 sky130_rom_krom_rom_base_one_cell_958/S
+ bl_0_64 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_479 wl_0_4 sky130_rom_krom_rom_base_one_cell_573/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_468 wl_0_4 sky130_rom_krom_rom_base_zero_cell_57/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_457 wl_0_4 sky130_rom_krom_rom_base_one_cell_917/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_446 wl_0_4 sky130_rom_krom_rom_base_one_cell_437/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_435 wl_0_4 sky130_rom_krom_rom_base_one_cell_423/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_424 wl_0_4 sky130_rom_krom_rom_base_one_cell_766/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_413 wl_0_4 sky130_rom_krom_rom_base_one_cell_880/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_402 wl_0_4 sky130_rom_krom_rom_base_one_cell_746/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_904 wl_0_2 sky130_rom_krom_rom_base_one_cell_904/D
+ bl_0_173 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_980 wl_0_0 bl_0_150 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_991 wl_0_0 bl_0_128 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_959 wl_0_2 sky130_rom_krom_rom_base_one_cell_959/D
+ sky130_rom_krom_rom_base_one_cell_959/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_948 wl_0_2 sky130_rom_krom_rom_base_one_cell_948/D
+ sky130_rom_krom_rom_base_one_cell_948/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_937 wl_0_2 sky130_rom_krom_rom_base_one_cell_937/D
+ bl_0_97 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_926 wl_0_2 sky130_rom_krom_rom_base_zero_cell_59/S
+ bl_0_124 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_915 wl_0_2 sky130_rom_krom_rom_base_one_cell_915/D
+ bl_0_148 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1035 wl_0_1 sky130_rom_krom_rom_base_one_cell_543/S
+ bl_0_174 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1024 wl_0_1 sky130_rom_krom_rom_base_one_cell_895/S
+ sky130_rom_krom_rom_base_one_cell_1149/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1013 wl_0_1 sky130_rom_krom_rom_base_one_cell_646/S
+ sky130_rom_krom_rom_base_one_cell_1138/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1002 wl_0_1 sky130_rom_krom_rom_base_one_cell_872/S
+ bl_0_236 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_210 wl_0_6 sky130_rom_krom_rom_base_one_cell_826/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_221 wl_0_6 sky130_rom_krom_rom_base_one_cell_957/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_232 wl_0_6 sky130_rom_krom_rom_base_one_cell_722/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_243 wl_0_6 sky130_rom_krom_rom_base_one_cell_615/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_254 wl_0_6 sky130_rom_krom_rom_base_one_cell_623/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_265 wl_0_5 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_276 wl_0_5 sky130_rom_krom_rom_base_one_cell_273/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_287 wl_0_5 sky130_rom_krom_rom_base_one_cell_650/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_298 wl_0_5 sky130_rom_krom_rom_base_one_cell_660/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1079 wl_0_1 sky130_rom_krom_rom_base_one_cell_939/S
+ sky130_rom_krom_rom_base_one_cell_1200/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1068 wl_0_1 sky130_rom_krom_rom_base_one_cell_930/S
+ sky130_rom_krom_rom_base_one_cell_1191/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1057 wl_0_1 sky130_rom_krom_rom_base_one_cell_922/S
+ bl_0_133 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1046 wl_0_1 sky130_rom_krom_rom_base_one_cell_794/S
+ sky130_rom_krom_rom_base_one_cell_1171/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_11 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_11/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_22 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_22/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_33 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_33/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_44 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_44/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_55 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_55/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_66 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_66/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_77 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_77/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_88 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_88/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_99 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_99/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_745 wl_0_3 sky130_rom_krom_rom_base_one_cell_745/D
+ sky130_rom_krom_rom_base_one_cell_993/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_734 wl_0_4 sky130_rom_krom_rom_base_one_cell_734/D
+ sky130_rom_krom_rom_base_one_cell_984/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_723 wl_0_4 sky130_rom_krom_rom_base_one_cell_723/D
+ sky130_rom_krom_rom_base_one_cell_970/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_712 wl_0_4 sky130_rom_krom_rom_base_one_cell_712/D
+ sky130_rom_krom_rom_base_one_cell_959/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_701 wl_0_4 sky130_rom_krom_rom_base_one_cell_701/D
+ sky130_rom_krom_rom_base_one_cell_824/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_789 wl_0_3 sky130_rom_krom_rom_base_one_cell_789/D
+ sky130_rom_krom_rom_base_one_cell_907/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_778 wl_0_3 sky130_rom_krom_rom_base_one_cell_778/D
+ sky130_rom_krom_rom_base_one_cell_778/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_767 wl_0_3 sky130_rom_krom_rom_base_one_cell_767/D
+ sky130_rom_krom_rom_base_one_cell_887/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_756 wl_0_3 sky130_rom_krom_rom_base_one_cell_756/D
+ sky130_rom_krom_rom_base_one_cell_756/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1001 wl_0_0 bl_0_106 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1012 wl_0_0 bl_0_82 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1045 wl_0_0 bl_0_21 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1034 wl_0_0 bl_0_43 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1023 wl_0_0 bl_0_62 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_520 wl_0_5 sky130_rom_krom_rom_base_zero_cell_8/S
+ sky130_rom_krom_rom_base_one_cell_753/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_531 wl_0_5 sky130_rom_krom_rom_base_one_cell_531/D
+ sky130_rom_krom_rom_base_one_cell_764/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_542 wl_0_5 sky130_rom_krom_rom_base_one_cell_542/D
+ sky130_rom_krom_rom_base_one_cell_786/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_553 wl_0_5 sky130_rom_krom_rom_base_one_cell_553/D
+ sky130_rom_krom_rom_base_one_cell_675/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_564 wl_0_5 sky130_rom_krom_rom_base_zero_cell_58/S
+ sky130_rom_krom_rom_base_one_cell_807/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_575 wl_0_5 sky130_rom_krom_rom_base_one_cell_575/D
+ sky130_rom_krom_rom_base_one_cell_691/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_597 wl_0_5 sky130_rom_krom_rom_base_zero_cell_91/S
+ sky130_rom_krom_rom_base_one_cell_713/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_586 wl_0_5 sky130_rom_krom_rom_base_zero_cell_77/S
+ sky130_rom_krom_rom_base_one_cell_700/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_809 wl_0_1 sky130_rom_krom_rom_base_one_cell_873/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_350 wl_0_7 sky130_rom_krom_rom_base_one_cell_350/D
+ sky130_rom_krom_rom_base_one_cell_590/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_361 wl_0_7 sky130_rom_krom_rom_base_one_cell_361/D
+ sky130_rom_krom_rom_base_one_cell_716/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_372 wl_0_7 sky130_rom_krom_rom_base_one_cell_372/D
+ sky130_rom_krom_rom_base_one_cell_500/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_383 wl_0_7 sky130_rom_krom_rom_base_one_cell_383/D
+ sky130_rom_krom_rom_base_one_cell_739/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_394 wl_0_6 sky130_rom_krom_rom_base_one_cell_394/D
+ sky130_rom_krom_rom_base_one_cell_629/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_639 wl_0_3 sky130_rom_krom_rom_base_one_cell_959/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_628 wl_0_3 sky130_rom_krom_rom_base_one_cell_950/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_617 wl_0_3 bl_0_98 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_606 wl_0_3 sky130_rom_krom_rom_base_one_cell_687/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_180 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_353/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_191 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_360/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1206 wl_0_0 sky130_rom_krom_rom_base_one_cell_945/S
+ bl_0_86 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1217 wl_0_0 sky130_rom_krom_rom_base_one_cell_1217/D
+ bl_0_63 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1239 wl_0_0 sky130_rom_krom_rom_base_one_cell_1239/D
+ bl_0_18 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1228 wl_0_0 sky130_rom_krom_rom_base_one_cell_974/S
+ bl_0_37 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_469 wl_0_4 sky130_rom_krom_rom_base_one_cell_563/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_458 wl_0_4 sky130_rom_krom_rom_base_one_cell_445/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_447 wl_0_4 sky130_rom_krom_rom_base_one_cell_309/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_436 wl_0_4 sky130_rom_krom_rom_base_one_cell_782/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_425 wl_0_4 sky130_rom_krom_rom_base_one_cell_52/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_414 wl_0_4 sky130_rom_krom_rom_base_one_cell_273/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_403 wl_0_4 sky130_rom_krom_rom_base_one_cell_747/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_938 wl_0_2 sky130_rom_krom_rom_base_one_cell_938/D
+ sky130_rom_krom_rom_base_one_cell_938/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_927 wl_0_2 sky130_rom_krom_rom_base_one_cell_927/D
+ sky130_rom_krom_rom_base_one_cell_927/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_916 wl_0_2 sky130_rom_krom_rom_base_one_cell_916/D
+ sky130_rom_krom_rom_base_one_cell_916/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_905 wl_0_2 sky130_rom_krom_rom_base_one_cell_905/D
+ sky130_rom_krom_rom_base_one_cell_905/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_970 wl_0_0 bl_0_170 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_981 wl_0_0 bl_0_149 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_992 wl_0_0 bl_0_127 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_949 wl_0_2 sky130_rom_krom_rom_base_one_cell_949/D
+ bl_0_79 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_200 wl_0_6 sky130_rom_krom_rom_base_one_cell_574/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_211 wl_0_6 sky130_rom_krom_rom_base_zero_cell_80/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1058 wl_0_1 sky130_rom_krom_rom_base_one_cell_924/S
+ sky130_rom_krom_rom_base_one_cell_1183/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1047 wl_0_1 sky130_rom_krom_rom_base_zero_cell_46/S
+ bl_0_153 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1036 wl_0_1 sky130_rom_krom_rom_base_one_cell_905/S
+ bl_0_172 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1025 wl_0_1 sky130_rom_krom_rom_base_one_cell_897/S
+ sky130_rom_krom_rom_base_one_cell_1151/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1014 wl_0_1 sky130_rom_krom_rom_base_one_cell_883/S
+ sky130_rom_krom_rom_base_one_cell_1139/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1003 wl_0_1 sky130_rom_krom_rom_base_one_cell_874/S
+ sky130_rom_krom_rom_base_one_cell_1129/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_222 wl_0_6 sky130_rom_krom_rom_base_zero_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_233 wl_0_6 sky130_rom_krom_rom_base_one_cell_725/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_244 wl_0_6 sky130_rom_krom_rom_base_one_cell_616/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_255 wl_0_6 sky130_rom_krom_rom_base_one_cell_624/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_266 wl_0_5 sky130_rom_krom_rom_base_zero_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_277 wl_0_5 sky130_rom_krom_rom_base_one_cell_758/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_288 wl_0_5 sky130_rom_krom_rom_base_one_cell_52/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_299 wl_0_5 sky130_rom_krom_rom_base_one_cell_781/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1069 wl_0_1 sky130_rom_krom_rom_base_one_cell_573/S
+ sky130_rom_krom_rom_base_one_cell_1193/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_12 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_5/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_23 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_23/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_34 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_34/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_45 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_45/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_56 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_56/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_67 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_67/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_78 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_78/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_89 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_89/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_779 wl_0_3 sky130_rom_krom_rom_base_one_cell_779/D
+ sky130_rom_krom_rom_base_one_cell_899/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_768 wl_0_3 sky130_rom_krom_rom_base_one_cell_52/S
+ sky130_rom_krom_rom_base_one_cell_888/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_757 wl_0_3 sky130_rom_krom_rom_base_one_cell_757/D
+ bl_0_225 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_746 wl_0_3 sky130_rom_krom_rom_base_one_cell_746/D
+ sky130_rom_krom_rom_base_one_cell_994/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_735 wl_0_4 sky130_rom_krom_rom_base_one_cell_735/D
+ sky130_rom_krom_rom_base_one_cell_856/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_724 wl_0_4 sky130_rom_krom_rom_base_one_cell_724/D
+ sky130_rom_krom_rom_base_one_cell_971/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_713 wl_0_4 sky130_rom_krom_rom_base_one_cell_713/D
+ sky130_rom_krom_rom_base_one_cell_836/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_702 wl_0_4 sky130_rom_krom_rom_base_zero_cell_78/S
+ sky130_rom_krom_rom_base_one_cell_825/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1002 wl_0_0 bl_0_104 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1046 wl_0_0 bl_0_16 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1035 wl_0_0 bl_0_41 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1024 wl_0_0 bl_0_56 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1013 wl_0_0 bl_0_80 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_510 wl_0_6 sky130_rom_krom_rom_base_one_cell_510/D
+ sky130_rom_krom_rom_base_one_cell_613/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_521 wl_0_5 sky130_rom_krom_rom_base_one_cell_521/D
+ sky130_rom_krom_rom_base_one_cell_879/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_532 wl_0_5 sky130_rom_krom_rom_base_one_cell_532/D
+ sky130_rom_krom_rom_base_one_cell_651/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_543 wl_0_5 sky130_rom_krom_rom_base_one_cell_81/S
+ sky130_rom_krom_rom_base_one_cell_543/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_554 wl_0_5 sky130_rom_krom_rom_base_one_cell_554/D
+ sky130_rom_krom_rom_base_one_cell_677/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_565 wl_0_5 sky130_rom_krom_rom_base_zero_cell_60/S
+ sky130_rom_krom_rom_base_one_cell_809/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_576 wl_0_5 sky130_rom_krom_rom_base_one_cell_576/D
+ sky130_rom_krom_rom_base_one_cell_817/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_598 wl_0_5 sky130_rom_krom_rom_base_one_cell_598/D
+ sky130_rom_krom_rom_base_one_cell_717/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_587 wl_0_5 sky130_rom_krom_rom_base_one_cell_587/D
+ sky130_rom_krom_rom_base_one_cell_701/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_0 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_0/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_340 wl_0_7 sky130_rom_krom_rom_base_one_cell_340/D
+ sky130_rom_krom_rom_base_one_cell_466/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_351 wl_0_7 sky130_rom_krom_rom_base_one_cell_351/D
+ sky130_rom_krom_rom_base_one_cell_707/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_362 wl_0_7 sky130_rom_krom_rom_base_one_cell_362/D
+ sky130_rom_krom_rom_base_one_cell_486/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_373 wl_0_7 sky130_rom_krom_rom_base_one_cell_373/D
+ sky130_rom_krom_rom_base_one_cell_501/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_384 wl_0_7 sky130_rom_krom_rom_base_one_cell_384/D
+ sky130_rom_krom_rom_base_one_cell_618/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_395 wl_0_6 sky130_rom_krom_rom_base_one_cell_395/D
+ sky130_rom_krom_rom_base_one_cell_630/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_170 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_78/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_629 wl_0_3 sky130_rom_krom_rom_base_one_cell_952/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_618 wl_0_3 sky130_rom_krom_rom_base_one_cell_937/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_607 wl_0_3 bl_0_115 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_181 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_354/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_192 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_87/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1207 wl_0_0 sky130_rom_krom_rom_base_one_cell_946/S
+ bl_0_85 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1229 wl_0_0 sky130_rom_krom_rom_base_one_cell_975/S
+ bl_0_36 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1218 wl_0_0 sky130_rom_krom_rom_base_one_cell_835/S
+ bl_0_61 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_459 wl_0_4 bl_0_141 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_448 wl_0_4 bl_0_158 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_437 wl_0_4 sky130_rom_krom_rom_base_one_cell_784/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_426 wl_0_4 sky130_rom_krom_rom_base_one_cell_770/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_415 wl_0_4 sky130_rom_krom_rom_base_one_cell_881/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_404 wl_0_4 sky130_rom_krom_rom_base_one_cell_749/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_939 wl_0_2 sky130_rom_krom_rom_base_one_cell_939/D
+ sky130_rom_krom_rom_base_one_cell_939/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_928 wl_0_2 sky130_rom_krom_rom_base_one_cell_928/D
+ sky130_rom_krom_rom_base_one_cell_928/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_917 wl_0_2 sky130_rom_krom_rom_base_one_cell_917/D
+ sky130_rom_krom_rom_base_one_cell_917/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_906 wl_0_2 sky130_rom_krom_rom_base_one_cell_906/D
+ sky130_rom_krom_rom_base_one_cell_906/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_960 wl_0_0 bl_0_191 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_971 wl_0_0 bl_0_166 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_982 wl_0_0 bl_0_148 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_993 wl_0_0 bl_0_124 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_201 wl_0_6 sky130_rom_krom_rom_base_zero_cell_69/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_212 wl_0_6 sky130_rom_krom_rom_base_one_cell_590/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_223 wl_0_6 sky130_rom_krom_rom_base_zero_cell_89/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_234 wl_0_6 sky130_rom_krom_rom_base_one_cell_845/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_245 wl_0_6 sky130_rom_krom_rom_base_one_cell_617/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1059 wl_0_1 sky130_rom_krom_rom_base_one_cell_563/S
+ bl_0_128 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1048 wl_0_1 sky130_rom_krom_rom_base_one_cell_796/S
+ bl_0_151 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1037 wl_0_1 sky130_rom_krom_rom_base_one_cell_787/S
+ bl_0_171 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1026 wl_0_1 sky130_rom_krom_rom_base_one_cell_775/S
+ bl_0_191 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1015 wl_0_1 sky130_rom_krom_rom_base_one_cell_884/S
+ bl_0_212 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1004 wl_0_1 sky130_rom_krom_rom_base_one_cell_878/S
+ bl_0_229 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_13 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_6/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_256 wl_0_5 sky130_rom_krom_rom_base_one_cell_625/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_267 wl_0_5 sky130_rom_krom_rom_base_one_cell_754/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_278 wl_0_5 sky130_rom_krom_rom_base_one_cell_34/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_289 wl_0_5 sky130_rom_krom_rom_base_one_cell_771/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_precharge_array_0 bl_0_0 bl_0_1 bl_0_3 bl_0_6 bl_0_8 bl_0_9 bl_0_10
+ bl_0_13 bl_0_15 bl_0_16 bl_0_22 bl_0_24 bl_0_26 bl_0_29 bl_0_31 bl_0_33 bl_0_34
+ bl_0_36 bl_0_38 bl_0_40 bl_0_43 bl_0_44 bl_0_46 bl_0_47 bl_0_52 bl_0_53 bl_0_54
+ bl_0_56 bl_0_58 bl_0_59 bl_0_60 bl_0_61 bl_0_62 bl_0_65 bl_0_68 bl_0_70 bl_0_71
+ bl_0_74 bl_0_77 bl_0_79 bl_0_80 bl_0_81 bl_0_83 bl_0_86 bl_0_88 bl_0_89 bl_0_90
+ bl_0_91 bl_0_95 bl_0_97 bl_0_98 bl_0_102 bl_0_104 bl_0_106 bl_0_109 bl_0_111 bl_0_113
+ bl_0_114 bl_0_116 bl_0_118 bl_0_120 bl_0_123 bl_0_124 bl_0_127 bl_0_132 bl_0_133
+ bl_0_134 bl_0_139 bl_0_141 bl_0_142 bl_0_143 bl_0_144 bl_0_145 bl_0_148 bl_0_150
+ bl_0_151 bl_0_153 bl_0_156 bl_0_157 bl_0_160 bl_0_162 bl_0_163 bl_0_165 bl_0_166
+ bl_0_167 bl_0_172 bl_0_174 bl_0_175 bl_0_177 bl_0_181 bl_0_183 bl_0_184 bl_0_185
+ bl_0_186 bl_0_190 bl_0_192 bl_0_193 bl_0_195 bl_0_196 bl_0_202 bl_0_204 bl_0_206
+ bl_0_209 bl_0_211 bl_0_213 bl_0_214 bl_0_215 bl_0_218 bl_0_220 bl_0_222 bl_0_223
+ bl_0_224 bl_0_227 bl_0_229 bl_0_232 bl_0_233 bl_0_234 bl_0_239 bl_0_241 bl_0_242
+ bl_0_243 bl_0_245 bl_0_248 bl_0_250 bl_0_251 bl_0_252 bl_0_254 precharge bl_0_197
+ bl_0_158 bl_0_188 bl_0_146 bl_0_72 bl_0_216 bl_0_179 bl_0_45 bl_0_125 bl_0_27 bl_0_107
+ bl_0_155 bl_0_20 bl_0_137 bl_0_100 bl_0_50 bl_0_63 bl_0_130 bl_0_93 bl_0_225 bl_0_207
+ bl_0_170 bl_0_237 bl_0_200 bl_0_246 bl_0_18 bl_0_230 bl_0_48 bl_0_11 bl_0_128 bl_0_41
+ bl_0_4 bl_0_121 bl_0_168 bl_0_84 bl_0_66 bl_0_198 bl_0_161 bl_0_255 bl_0_96 bl_0_228
+ bl_0_191 bl_0_126 bl_0_39 bl_0_221 bl_0_2 bl_0_119 bl_0_82 bl_0_32 bl_0_149 bl_0_112
+ bl_0_244 bl_0_75 bl_0_159 bl_0_25 bl_0_253 bl_0_226 bl_0_57 bl_0_189 bl_0_105 bl_0_7
+ bl_0_55 bl_0_87 bl_0_37 bl_0_135 bl_0_219 bl_0_182 bl_0_117 bl_0_212 bl_0_30 bl_0_147
+ bl_0_110 bl_0_73 bl_0_205 bl_0_23 bl_0_140 bl_0_187 bl_0_103 bl_0_235 bl_0_217 bl_0_180
+ bl_0_78 bl_0_210 bl_0_28 bl_0_173 bl_0_108 bl_0_240 bl_0_203 bl_0_249 bl_0_21 bl_0_138
+ bl_0_101 bl_0_51 bl_0_64 bl_0_14 bl_0_131 bl_0_178 bl_0_94 bl_0_76 bl_0_208 bl_0_171
+ bl_0_238 bl_0_154 bl_0_69 bl_0_19 bl_0_201 bl_0_247 bl_0_136 bl_0_164 bl_0_99 bl_0_231
+ bl_0_49 bl_0_194 bl_0_12 bl_0_129 bl_0_176 bl_0_92 bl_0_42 bl_0_5 bl_0_122 bl_0_85
+ bl_0_169 bl_0_35 bl_0_236 bl_0_152 bl_0_67 vdd bl_0_199 bl_0_115 bl_0_17 sky130_rom_krom_rom_precharge_array
Xsky130_rom_krom_rom_base_one_cell_24 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_24/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_35 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_35/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_46 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_46/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_57 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_57/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_68 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_68/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_79 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_79/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_790 wl_0_2 sky130_rom_krom_rom_base_one_cell_854/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_769 wl_0_3 sky130_rom_krom_rom_base_one_cell_769/D
+ sky130_rom_krom_rom_base_one_cell_889/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_758 wl_0_3 sky130_rom_krom_rom_base_one_cell_758/D
+ sky130_rom_krom_rom_base_one_cell_882/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_747 wl_0_3 sky130_rom_krom_rom_base_one_cell_747/D
+ sky130_rom_krom_rom_base_one_cell_866/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_736 wl_0_4 sky130_rom_krom_rom_base_one_cell_736/D
+ sky130_rom_krom_rom_base_one_cell_857/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_725 wl_0_4 sky130_rom_krom_rom_base_one_cell_725/D
+ sky130_rom_krom_rom_base_one_cell_972/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_714 wl_0_4 sky130_rom_krom_rom_base_one_cell_714/D
+ sky130_rom_krom_rom_base_one_cell_960/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_703 wl_0_4 sky130_rom_krom_rom_base_one_cell_703/D
+ sky130_rom_krom_rom_base_one_cell_703/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1003 wl_0_0 bl_0_101 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1047 wl_0_0 bl_0_15 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1036 wl_0_0 bl_0_40 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1025 wl_0_0 bl_0_53 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1014 wl_0_0 bl_0_79 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_500 wl_0_6 sky130_rom_krom_rom_base_one_cell_500/D
+ sky130_rom_krom_rom_base_one_cell_607/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_511 wl_0_6 sky130_rom_krom_rom_base_one_cell_511/D
+ sky130_rom_krom_rom_base_one_cell_614/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_522 wl_0_5 sky130_rom_krom_rom_base_one_cell_522/D
+ sky130_rom_krom_rom_base_one_cell_640/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_533 wl_0_5 sky130_rom_krom_rom_base_one_cell_533/D
+ sky130_rom_krom_rom_base_one_cell_770/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_544 wl_0_5 sky130_rom_krom_rom_base_one_cell_544/D
+ sky130_rom_krom_rom_base_one_cell_904/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_555 wl_0_5 sky130_rom_krom_rom_base_zero_cell_49/S
+ sky130_rom_krom_rom_base_one_cell_917/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_566 wl_0_5 sky130_rom_krom_rom_base_one_cell_566/D
+ sky130_rom_krom_rom_base_one_cell_683/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_577 wl_0_5 sky130_rom_krom_rom_base_one_cell_577/D
+ sky130_rom_krom_rom_base_one_cell_818/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_599 wl_0_5 sky130_rom_krom_rom_base_zero_cell_97/S
+ sky130_rom_krom_rom_base_one_cell_718/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_588 wl_0_5 sky130_rom_krom_rom_base_one_cell_588/D
+ sky130_rom_krom_rom_base_one_cell_703/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_1/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_330 wl_0_7 sky130_rom_krom_rom_base_one_cell_330/D
+ sky130_rom_krom_rom_base_one_cell_566/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_341 wl_0_7 sky130_rom_krom_rom_base_one_cell_341/D
+ sky130_rom_krom_rom_base_one_cell_582/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_352 wl_0_7 sky130_rom_krom_rom_base_one_cell_352/D
+ sky130_rom_krom_rom_base_one_cell_476/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_363 wl_0_7 sky130_rom_krom_rom_base_one_cell_363/D
+ sky130_rom_krom_rom_base_one_cell_840/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_374 wl_0_7 sky130_rom_krom_rom_base_one_cell_374/D
+ sky130_rom_krom_rom_base_one_cell_503/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_385 wl_0_7 sky130_rom_krom_rom_base_one_cell_385/D
+ sky130_rom_krom_rom_base_one_cell_619/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_396 wl_0_6 sky130_rom_krom_rom_base_one_cell_396/D
+ sky130_rom_krom_rom_base_one_cell_749/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_160 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_342/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_171 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_348/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_182 precharge gnd_uq0 bl_0_73 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_193 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_88/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_619 wl_0_3 sky130_rom_krom_rom_base_one_cell_939/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_608 wl_0_3 sky130_rom_krom_rom_base_one_cell_929/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1219 wl_0_0 sky130_rom_krom_rom_base_one_cell_959/S
+ bl_0_60 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1208 wl_0_0 sky130_rom_krom_rom_base_one_cell_703/S
+ bl_0_83 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_427 wl_0_4 sky130_rom_krom_rom_base_one_cell_771/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_416 wl_0_4 sky130_rom_krom_rom_base_one_cell_758/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_405 wl_0_4 sky130_rom_krom_rom_base_zero_cell_6/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_449 wl_0_4 sky130_rom_krom_rom_base_one_cell_98/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_438 wl_0_4 sky130_rom_krom_rom_base_one_cell_785/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_950 wl_0_0 bl_0_215 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_961 wl_0_0 bl_0_190 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_972 wl_0_0 bl_0_165 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_983 wl_0_0 bl_0_147 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_929 wl_0_2 sky130_rom_krom_rom_base_one_cell_929/D
+ sky130_rom_krom_rom_base_one_cell_929/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_918 wl_0_2 sky130_rom_krom_rom_base_one_cell_918/D
+ sky130_rom_krom_rom_base_one_cell_918/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_907 wl_0_2 sky130_rom_krom_rom_base_one_cell_907/D
+ sky130_rom_krom_rom_base_one_cell_907/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_0 wl_0_7 sky130_rom_krom_rom_base_one_cell_0/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_994 wl_0_0 bl_0_122 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_202 wl_0_6 sky130_rom_krom_rom_base_zero_cell_72/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_213 wl_0_6 sky130_rom_krom_rom_base_one_cell_707/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_224 wl_0_6 sky130_rom_krom_rom_base_zero_cell_91/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_235 wl_0_6 sky130_rom_krom_rom_base_one_cell_726/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_246 wl_0_6 sky130_rom_krom_rom_base_one_cell_988/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_257 wl_0_5 sky130_rom_krom_rom_base_one_cell_626/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_268 wl_0_5 sky130_rom_krom_rom_base_one_cell_635/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_279 wl_0_5 sky130_rom_krom_rom_base_one_cell_643/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1049 wl_0_1 sky130_rom_krom_rom_base_one_cell_441/S
+ bl_0_149 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1038 wl_0_1 sky130_rom_krom_rom_base_one_cell_906/S
+ bl_0_170 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1027 wl_0_1 sky130_rom_krom_rom_base_one_cell_777/S
+ sky130_rom_krom_rom_base_one_cell_1152/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1016 wl_0_1 sky130_rom_krom_rom_base_one_cell_648/S
+ bl_0_210 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1005 wl_0_1 sky130_rom_krom_rom_base_one_cell_756/S
+ sky130_rom_krom_rom_base_one_cell_1131/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_14 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_14/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_25 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_25/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_36 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_36/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_47 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_47/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_58 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_58/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_69 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_69/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_791 wl_0_2 sky130_rom_krom_rom_base_one_cell_857/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_780 wl_0_2 sky130_rom_krom_rom_base_one_cell_845/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_759 wl_0_3 sky130_rom_krom_rom_base_one_cell_759/D
+ sky130_rom_krom_rom_base_one_cell_759/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_748 wl_0_3 sky130_rom_krom_rom_base_one_cell_748/D
+ sky130_rom_krom_rom_base_one_cell_867/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_737 wl_0_4 sky130_rom_krom_rom_base_one_cell_737/D
+ sky130_rom_krom_rom_base_one_cell_737/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_726 wl_0_4 sky130_rom_krom_rom_base_one_cell_726/D
+ sky130_rom_krom_rom_base_one_cell_976/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_715 wl_0_4 sky130_rom_krom_rom_base_one_cell_715/D
+ bl_0_56 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_704 wl_0_4 sky130_rom_krom_rom_base_zero_cell_80/S
+ sky130_rom_krom_rom_base_one_cell_704/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1004 wl_0_0 bl_0_100 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1048 wl_0_0 bl_0_14 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1037 wl_0_0 bl_0_38 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1026 wl_0_0 bl_0_52 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1015 wl_0_0 bl_0_78 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_501 wl_0_6 sky130_rom_krom_rom_base_one_cell_501/D
+ sky130_rom_krom_rom_base_one_cell_609/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_512 wl_0_5 sky130_rom_krom_rom_base_one_cell_512/D
+ sky130_rom_krom_rom_base_one_cell_742/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_523 wl_0_5 sky130_rom_krom_rom_base_one_cell_523/D
+ sky130_rom_krom_rom_base_one_cell_881/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_534 wl_0_5 sky130_rom_krom_rom_base_one_cell_534/D
+ sky130_rom_krom_rom_base_one_cell_892/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_545 wl_0_5 sky130_rom_krom_rom_base_one_cell_545/D
+ sky130_rom_krom_rom_base_one_cell_789/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_556 wl_0_5 sky130_rom_krom_rom_base_one_cell_556/D
+ sky130_rom_krom_rom_base_one_cell_679/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_567 wl_0_5 sky130_rom_krom_rom_base_one_cell_567/D
+ sky130_rom_krom_rom_base_one_cell_684/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_578 wl_0_5 sky130_rom_krom_rom_base_one_cell_578/D
+ sky130_rom_krom_rom_base_one_cell_692/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_589 wl_0_5 sky130_rom_krom_rom_base_one_cell_589/D
+ sky130_rom_krom_rom_base_one_cell_705/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_90 wl_0_7 sky130_rom_krom_rom_base_zero_cell_90/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_2 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_2/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_320 wl_0_7 sky130_rom_krom_rom_base_one_cell_320/D
+ sky130_rom_krom_rom_base_one_cell_556/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_331 wl_0_7 sky130_rom_krom_rom_base_one_cell_331/D
+ sky130_rom_krom_rom_base_one_cell_569/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_342 wl_0_7 sky130_rom_krom_rom_base_one_cell_342/D
+ sky130_rom_krom_rom_base_one_cell_697/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_353 wl_0_7 sky130_rom_krom_rom_base_one_cell_353/D
+ sky130_rom_krom_rom_base_one_cell_591/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_364 wl_0_7 sky130_rom_krom_rom_base_one_cell_364/D
+ sky130_rom_krom_rom_base_one_cell_602/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_375 wl_0_7 sky130_rom_krom_rom_base_one_cell_375/D
+ sky130_rom_krom_rom_base_one_cell_504/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_386 wl_0_7 sky130_rom_krom_rom_base_one_cell_386/D
+ sky130_rom_krom_rom_base_one_cell_620/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_397 wl_0_6 sky130_rom_krom_rom_base_one_cell_397/D
+ sky130_rom_krom_rom_base_one_cell_751/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_609 wl_0_3 sky130_rom_krom_rom_base_one_cell_457/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_150 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_336/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_161 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_343/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_172 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_79/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_183 precharge gnd_uq0 bl_0_72 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_194 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_89/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1209 wl_0_0 sky130_rom_krom_rom_base_one_cell_948/S
+ bl_0_81 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_439 wl_0_4 sky130_rom_krom_rom_base_one_cell_786/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_428 wl_0_4 sky130_rom_krom_rom_base_one_cell_892/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_417 wl_0_4 sky130_rom_krom_rom_base_one_cell_760/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_406 wl_0_4 sky130_rom_krom_rom_base_one_cell_870/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_940 wl_0_0 bl_0_233 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_951 wl_0_0 bl_0_212 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_962 wl_0_0 bl_0_188 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_973 wl_0_0 bl_0_164 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_984 wl_0_0 bl_0_145 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_995 wl_0_0 bl_0_120 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_919 wl_0_2 sky130_rom_krom_rom_base_one_cell_919/D
+ bl_0_136 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_908 wl_0_2 sky130_rom_krom_rom_base_one_cell_908/D
+ sky130_rom_krom_rom_base_one_cell_908/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1 wl_0_7 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1017 wl_0_1 sky130_rom_krom_rom_base_one_cell_885/S
+ sky130_rom_krom_rom_base_one_cell_1141/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1006 wl_0_1 sky130_rom_krom_rom_base_one_cell_273/S
+ sky130_rom_krom_rom_base_one_cell_1132/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_203 wl_0_6 sky130_rom_krom_rom_base_zero_cell_73/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_214 wl_0_6 sky130_rom_krom_rom_base_zero_cell_82/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_225 wl_0_6 sky130_rom_krom_rom_base_zero_cell_93/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_236 wl_0_6 sky130_rom_krom_rom_base_one_cell_606/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_247 wl_0_6 sky130_rom_krom_rom_base_one_cell_989/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_258 wl_0_5 sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_269 wl_0_5 sky130_rom_krom_rom_base_one_cell_755/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1039 wl_0_1 sky130_rom_krom_rom_base_one_cell_910/S
+ bl_0_164 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1028 wl_0_1 sky130_rom_krom_rom_base_one_cell_778/S
+ bl_0_188 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_15 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_15/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_26 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_26/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_37 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_37/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_48 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_48/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_59 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_59/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_727 wl_0_4 sky130_rom_krom_rom_base_one_cell_727/D
+ sky130_rom_krom_rom_base_one_cell_846/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_716 wl_0_4 sky130_rom_krom_rom_base_one_cell_716/D
+ sky130_rom_krom_rom_base_one_cell_962/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_705 wl_0_4 sky130_rom_krom_rom_base_one_cell_705/D
+ sky130_rom_krom_rom_base_one_cell_828/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_792 wl_0_2 sky130_rom_krom_rom_base_one_cell_737/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_781 wl_0_2 sky130_rom_krom_rom_base_one_cell_847/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_770 wl_0_2 sky130_rom_krom_rom_base_one_cell_711/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_749 wl_0_3 sky130_rom_krom_rom_base_one_cell_749/D
+ sky130_rom_krom_rom_base_one_cell_868/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_738 wl_0_4 sky130_rom_krom_rom_base_one_cell_738/D
+ bl_0_10 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1005 wl_0_0 bl_0_99 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1049 wl_0_0 bl_0_12 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1038 wl_0_0 bl_0_34 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1027 wl_0_0 bl_0_51 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1016 wl_0_0 bl_0_75 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_502 wl_0_6 sky130_rom_krom_rom_base_one_cell_502/D
+ sky130_rom_krom_rom_base_one_cell_730/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_513 wl_0_5 sky130_rom_krom_rom_base_one_cell_513/D
+ sky130_rom_krom_rom_base_one_cell_744/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_524 wl_0_5 sky130_rom_krom_rom_base_one_cell_524/D
+ sky130_rom_krom_rom_base_one_cell_642/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_535 wl_0_5 sky130_rom_krom_rom_base_one_cell_535/D
+ sky130_rom_krom_rom_base_one_cell_773/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_546 wl_0_5 sky130_rom_krom_rom_base_one_cell_546/D
+ sky130_rom_krom_rom_base_one_cell_791/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_557 wl_0_5 sky130_rom_krom_rom_base_zero_cell_51/S
+ sky130_rom_krom_rom_base_one_cell_801/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_568 wl_0_5 sky130_rom_krom_rom_base_zero_cell_62/S
+ sky130_rom_krom_rom_base_one_cell_685/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_579 wl_0_5 sky130_rom_krom_rom_base_zero_cell_72/S
+ sky130_rom_krom_rom_base_one_cell_694/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_80 wl_0_7 sky130_rom_krom_rom_base_zero_cell_80/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_91 wl_0_7 sky130_rom_krom_rom_base_zero_cell_91/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_3 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_3/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_310 wl_0_7 sky130_rom_krom_rom_base_one_cell_99/S
+ sky130_rom_krom_rom_base_one_cell_673/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_321 wl_0_7 sky130_rom_krom_rom_base_one_cell_321/D
+ sky130_rom_krom_rom_base_one_cell_447/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_332 wl_0_7 sky130_rom_krom_rom_base_one_cell_332/D
+ bl_0_115 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_343 wl_0_7 sky130_rom_krom_rom_base_one_cell_343/D
+ sky130_rom_krom_rom_base_one_cell_467/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_354 wl_0_7 sky130_rom_krom_rom_base_one_cell_354/D
+ sky130_rom_krom_rom_base_one_cell_477/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_365 wl_0_7 sky130_rom_krom_rom_base_one_cell_365/D
+ sky130_rom_krom_rom_base_one_cell_490/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_376 wl_0_7 sky130_rom_krom_rom_base_one_cell_376/D
+ sky130_rom_krom_rom_base_one_cell_610/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_387 wl_0_7 sky130_rom_krom_rom_base_one_cell_387/D
+ sky130_rom_krom_rom_base_one_cell_621/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_398 wl_0_6 sky130_rom_krom_rom_base_one_cell_398/D
+ sky130_rom_krom_rom_base_one_cell_519/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_140 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_332/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_151 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_337/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_162 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_344/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_173 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_80/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_184 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_85/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_195 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_90/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_429 wl_0_4 sky130_rom_krom_rom_base_one_cell_772/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_418 wl_0_4 sky130_rom_krom_rom_base_one_cell_761/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_407 wl_0_4 sky130_rom_krom_rom_base_one_cell_751/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_909 wl_0_2 sky130_rom_krom_rom_base_one_cell_909/D
+ bl_0_166 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_2 wl_0_7 sky130_rom_krom_rom_base_one_cell_4/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_930 wl_0_0 bl_0_254 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_941 wl_0_0 bl_0_232 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_952 wl_0_0 bl_0_210 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_963 wl_0_0 bl_0_185 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_974 wl_0_0 bl_0_161 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_985 wl_0_0 bl_0_142 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_996 wl_0_0 bl_0_119 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1029 wl_0_1 sky130_rom_krom_rom_base_one_cell_899/S
+ sky130_rom_krom_rom_base_one_cell_1153/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1018 wl_0_1 sky130_rom_krom_rom_base_one_cell_766/S
+ sky130_rom_krom_rom_base_one_cell_1142/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1007 wl_0_1 sky130_rom_krom_rom_base_one_cell_881/S
+ sky130_rom_krom_rom_base_one_cell_1133/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_204 wl_0_6 sky130_rom_krom_rom_base_one_cell_582/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_215 wl_0_6 sky130_rom_krom_rom_base_one_cell_591/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_226 wl_0_6 sky130_rom_krom_rom_base_one_cell_716/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_237 wl_0_6 sky130_rom_krom_rom_base_one_cell_608/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_248 wl_0_6 sky130_rom_krom_rom_base_one_cell_739/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_259 wl_0_5 sky130_rom_krom_rom_base_one_cell_747/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_16 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_27 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_27/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_38 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_38/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_49 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_49/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_739 wl_0_4 sky130_rom_krom_rom_base_one_cell_739/D
+ sky130_rom_krom_rom_base_one_cell_739/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_728 wl_0_4 sky130_rom_krom_rom_base_one_cell_728/D
+ sky130_rom_krom_rom_base_one_cell_848/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_717 wl_0_4 sky130_rom_krom_rom_base_one_cell_717/D
+ sky130_rom_krom_rom_base_one_cell_963/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_706 wl_0_4 sky130_rom_krom_rom_base_one_cell_706/D
+ sky130_rom_krom_rom_base_one_cell_949/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_793 wl_0_2 bl_0_10 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_782 wl_0_2 sky130_rom_krom_rom_base_one_cell_849/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_771 wl_0_2 sky130_rom_krom_rom_base_one_cell_835/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_760 wl_0_2 sky130_rom_krom_rom_base_one_cell_703/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1006 wl_0_0 bl_0_98 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1028 wl_0_0 bl_0_50 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1017 wl_0_0 bl_0_73 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1039 wl_0_0 bl_0_33 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_503 wl_0_6 sky130_rom_krom_rom_base_one_cell_503/D
+ sky130_rom_krom_rom_base_one_cell_503/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_514 wl_0_5 sky130_rom_krom_rom_base_one_cell_514/D
+ sky130_rom_krom_rom_base_one_cell_627/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_525 wl_0_5 sky130_rom_krom_rom_base_one_cell_525/D
+ sky130_rom_krom_rom_base_one_cell_644/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_536 wl_0_5 sky130_rom_krom_rom_base_one_cell_536/D
+ sky130_rom_krom_rom_base_one_cell_655/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_547 wl_0_5 sky130_rom_krom_rom_base_one_cell_547/D
+ sky130_rom_krom_rom_base_one_cell_671/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_558 wl_0_5 sky130_rom_krom_rom_base_one_cell_558/D
+ sky130_rom_krom_rom_base_one_cell_802/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_569 wl_0_5 sky130_rom_krom_rom_base_one_cell_569/D
+ sky130_rom_krom_rom_base_one_cell_687/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_590 wl_0_3 bl_0_145 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_70 wl_0_7 sky130_rom_krom_rom_base_zero_cell_70/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_81 wl_0_7 sky130_rom_krom_rom_base_zero_cell_81/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_92 wl_0_7 sky130_rom_krom_rom_base_zero_cell_92/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_4 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_4/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_300 wl_0_7 sky130_rom_krom_rom_base_one_cell_76/S
+ sky130_rom_krom_rom_base_one_cell_784/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_311 wl_0_7 sky130_rom_krom_rom_base_one_cell_311/D
+ sky130_rom_krom_rom_base_one_cell_439/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_322 wl_0_7 sky130_rom_krom_rom_base_one_cell_322/D
+ sky130_rom_krom_rom_base_one_cell_448/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_333 wl_0_7 sky130_rom_krom_rom_base_one_cell_333/D
+ sky130_rom_krom_rom_base_one_cell_572/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_344 wl_0_7 sky130_rom_krom_rom_base_one_cell_344/D
+ sky130_rom_krom_rom_base_one_cell_468/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_355 wl_0_7 sky130_rom_krom_rom_base_one_cell_355/D
+ sky130_rom_krom_rom_base_one_cell_478/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_366 wl_0_7 sky130_rom_krom_rom_base_one_cell_366/D
+ sky130_rom_krom_rom_base_one_cell_491/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_377 wl_0_7 sky130_rom_krom_rom_base_one_cell_377/D
+ sky130_rom_krom_rom_base_one_cell_731/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_388 wl_0_7 sky130_rom_krom_rom_base_one_cell_388/D
+ sky130_rom_krom_rom_base_one_cell_622/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_399 wl_0_6 sky130_rom_krom_rom_base_one_cell_20/S
+ sky130_rom_krom_rom_base_one_cell_754/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1190 wl_0_0 sky130_rom_krom_rom_base_one_cell_1190/D
+ bl_0_113 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_130 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_58/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_141 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_64/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_152 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_70/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_163 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_345/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_174 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_349/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_185 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_355/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_196 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_91/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_419 wl_0_4 sky130_rom_krom_rom_base_one_cell_762/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_408 wl_0_4 sky130_rom_krom_rom_base_one_cell_753/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_920 wl_0_1 sky130_rom_krom_rom_base_one_cell_983/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_931 wl_0_0 bl_0_248 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_3 wl_0_7 sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_942 wl_0_0 bl_0_231 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_953 wl_0_0 bl_0_209 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_964 wl_0_0 bl_0_181 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_975 wl_0_0 bl_0_158 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_986 wl_0_0 bl_0_141 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_997 wl_0_0 bl_0_117 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_205 wl_0_6 sky130_rom_krom_rom_base_one_cell_697/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_216 wl_0_6 bl_0_73 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_227 wl_0_6 sky130_rom_krom_rom_base_zero_cell_96/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1019 wl_0_1 sky130_rom_krom_rom_base_one_cell_887/S
+ sky130_rom_krom_rom_base_one_cell_1143/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1008 wl_0_1 sky130_rom_krom_rom_base_one_cell_641/S
+ sky130_rom_krom_rom_base_one_cell_1134/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_238 wl_0_6 sky130_rom_krom_rom_base_one_cell_851/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_249 wl_0_6 sky130_rom_krom_rom_base_one_cell_618/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_17 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_17/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_28 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_28/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_39 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_39/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_783 wl_0_2 sky130_rom_krom_rom_base_one_cell_609/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_772 wl_0_2 sky130_rom_krom_rom_base_one_cell_836/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_761 wl_0_2 sky130_rom_krom_rom_base_one_cell_704/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_750 wl_0_2 sky130_rom_krom_rom_base_one_cell_573/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_729 wl_0_4 sky130_rom_krom_rom_base_one_cell_729/D
+ sky130_rom_krom_rom_base_one_cell_849/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_718 wl_0_4 sky130_rom_krom_rom_base_one_cell_718/D
+ sky130_rom_krom_rom_base_one_cell_839/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_707 wl_0_4 sky130_rom_krom_rom_base_one_cell_707/D
+ sky130_rom_krom_rom_base_one_cell_829/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_794 wl_0_2 sky130_rom_krom_rom_base_one_cell_739/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1007 wl_0_0 bl_0_97 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1029 wl_0_0 bl_0_49 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1018 wl_0_0 bl_0_72 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_504 wl_0_6 sky130_rom_krom_rom_base_one_cell_504/D
+ sky130_rom_krom_rom_base_one_cell_852/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_515 wl_0_5 sky130_rom_krom_rom_base_one_cell_515/D
+ sky130_rom_krom_rom_base_one_cell_746/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_526 wl_0_5 sky130_rom_krom_rom_base_one_cell_526/D
+ sky130_rom_krom_rom_base_one_cell_761/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_537 wl_0_5 sky130_rom_krom_rom_base_one_cell_537/D
+ sky130_rom_krom_rom_base_one_cell_656/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_548 wl_0_5 sky130_rom_krom_rom_base_one_cell_95/S
+ sky130_rom_krom_rom_base_one_cell_672/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_559 wl_0_5 sky130_rom_krom_rom_base_one_cell_559/D
+ sky130_rom_krom_rom_base_one_cell_803/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_591 wl_0_3 sky130_rom_krom_rom_base_one_cell_917/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_580 wl_0_3 sky130_rom_krom_rom_base_one_cell_911/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_60 wl_0_7 sky130_rom_krom_rom_base_zero_cell_60/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_71 wl_0_7 sky130_rom_krom_rom_base_zero_cell_71/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_82 wl_0_7 sky130_rom_krom_rom_base_zero_cell_82/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_93 wl_0_7 sky130_rom_krom_rom_base_zero_cell_93/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_5 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_301 wl_0_7 sky130_rom_krom_rom_base_one_cell_78/S
+ sky130_rom_krom_rom_base_one_cell_542/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_312 wl_0_7 sky130_rom_krom_rom_base_one_cell_312/D
+ sky130_rom_krom_rom_base_one_cell_440/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_323 wl_0_7 sky130_rom_krom_rom_base_one_cell_323/D
+ sky130_rom_krom_rom_base_one_cell_450/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_334 wl_0_7 sky130_rom_krom_rom_base_one_cell_334/D
+ sky130_rom_krom_rom_base_one_cell_459/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_345 wl_0_7 sky130_rom_krom_rom_base_one_cell_345/D
+ sky130_rom_krom_rom_base_one_cell_469/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1180 wl_0_0 sky130_rom_krom_rom_base_one_cell_921/S
+ bl_0_134 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_356 wl_0_7 sky130_rom_krom_rom_base_one_cell_356/D
+ sky130_rom_krom_rom_base_one_cell_594/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_367 wl_0_7 sky130_rom_krom_rom_base_one_cell_367/D
+ sky130_rom_krom_rom_base_one_cell_492/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_378 wl_0_7 sky130_rom_krom_rom_base_one_cell_378/D
+ sky130_rom_krom_rom_base_one_cell_611/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_389 wl_0_6 sky130_rom_krom_rom_base_one_cell_0/S
+ sky130_rom_krom_rom_base_one_cell_625/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1191 wl_0_0 sky130_rom_krom_rom_base_one_cell_1191/D
+ bl_0_112 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_890 wl_0_2 sky130_rom_krom_rom_base_one_cell_890/D
+ bl_0_200 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_120 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_53/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_131 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_59/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_142 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_65/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_153 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_338/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_164 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_74/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_175 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_81/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_186 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_86/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_197 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_92/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_409 wl_0_4 sky130_rom_krom_rom_base_one_cell_754/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_910 wl_0_1 sky130_rom_krom_rom_base_one_cell_845/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_921 wl_0_1 bl_0_16 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_932 wl_0_0 bl_0_247 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_943 wl_0_0 bl_0_230 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_954 wl_0_0 bl_0_208 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_965 wl_0_0 bl_0_177 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_4 wl_0_7 sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_976 wl_0_0 bl_0_156 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_987 wl_0_0 bl_0_136 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_998 wl_0_0 bl_0_115 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_206 wl_0_6 sky130_rom_krom_rom_base_zero_cell_75/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_217 wl_0_6 bl_0_72 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_228 wl_0_6 sky130_rom_krom_rom_base_zero_cell_97/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_239 wl_0_6 sky130_rom_krom_rom_base_one_cell_610/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1009 wl_0_1 sky130_rom_krom_rom_base_one_cell_759/S
+ sky130_rom_krom_rom_base_one_cell_1135/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_18 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_8/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_29 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_29/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_795 wl_0_2 sky130_rom_krom_rom_base_one_cell_740/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_784 wl_0_2 sky130_rom_krom_rom_base_one_cell_850/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_773 wl_0_2 bl_0_56 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_762 wl_0_2 bl_0_80 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_751 wl_0_2 sky130_rom_krom_rom_base_one_cell_459/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_740 wl_0_2 sky130_rom_krom_rom_base_one_cell_807/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_719 wl_0_4 sky130_rom_krom_rom_base_one_cell_719/D
+ sky130_rom_krom_rom_base_one_cell_965/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_708 wl_0_4 sky130_rom_krom_rom_base_one_cell_708/D
+ sky130_rom_krom_rom_base_one_cell_950/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1008 wl_0_0 bl_0_90 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1019 wl_0_0 bl_0_71 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_505 wl_0_6 sky130_rom_krom_rom_base_one_cell_505/D
+ sky130_rom_krom_rom_base_one_cell_980/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_516 wl_0_5 sky130_rom_krom_rom_base_one_cell_7/S
+ sky130_rom_krom_rom_base_one_cell_628/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_527 wl_0_5 sky130_rom_krom_rom_base_one_cell_527/D
+ sky130_rom_krom_rom_base_one_cell_647/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_538 wl_0_5 sky130_rom_krom_rom_base_one_cell_68/S
+ sky130_rom_krom_rom_base_one_cell_658/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_549 wl_0_5 sky130_rom_krom_rom_base_one_cell_97/S
+ bl_0_158 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_592 wl_0_3 sky130_rom_krom_rom_base_one_cell_445/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_581 wl_0_3 sky130_rom_krom_rom_base_one_cell_437/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_570 wl_0_3 sky130_rom_krom_rom_base_one_cell_423/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_50 wl_0_7 sky130_rom_krom_rom_base_zero_cell_50/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_61 wl_0_7 sky130_rom_krom_rom_base_zero_cell_61/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_72 wl_0_7 sky130_rom_krom_rom_base_zero_cell_72/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_83 wl_0_7 bl_0_73 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_94 wl_0_7 sky130_rom_krom_rom_base_zero_cell_94/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_6 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_6/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_302 wl_0_7 sky130_rom_krom_rom_base_one_cell_79/S
+ sky130_rom_krom_rom_base_one_cell_663/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_313 wl_0_7 sky130_rom_krom_rom_base_one_cell_313/D
+ sky130_rom_krom_rom_base_one_cell_552/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_324 wl_0_7 sky130_rom_krom_rom_base_one_cell_324/D
+ sky130_rom_krom_rom_base_one_cell_561/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_335 wl_0_7 sky130_rom_krom_rom_base_one_cell_335/D
+ sky130_rom_krom_rom_base_one_cell_574/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_346 wl_0_7 sky130_rom_krom_rom_base_one_cell_346/D
+ sky130_rom_krom_rom_base_one_cell_472/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_357 wl_0_7 sky130_rom_krom_rom_base_one_cell_357/D
+ sky130_rom_krom_rom_base_one_cell_480/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_368 wl_0_7 sky130_rom_krom_rom_base_one_cell_368/D
+ sky130_rom_krom_rom_base_one_cell_725/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1170 wl_0_0 sky130_rom_krom_rom_base_one_cell_1170/D
+ bl_0_157 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1181 wl_0_0 sky130_rom_krom_rom_base_one_cell_561/S
+ bl_0_132 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1192 wl_0_0 sky130_rom_krom_rom_base_one_cell_457/S
+ bl_0_111 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_379 wl_0_7 sky130_rom_krom_rom_base_one_cell_379/D
+ sky130_rom_krom_rom_base_one_cell_612/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_891 wl_0_2 sky130_rom_krom_rom_base_one_cell_891/D
+ sky130_rom_krom_rom_base_one_cell_891/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_880 wl_0_2 sky130_rom_krom_rom_base_one_cell_880/D
+ bl_0_227 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_110 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_317/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_121 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_323/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_132 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_328/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_143 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_333/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_154 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_71/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_165 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_75/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_176 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_350/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_187 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_356/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_198 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_93/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_900 wl_0_1 sky130_rom_krom_rom_base_one_cell_720/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_911 wl_0_1 bl_0_34 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_922 wl_0_1 bl_0_14 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_933 wl_0_0 bl_0_246 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_944 wl_0_0 bl_0_229 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_955 wl_0_0 bl_0_206 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_966 wl_0_0 bl_0_174 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_977 wl_0_0 bl_0_153 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_988 wl_0_0 bl_0_135 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_999 wl_0_0 bl_0_114 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_5 wl_0_7 sky130_rom_krom_rom_base_zero_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_207 wl_0_6 sky130_rom_krom_rom_base_zero_cell_77/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_218 wl_0_6 sky130_rom_krom_rom_base_zero_cell_85/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_229 wl_0_6 sky130_rom_krom_rom_base_one_cell_601/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_19 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_9/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_709 wl_0_4 sky130_rom_krom_rom_base_one_cell_709/D
+ sky130_rom_krom_rom_base_one_cell_832/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_796 wl_0_2 sky130_rom_krom_rom_base_one_cell_858/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_785 wl_0_2 sky130_rom_krom_rom_base_one_cell_851/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_774 wl_0_2 sky130_rom_krom_rom_base_one_cell_837/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_763 wl_0_2 sky130_rom_krom_rom_base_one_cell_829/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_752 wl_0_2 bl_0_106 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_741 wl_0_2 sky130_rom_krom_rom_base_one_cell_808/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_730 wl_0_2 sky130_rom_krom_rom_base_one_cell_445/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_1009 wl_0_0 bl_0_88 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_506 wl_0_6 sky130_rom_krom_rom_base_one_cell_506/D
+ sky130_rom_krom_rom_base_one_cell_732/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_517 wl_0_5 sky130_rom_krom_rom_base_zero_cell_5/S
+ sky130_rom_krom_rom_base_one_cell_631/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_528 wl_0_5 sky130_rom_krom_rom_base_one_cell_528/D
+ sky130_rom_krom_rom_base_one_cell_528/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_539 wl_0_5 sky130_rom_krom_rom_base_one_cell_539/D
+ sky130_rom_krom_rom_base_one_cell_659/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_593 wl_0_3 bl_0_141 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_582 wl_0_3 sky130_rom_krom_rom_base_one_cell_912/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_571 wl_0_3 bl_0_181 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_560 wl_0_3 sky130_rom_krom_rom_base_one_cell_883/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_40 wl_0_7 sky130_rom_krom_rom_base_one_cell_92/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_51 wl_0_7 sky130_rom_krom_rom_base_zero_cell_51/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_62 wl_0_7 sky130_rom_krom_rom_base_zero_cell_62/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_73 wl_0_7 sky130_rom_krom_rom_base_zero_cell_73/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_84 wl_0_7 bl_0_72 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_95 wl_0_7 sky130_rom_krom_rom_base_zero_cell_95/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_7 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_303 wl_0_7 sky130_rom_krom_rom_base_one_cell_82/S
+ sky130_rom_krom_rom_base_one_cell_544/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_314 wl_0_7 sky130_rom_krom_rom_base_one_cell_314/D
+ sky130_rom_krom_rom_base_one_cell_441/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_325 wl_0_7 sky130_rom_krom_rom_base_one_cell_325/D
+ sky130_rom_krom_rom_base_one_cell_453/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_336 wl_0_7 sky130_rom_krom_rom_base_one_cell_336/D
+ sky130_rom_krom_rom_base_one_cell_460/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_347 wl_0_7 sky130_rom_krom_rom_base_one_cell_347/D
+ sky130_rom_krom_rom_base_one_cell_945/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_358 wl_0_7 sky130_rom_krom_rom_base_one_cell_358/D
+ sky130_rom_krom_rom_base_one_cell_956/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_369 wl_0_7 sky130_rom_krom_rom_base_one_cell_369/D
+ sky130_rom_krom_rom_base_one_cell_495/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1160 wl_0_0 sky130_rom_krom_rom_base_one_cell_785/S
+ bl_0_178 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1171 wl_0_0 sky130_rom_krom_rom_base_one_cell_1171/D
+ bl_0_155 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1182 wl_0_0 sky130_rom_krom_rom_base_one_cell_923/S
+ bl_0_131 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1193 wl_0_0 sky130_rom_krom_rom_base_one_cell_1193/D
+ bl_0_110 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_390 wl_0_5 sky130_rom_krom_rom_base_one_cell_980/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_892 wl_0_2 sky130_rom_krom_rom_base_one_cell_892/D
+ sky130_rom_krom_rom_base_one_cell_892/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_881 wl_0_2 sky130_rom_krom_rom_base_one_cell_881/D
+ sky130_rom_krom_rom_base_one_cell_881/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_870 wl_0_2 sky130_rom_krom_rom_base_one_cell_870/D
+ bl_0_241 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_100 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_45/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_111 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_49/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_122 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_54/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_133 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_60/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_144 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_66/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_155 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_339/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_166 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_76/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_177 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_351/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_188 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_357/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_199 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_94/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_6 wl_0_7 sky130_rom_krom_rom_base_zero_cell_6/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_901 wl_0_1 bl_0_47 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_912 wl_0_1 bl_0_33 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_923 wl_0_1 sky130_rom_krom_rom_base_one_cell_987/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_934 wl_0_0 bl_0_245 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_945 wl_0_0 bl_0_227 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_956 wl_0_0 bl_0_203 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_967 wl_0_0 bl_0_173 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_978 wl_0_0 bl_0_152 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_989 wl_0_0 bl_0_133 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_208 wl_0_6 sky130_rom_krom_rom_base_one_cell_945/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_219 wl_0_6 sky130_rom_krom_rom_base_one_cell_594/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_731 wl_0_2 bl_0_142 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_720 wl_0_2 bl_0_158 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_797 wl_0_2 bl_0_4 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_786 wl_0_2 sky130_rom_krom_rom_base_one_cell_503/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_775 wl_0_2 sky130_rom_krom_rom_base_one_cell_838/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_764 wl_0_2 bl_0_75 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_753 wl_0_2 sky130_rom_krom_rom_base_one_cell_816/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_742 wl_0_2 sky130_rom_krom_rom_base_one_cell_810/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_507 wl_0_6 sky130_rom_krom_rom_base_one_cell_507/D
+ sky130_rom_krom_rom_base_one_cell_853/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_518 wl_0_5 sky130_rom_krom_rom_base_one_cell_518/D
+ sky130_rom_krom_rom_base_one_cell_870/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_529 wl_0_5 sky130_rom_krom_rom_base_one_cell_45/S
+ sky130_rom_krom_rom_base_one_cell_648/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_572 wl_0_3 sky130_rom_krom_rom_base_one_cell_663/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_561 wl_0_3 sky130_rom_krom_rom_base_one_cell_528/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_550 wl_0_3 sky130_rom_krom_rom_base_one_cell_878/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_594 wl_0_3 sky130_rom_krom_rom_base_one_cell_679/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_583 wl_0_3 sky130_rom_krom_rom_base_one_cell_309/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_30 wl_0_7 sky130_rom_krom_rom_base_one_cell_72/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_41 wl_0_7 sky130_rom_krom_rom_base_one_cell_94/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_52 wl_0_7 sky130_rom_krom_rom_base_zero_cell_52/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_63 wl_0_7 sky130_rom_krom_rom_base_zero_cell_63/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_74 wl_0_7 sky130_rom_krom_rom_base_zero_cell_74/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_85 wl_0_7 sky130_rom_krom_rom_base_zero_cell_85/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_96 wl_0_7 sky130_rom_krom_rom_base_zero_cell_96/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_8 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_8/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_304 wl_0_7 sky130_rom_krom_rom_base_one_cell_83/S
+ sky130_rom_krom_rom_base_one_cell_428/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_315 wl_0_7 sky130_rom_krom_rom_base_one_cell_315/D
+ sky130_rom_krom_rom_base_one_cell_553/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_326 wl_0_7 sky130_rom_krom_rom_base_one_cell_326/D
+ sky130_rom_krom_rom_base_one_cell_806/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_337 wl_0_7 sky130_rom_krom_rom_base_one_cell_337/D
+ sky130_rom_krom_rom_base_one_cell_461/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_348 wl_0_7 sky130_rom_krom_rom_base_one_cell_348/D
+ sky130_rom_krom_rom_base_one_cell_826/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_359 wl_0_7 sky130_rom_krom_rom_base_one_cell_359/D
+ sky130_rom_krom_rom_base_one_cell_957/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1150 wl_0_0 sky130_rom_krom_rom_base_one_cell_896/S
+ bl_0_193 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1161 wl_0_0 sky130_rom_krom_rom_base_one_cell_1161/D
+ bl_0_176 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1172 wl_0_0 sky130_rom_krom_rom_base_one_cell_913/S
+ bl_0_154 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1183 wl_0_0 sky130_rom_krom_rom_base_one_cell_1183/D
+ bl_0_130 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1194 wl_0_0 sky130_rom_krom_rom_base_one_cell_1194/D
+ bl_0_108 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_391 wl_0_5 sky130_rom_krom_rom_base_one_cell_731/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_380 wl_0_5 sky130_rom_krom_rom_base_one_cell_973/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_893 wl_0_2 sky130_rom_krom_rom_base_one_cell_893/D
+ sky130_rom_krom_rom_base_one_cell_893/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_882 wl_0_2 sky130_rom_krom_rom_base_one_cell_882/D
+ bl_0_222 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_871 wl_0_2 sky130_rom_krom_rom_base_one_cell_871/D
+ sky130_rom_krom_rom_base_one_cell_871/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_860 wl_0_3 sky130_rom_krom_rom_base_one_cell_860/D
+ sky130_rom_krom_rom_base_one_cell_860/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_101 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_311/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_112 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_318/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_123 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_324/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_134 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_329/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_145 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_67/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_156 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_72/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_167 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_77/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_178 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_352/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_189 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_358/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_690 wl_0_4 sky130_rom_krom_rom_base_zero_cell_69/S
+ bl_0_106 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_902 wl_0_1 bl_0_46 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_913 wl_0_1 bl_0_31 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_7 wl_0_7 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_924 wl_0_1 bl_0_10 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_935 wl_0_0 bl_0_243 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_946 wl_0_0 bl_0_225 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_957 wl_0_0 bl_0_201 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_968 wl_0_0 bl_0_172 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_979 wl_0_0 bl_0_151 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_209 wl_0_6 sky130_rom_krom_rom_base_zero_cell_78/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_765 wl_0_2 bl_0_73 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_754 wl_0_2 sky130_rom_krom_rom_base_one_cell_818/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_743 wl_0_2 sky130_rom_krom_rom_base_one_cell_684/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_732 wl_0_2 bl_0_141 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_721 wl_0_2 sky130_rom_krom_rom_base_one_cell_793/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_710 wl_0_2 sky130_rom_krom_rom_base_one_cell_785/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_798 wl_0_2 sky130_rom_krom_rom_base_one_cell_860/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_787 wl_0_2 sky130_rom_krom_rom_base_one_cell_852/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_776 wl_0_2 bl_0_51 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_508 wl_0_6 sky130_rom_krom_rom_base_one_cell_508/D
+ sky130_rom_krom_rom_base_one_cell_854/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_519 wl_0_5 sky130_rom_krom_rom_base_one_cell_519/D
+ sky130_rom_krom_rom_base_one_cell_633/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_595 wl_0_3 sky130_rom_krom_rom_base_one_cell_680/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_584 wl_0_3 bl_0_158 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_573 wl_0_3 sky130_rom_krom_rom_base_one_cell_664/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_562 wl_0_3 sky130_rom_krom_rom_base_one_cell_648/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_551 wl_0_3 sky130_rom_krom_rom_base_one_cell_879/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_540 wl_0_3 sky130_rom_krom_rom_base_one_cell_865/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_20 wl_0_7 sky130_rom_krom_rom_base_one_cell_52/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_31 wl_0_7 sky130_rom_krom_rom_base_one_cell_74/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_42 wl_0_7 sky130_rom_krom_rom_base_one_cell_95/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_53 wl_0_7 sky130_rom_krom_rom_base_zero_cell_53/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_64 wl_0_7 sky130_rom_krom_rom_base_zero_cell_64/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_75 wl_0_7 sky130_rom_krom_rom_base_zero_cell_75/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_86 wl_0_7 sky130_rom_krom_rom_base_zero_cell_86/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_97 wl_0_7 sky130_rom_krom_rom_base_zero_cell_97/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_9 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_9/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_305 wl_0_7 sky130_rom_krom_rom_base_one_cell_88/S
+ sky130_rom_krom_rom_base_one_cell_432/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_316 wl_0_7 sky130_rom_krom_rom_base_one_cell_316/D
+ sky130_rom_krom_rom_base_one_cell_443/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_327 wl_0_7 sky130_rom_krom_rom_base_one_cell_327/D
+ sky130_rom_krom_rom_base_one_cell_327/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1140 wl_0_0 sky130_rom_krom_rom_base_one_cell_528/S
+ bl_0_211 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1151 wl_0_0 sky130_rom_krom_rom_base_one_cell_1151/D
+ bl_0_192 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1162 wl_0_0 sky130_rom_krom_rom_base_one_cell_664/S
+ bl_0_175 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_338 wl_0_7 sky130_rom_krom_rom_base_one_cell_338/D
+ sky130_rom_krom_rom_base_one_cell_463/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_349 wl_0_7 sky130_rom_krom_rom_base_one_cell_349/D
+ sky130_rom_krom_rom_base_one_cell_474/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1173 wl_0_0 sky130_rom_krom_rom_base_one_cell_799/S
+ bl_0_146 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1184 wl_0_0 sky130_rom_krom_rom_base_one_cell_327/S
+ bl_0_126 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1195 wl_0_0 sky130_rom_krom_rom_base_one_cell_1195/D
+ bl_0_107 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_392 wl_0_5 sky130_rom_krom_rom_base_one_cell_732/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_381 wl_0_5 sky130_rom_krom_rom_base_one_cell_974/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_370 wl_0_5 sky130_rom_krom_rom_base_one_cell_716/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_872 wl_0_2 sky130_rom_krom_rom_base_one_cell_872/D
+ sky130_rom_krom_rom_base_one_cell_872/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_861 wl_0_3 sky130_rom_krom_rom_base_one_cell_861/D
+ sky130_rom_krom_rom_base_one_cell_861/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_850 wl_0_3 sky130_rom_krom_rom_base_one_cell_850/D
+ sky130_rom_krom_rom_base_one_cell_850/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_894 wl_0_2 sky130_rom_krom_rom_base_one_cell_894/D
+ sky130_rom_krom_rom_base_one_cell_894/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_883 wl_0_2 sky130_rom_krom_rom_base_one_cell_883/D
+ sky130_rom_krom_rom_base_one_cell_883/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_102 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_46/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_113 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_50/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_124 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_55/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_135 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_330/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_146 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_68/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_157 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_340/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_168 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_346/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_179 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_82/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_691 wl_0_4 sky130_rom_krom_rom_base_one_cell_691/D
+ sky130_rom_krom_rom_base_one_cell_816/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_680 wl_0_4 sky130_rom_krom_rom_base_one_cell_680/D
+ sky130_rom_krom_rom_base_one_cell_680/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_903 wl_0_1 bl_0_45 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_914 wl_0_1 sky130_rom_krom_rom_base_one_cell_849/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_925 wl_0_1 sky130_rom_krom_rom_base_one_cell_988/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_936 wl_0_0 bl_0_241 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_947 wl_0_0 bl_0_222 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_8 wl_0_7 sky130_rom_krom_rom_base_zero_cell_8/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_958 wl_0_0 bl_0_200 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_969 wl_0_0 bl_0_171 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_788 wl_0_2 bl_0_22 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_777 wl_0_2 sky130_rom_krom_rom_base_one_cell_720/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_766 wl_0_2 bl_0_72 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_755 wl_0_2 sky130_rom_krom_rom_base_one_cell_692/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_744 wl_0_2 sky130_rom_krom_rom_base_one_cell_811/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_733 wl_0_2 sky130_rom_krom_rom_base_one_cell_679/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_722 wl_0_2 sky130_rom_krom_rom_base_one_cell_673/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_711 wl_0_2 sky130_rom_krom_rom_base_one_cell_663/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_700 wl_0_2 bl_0_201 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_799 wl_0_2 sky130_rom_krom_rom_base_one_cell_861/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_509 wl_0_6 sky130_rom_krom_rom_base_one_cell_509/D
+ sky130_rom_krom_rom_base_one_cell_985/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_596 wl_0_3 sky130_rom_krom_rom_base_one_cell_920/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_585 wl_0_3 sky130_rom_krom_rom_base_one_cell_673/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_574 wl_0_3 sky130_rom_krom_rom_base_one_cell_543/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_563 wl_0_3 bl_0_208 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_552 wl_0_3 sky130_rom_krom_rom_base_one_cell_880/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_541 wl_0_3 sky130_rom_krom_rom_base_one_cell_995/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_530 wl_0_4 sky130_rom_krom_rom_base_one_cell_986/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_10 wl_0_7 sky130_rom_krom_rom_base_one_cell_20/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_21 wl_0_7 sky130_rom_krom_rom_base_one_cell_53/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_32 wl_0_7 sky130_rom_krom_rom_base_one_cell_77/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_43 wl_0_7 sky130_rom_krom_rom_base_one_cell_97/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_54 wl_0_7 sky130_rom_krom_rom_base_zero_cell_54/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_65 wl_0_7 sky130_rom_krom_rom_base_zero_cell_65/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_76 wl_0_7 sky130_rom_krom_rom_base_zero_cell_76/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_87 wl_0_7 sky130_rom_krom_rom_base_zero_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_98 wl_0_7 sky130_rom_krom_rom_base_zero_cell_98/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_306 wl_0_7 sky130_rom_krom_rom_base_one_cell_90/S
+ sky130_rom_krom_rom_base_one_cell_434/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_317 wl_0_7 sky130_rom_krom_rom_base_one_cell_317/D
+ sky130_rom_krom_rom_base_one_cell_444/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_328 wl_0_7 sky130_rom_krom_rom_base_one_cell_328/D
+ sky130_rom_krom_rom_base_one_cell_808/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_339 wl_0_7 sky130_rom_krom_rom_base_one_cell_339/D
+ sky130_rom_krom_rom_base_one_cell_465/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1130 wl_0_0 sky130_rom_krom_rom_base_one_cell_879/S
+ bl_0_228 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1141 wl_0_0 sky130_rom_krom_rom_base_one_cell_1141/D
+ bl_0_207 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1152 wl_0_0 sky130_rom_krom_rom_base_one_cell_1152/D
+ bl_0_189 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1163 wl_0_0 sky130_rom_krom_rom_base_one_cell_907/S
+ bl_0_169 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1174 wl_0_0 sky130_rom_krom_rom_base_one_cell_1174/D
+ bl_0_144 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1185 wl_0_0 sky130_rom_krom_rom_base_one_cell_807/S
+ bl_0_125 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1196 wl_0_0 sky130_rom_krom_rom_base_one_cell_933/S
+ bl_0_105 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_393 wl_0_5 sky130_rom_krom_rom_base_one_cell_853/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_382 wl_0_5 sky130_rom_krom_rom_base_one_cell_975/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_371 wl_0_5 sky130_rom_krom_rom_base_one_cell_837/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_360 wl_0_5 sky130_rom_krom_rom_base_one_cell_709/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_895 wl_0_2 sky130_rom_krom_rom_base_one_cell_895/D
+ sky130_rom_krom_rom_base_one_cell_895/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_884 wl_0_2 sky130_rom_krom_rom_base_one_cell_884/D
+ sky130_rom_krom_rom_base_one_cell_884/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_873 wl_0_2 sky130_rom_krom_rom_base_one_cell_873/D
+ sky130_rom_krom_rom_base_one_cell_873/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_862 wl_0_3 sky130_rom_krom_rom_base_one_cell_862/D
+ sky130_rom_krom_rom_base_one_cell_990/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_851 wl_0_3 sky130_rom_krom_rom_base_one_cell_851/D
+ sky130_rom_krom_rom_base_one_cell_851/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_840 wl_0_3 sky130_rom_krom_rom_base_one_cell_840/D
+ sky130_rom_krom_rom_base_one_cell_966/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_103 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_47/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_114 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_319/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_125 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_56/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_136 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_61/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_147 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_334/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_158 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_73/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_169 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_347/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_190 wl_0_6 sky130_rom_krom_rom_base_one_cell_808/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_692 wl_0_4 sky130_rom_krom_rom_base_one_cell_692/D
+ sky130_rom_krom_rom_base_one_cell_692/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_681 wl_0_4 sky130_rom_krom_rom_base_one_cell_681/D
+ sky130_rom_krom_rom_base_one_cell_921/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_670 wl_0_4 sky130_rom_krom_rom_base_one_cell_670/D
+ sky130_rom_krom_rom_base_one_cell_792/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_904 wl_0_1 bl_0_44 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_915 wl_0_1 sky130_rom_krom_rom_base_one_cell_851/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_926 wl_0_1 bl_0_4 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_937 wl_0_0 bl_0_240 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_948 wl_0_0 bl_0_219 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_959 wl_0_0 bl_0_196 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_9 wl_0_7 sky130_rom_krom_rom_base_zero_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_789 wl_0_2 bl_0_21 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_778 wl_0_2 bl_0_45 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_767 wl_0_2 sky130_rom_krom_rom_base_one_cell_833/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_756 wl_0_2 bl_0_98 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_745 wl_0_2 sky130_rom_krom_rom_base_one_cell_812/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_734 wl_0_2 sky130_rom_krom_rom_base_one_cell_801/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_723 wl_0_2 sky130_rom_krom_rom_base_one_cell_794/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_712 wl_0_2 sky130_rom_krom_rom_base_one_cell_664/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_701 wl_0_2 bl_0_196 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_531 wl_0_4 sky130_rom_krom_rom_base_one_cell_988/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_520 wl_0_4 sky130_rom_krom_rom_base_one_cell_979/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_597 wl_0_3 sky130_rom_krom_rom_base_one_cell_921/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_586 wl_0_3 sky130_rom_krom_rom_base_one_cell_913/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_575 wl_0_3 sky130_rom_krom_rom_base_one_cell_904/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_564 wl_0_3 sky130_rom_krom_rom_base_one_cell_891/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_553 wl_0_3 sky130_rom_krom_rom_base_one_cell_273/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_542 wl_0_3 sky130_rom_krom_rom_base_zero_cell_6/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_11 wl_0_7 sky130_rom_krom_rom_base_one_cell_24/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_22 wl_0_7 sky130_rom_krom_rom_base_one_cell_60/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_33 wl_0_7 sky130_rom_krom_rom_base_one_cell_80/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_44 wl_0_7 sky130_rom_krom_rom_base_one_cell_98/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_55 wl_0_7 sky130_rom_krom_rom_base_zero_cell_55/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_66 wl_0_7 sky130_rom_krom_rom_base_zero_cell_66/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_77 wl_0_7 sky130_rom_krom_rom_base_zero_cell_77/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_88 wl_0_7 sky130_rom_krom_rom_base_zero_cell_88/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_99 wl_0_7 sky130_rom_krom_rom_base_zero_cell_99/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_307 wl_0_7 sky130_rom_krom_rom_base_one_cell_91/S
+ sky130_rom_krom_rom_base_one_cell_435/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_318 wl_0_7 sky130_rom_krom_rom_base_one_cell_318/D
+ sky130_rom_krom_rom_base_one_cell_445/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_329 wl_0_7 sky130_rom_krom_rom_base_one_cell_329/D
+ sky130_rom_krom_rom_base_one_cell_454/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1120 wl_0_0 sky130_rom_krom_rom_base_one_cell_864/S
+ bl_0_252 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1131 wl_0_0 sky130_rom_krom_rom_base_one_cell_1131/D
+ bl_0_226 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1142 wl_0_0 sky130_rom_krom_rom_base_one_cell_1142/D
+ bl_0_205 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1153 wl_0_0 sky130_rom_krom_rom_base_one_cell_1153/D
+ bl_0_187 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1164 wl_0_0 sky130_rom_krom_rom_base_one_cell_87/S
+ bl_0_168 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1175 wl_0_0 sky130_rom_krom_rom_base_one_cell_1175/D
+ bl_0_143 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1186 wl_0_0 sky130_rom_krom_rom_base_one_cell_808/S
+ bl_0_123 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1197 wl_0_0 sky130_rom_krom_rom_base_one_cell_1197/D
+ bl_0_103 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_372 wl_0_5 sky130_rom_krom_rom_base_zero_cell_96/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_361 wl_0_5 sky130_rom_krom_rom_base_one_cell_480/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_350 wl_0_5 sky130_rom_krom_rom_base_zero_cell_78/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_394 wl_0_5 sky130_rom_krom_rom_base_one_cell_854/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_383 wl_0_5 sky130_rom_krom_rom_base_one_cell_845/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_896 wl_0_2 sky130_rom_krom_rom_base_one_cell_62/S
+ sky130_rom_krom_rom_base_one_cell_896/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_885 wl_0_2 sky130_rom_krom_rom_base_one_cell_885/D
+ sky130_rom_krom_rom_base_one_cell_885/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_874 wl_0_2 sky130_rom_krom_rom_base_one_cell_874/D
+ sky130_rom_krom_rom_base_one_cell_874/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_863 wl_0_3 sky130_rom_krom_rom_base_one_cell_863/D
+ sky130_rom_krom_rom_base_one_cell_991/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_852 wl_0_3 sky130_rom_krom_rom_base_one_cell_852/D
+ sky130_rom_krom_rom_base_one_cell_852/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_841 wl_0_3 sky130_rom_krom_rom_base_one_cell_841/D
+ sky130_rom_krom_rom_base_one_cell_967/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_830 wl_0_3 sky130_rom_krom_rom_base_zero_cell_82/S
+ sky130_rom_krom_rom_base_one_cell_951/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_104 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_312/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_115 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_320/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_126 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_57/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_137 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_62/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_148 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_335/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_159 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_341/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_180 wl_0_6 sky130_rom_krom_rom_base_one_cell_556/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_191 wl_0_6 sky130_rom_krom_rom_base_zero_cell_60/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_693 wl_0_4 sky130_rom_krom_rom_base_one_cell_693/D
+ sky130_rom_krom_rom_base_one_cell_935/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_682 wl_0_4 sky130_rom_krom_rom_base_one_cell_682/D
+ sky130_rom_krom_rom_base_one_cell_810/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_671 wl_0_4 sky130_rom_krom_rom_base_one_cell_671/D
+ sky130_rom_krom_rom_base_one_cell_911/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_660 wl_0_4 sky130_rom_krom_rom_base_one_cell_660/D
+ sky130_rom_krom_rom_base_one_cell_901/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_490 wl_0_6 sky130_rom_krom_rom_base_one_cell_490/D
+ sky130_rom_krom_rom_base_one_cell_603/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_905 wl_0_1 bl_0_41 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_916 wl_0_1 sky130_rom_krom_rom_base_one_cell_980/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_927 wl_0_1 sky130_rom_krom_rom_base_one_cell_860/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_938 wl_0_0 bl_0_237 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_949 wl_0_0 bl_0_218 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_713 wl_0_2 sky130_rom_krom_rom_base_one_cell_543/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_702 wl_0_2 sky130_rom_krom_rom_base_one_cell_775/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_779 wl_0_2 sky130_rom_krom_rom_base_one_cell_494/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_768 wl_0_2 sky130_rom_krom_rom_base_one_cell_480/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_757 wl_0_2 sky130_rom_krom_rom_base_one_cell_584/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_746 wl_0_2 sky130_rom_krom_rom_base_one_cell_687/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_735 wl_0_2 sky130_rom_krom_rom_base_one_cell_680/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_724 wl_0_2 sky130_rom_krom_rom_base_zero_cell_46/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_554 wl_0_3 sky130_rom_krom_rom_base_one_cell_881/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_543 wl_0_3 sky130_rom_krom_rom_base_one_cell_870/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_532 wl_0_4 sky130_rom_krom_rom_base_one_cell_989/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_521 wl_0_4 sky130_rom_krom_rom_base_one_cell_609/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_510 wl_0_4 sky130_rom_krom_rom_base_one_cell_964/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_598 wl_0_3 sky130_rom_krom_rom_base_one_cell_561/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_587 wl_0_3 sky130_rom_krom_rom_base_zero_cell_46/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_576 wl_0_3 sky130_rom_krom_rom_base_one_cell_905/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_565 wl_0_3 sky130_rom_krom_rom_base_one_cell_892/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_12 wl_0_7 sky130_rom_krom_rom_base_one_cell_25/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_23 wl_0_7 sky130_rom_krom_rom_base_one_cell_61/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_34 wl_0_7 sky130_rom_krom_rom_base_one_cell_81/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_45 wl_0_7 sky130_rom_krom_rom_base_zero_cell_45/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_56 wl_0_7 sky130_rom_krom_rom_base_zero_cell_56/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_67 wl_0_7 sky130_rom_krom_rom_base_zero_cell_67/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_78 wl_0_7 sky130_rom_krom_rom_base_zero_cell_78/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_89 wl_0_7 sky130_rom_krom_rom_base_zero_cell_89/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1110 wl_0_1 sky130_rom_krom_rom_base_one_cell_985/S
+ bl_0_15 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_308 wl_0_7 sky130_rom_krom_rom_base_one_cell_93/S
+ sky130_rom_krom_rom_base_one_cell_547/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_319 wl_0_7 sky130_rom_krom_rom_base_one_cell_319/D
+ bl_0_141 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_340 wl_0_5 sky130_rom_krom_rom_base_zero_cell_68/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1121 wl_0_0 sky130_rom_krom_rom_base_one_cell_993/S
+ bl_0_251 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1132 wl_0_0 sky130_rom_krom_rom_base_one_cell_1132/D
+ bl_0_224 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1143 wl_0_0 sky130_rom_krom_rom_base_one_cell_1143/D
+ bl_0_204 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1154 wl_0_0 sky130_rom_krom_rom_base_one_cell_1154/D
+ bl_0_186 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1165 wl_0_0 sky130_rom_krom_rom_base_one_cell_908/S
+ bl_0_167 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1176 wl_0_0 sky130_rom_krom_rom_base_one_cell_1176/D
+ bl_0_140 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1187 wl_0_0 sky130_rom_krom_rom_base_one_cell_1187/D
+ bl_0_121 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1198 wl_0_0 sky130_rom_krom_rom_base_one_cell_1198/D
+ bl_0_102 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_395 wl_0_5 sky130_rom_krom_rom_base_one_cell_985/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_384 wl_0_5 sky130_rom_krom_rom_base_one_cell_726/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_373 wl_0_5 sky130_rom_krom_rom_base_one_cell_719/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_362 wl_0_5 sky130_rom_krom_rom_base_one_cell_956/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_351 wl_0_5 sky130_rom_krom_rom_base_one_cell_826/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_831 wl_0_3 sky130_rom_krom_rom_base_one_cell_831/D
+ bl_0_75 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_820 wl_0_3 sky130_rom_krom_rom_base_one_cell_820/D
+ sky130_rom_krom_rom_base_one_cell_938/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_897 wl_0_2 sky130_rom_krom_rom_base_one_cell_897/D
+ sky130_rom_krom_rom_base_one_cell_897/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_886 wl_0_2 sky130_rom_krom_rom_base_one_cell_886/D
+ bl_0_206 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_875 wl_0_2 sky130_rom_krom_rom_base_one_cell_875/D
+ bl_0_233 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_864 wl_0_2 sky130_rom_krom_rom_base_one_cell_864/D
+ sky130_rom_krom_rom_base_one_cell_864/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_853 wl_0_3 sky130_rom_krom_rom_base_one_cell_853/D
+ sky130_rom_krom_rom_base_one_cell_982/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_842 wl_0_3 sky130_rom_krom_rom_base_one_cell_842/D
+ bl_0_45 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_105 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_313/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_116 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_51/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_127 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_325/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_138 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_63/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_149 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_69/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_170 wl_0_6 sky130_rom_krom_rom_base_one_cell_309/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_181 wl_0_6 sky130_rom_krom_rom_base_zero_cell_51/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_192 wl_0_6 sky130_rom_krom_rom_base_one_cell_566/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_672 wl_0_4 sky130_rom_krom_rom_base_one_cell_672/D
+ sky130_rom_krom_rom_base_one_cell_912/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_661 wl_0_4 sky130_rom_krom_rom_base_one_cell_661/D
+ bl_0_181 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_650 wl_0_4 sky130_rom_krom_rom_base_one_cell_650/D
+ sky130_rom_krom_rom_base_one_cell_767/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_694 wl_0_4 sky130_rom_krom_rom_base_one_cell_694/D
+ sky130_rom_krom_rom_base_one_cell_819/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_683 wl_0_4 sky130_rom_krom_rom_base_one_cell_683/D
+ sky130_rom_krom_rom_base_one_cell_928/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_480 wl_0_6 sky130_rom_krom_rom_base_one_cell_480/D
+ sky130_rom_krom_rom_base_one_cell_480/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_491 wl_0_6 sky130_rom_krom_rom_base_one_cell_491/D
+ sky130_rom_krom_rom_base_one_cell_604/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_906 wl_0_1 bl_0_40 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_917 wl_0_1 bl_0_22 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_928 wl_0_1 sky130_rom_krom_rom_base_one_cell_861/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_939 wl_0_0 bl_0_236 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_747 wl_0_2 bl_0_115 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_736 wl_0_2 sky130_rom_krom_rom_base_one_cell_561/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_725 wl_0_2 bl_0_152 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_714 wl_0_2 sky130_rom_krom_rom_base_one_cell_787/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_703 wl_0_2 sky130_rom_krom_rom_base_one_cell_777/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_769 wl_0_2 sky130_rom_krom_rom_base_zero_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_758 wl_0_2 sky130_rom_krom_rom_base_one_cell_821/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_588 wl_0_3 sky130_rom_krom_rom_base_one_cell_441/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_577 wl_0_3 sky130_rom_krom_rom_base_one_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_566 wl_0_3 sky130_rom_krom_rom_base_one_cell_893/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_555 wl_0_3 sky130_rom_krom_rom_base_one_cell_641/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_544 wl_0_3 sky130_rom_krom_rom_base_one_cell_871/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_533 wl_0_4 sky130_rom_krom_rom_base_one_cell_858/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_522 wl_0_4 sky130_rom_krom_rom_base_one_cell_851/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_511 wl_0_4 sky130_rom_krom_rom_base_one_cell_840/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_500 wl_0_4 sky130_rom_krom_rom_base_one_cell_833/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_599 wl_0_3 sky130_rom_krom_rom_base_one_cell_923/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_13 wl_0_7 sky130_rom_krom_rom_base_one_cell_29/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_24 wl_0_7 sky130_rom_krom_rom_base_one_cell_62/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_35 wl_0_7 sky130_rom_krom_rom_base_one_cell_84/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_46 wl_0_7 sky130_rom_krom_rom_base_zero_cell_46/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_57 wl_0_7 sky130_rom_krom_rom_base_zero_cell_57/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_68 wl_0_7 sky130_rom_krom_rom_base_zero_cell_68/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_79 wl_0_7 sky130_rom_krom_rom_base_zero_cell_79/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_309 wl_0_7 sky130_rom_krom_rom_base_one_cell_96/S
+ sky130_rom_krom_rom_base_one_cell_309/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1100 wl_0_1 sky130_rom_krom_rom_base_one_cell_970/S
+ sky130_rom_krom_rom_base_one_cell_1226/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1111 wl_0_1 sky130_rom_krom_rom_base_one_cell_857/S
+ bl_0_12 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1122 wl_0_0 sky130_rom_krom_rom_base_one_cell_5/S
+ bl_0_250 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1133 wl_0_0 sky130_rom_krom_rom_base_one_cell_1133/D
+ bl_0_223 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1144 wl_0_0 sky130_rom_krom_rom_base_one_cell_889/S
+ bl_0_202 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_330 wl_0_5 sky130_rom_krom_rom_base_one_cell_923/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_341 wl_0_5 sky130_rom_krom_rom_base_one_cell_459/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1155 wl_0_0 sky130_rom_krom_rom_base_one_cell_902/S
+ bl_0_184 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1166 wl_0_0 sky130_rom_krom_rom_base_one_cell_1166/D
+ bl_0_163 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1177 wl_0_0 sky130_rom_krom_rom_base_one_cell_1177/D
+ bl_0_139 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1188 wl_0_0 sky130_rom_krom_rom_base_one_cell_811/S
+ bl_0_118 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1199 wl_0_0 sky130_rom_krom_rom_base_one_cell_938/S
+ bl_0_96 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_396 wl_0_5 sky130_rom_krom_rom_base_one_cell_988/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_385 wl_0_5 sky130_rom_krom_rom_base_one_cell_847/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_374 wl_0_5 sky130_rom_krom_rom_base_one_cell_840/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_363 wl_0_5 sky130_rom_krom_rom_base_one_cell_957/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_352 wl_0_5 sky130_rom_krom_rom_base_zero_cell_80/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_854 wl_0_3 sky130_rom_krom_rom_base_one_cell_854/D
+ sky130_rom_krom_rom_base_one_cell_854/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_843 wl_0_3 sky130_rom_krom_rom_base_one_cell_843/D
+ sky130_rom_krom_rom_base_one_cell_968/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_832 wl_0_3 sky130_rom_krom_rom_base_one_cell_832/D
+ sky130_rom_krom_rom_base_one_cell_954/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_821 wl_0_3 sky130_rom_krom_rom_base_one_cell_821/D
+ sky130_rom_krom_rom_base_one_cell_821/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_810 wl_0_3 sky130_rom_krom_rom_base_one_cell_810/D
+ sky130_rom_krom_rom_base_one_cell_810/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_898 wl_0_2 sky130_rom_krom_rom_base_one_cell_898/D
+ bl_0_190 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_887 wl_0_2 sky130_rom_krom_rom_base_one_cell_887/D
+ sky130_rom_krom_rom_base_one_cell_887/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_876 wl_0_2 sky130_rom_krom_rom_base_one_cell_24/S
+ bl_0_231 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_865 wl_0_2 sky130_rom_krom_rom_base_one_cell_865/D
+ bl_0_248 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_106 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_314/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_117 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_321/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_128 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_326/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_139 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_331/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_160 wl_0_6 sky130_rom_krom_rom_base_one_cell_660/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_171 wl_0_6 sky130_rom_krom_rom_base_one_cell_97/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_182 wl_0_6 sky130_rom_krom_rom_base_zero_cell_53/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_193 wl_0_6 sky130_rom_krom_rom_base_zero_cell_62/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_695 wl_0_4 sky130_rom_krom_rom_base_one_cell_695/D
+ bl_0_98 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_684 wl_0_4 sky130_rom_krom_rom_base_one_cell_684/D
+ sky130_rom_krom_rom_base_one_cell_684/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_673 wl_0_4 sky130_rom_krom_rom_base_one_cell_673/D
+ sky130_rom_krom_rom_base_one_cell_673/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_662 wl_0_4 sky130_rom_krom_rom_base_one_cell_662/D
+ sky130_rom_krom_rom_base_one_cell_783/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_651 wl_0_4 sky130_rom_krom_rom_base_one_cell_651/D
+ sky130_rom_krom_rom_base_one_cell_769/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_640 wl_0_4 sky130_rom_krom_rom_base_one_cell_640/D
+ sky130_rom_krom_rom_base_one_cell_757/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_907 wl_0_1 sky130_rom_krom_rom_base_one_cell_494/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_918 wl_0_1 bl_0_21 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_929 wl_0_1 bl_0_1 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_470 wl_0_6 sky130_rom_krom_rom_base_zero_cell_74/S
+ sky130_rom_krom_rom_base_one_cell_698/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_481 wl_0_6 sky130_rom_krom_rom_base_one_cell_481/D
+ sky130_rom_krom_rom_base_one_cell_595/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_492 wl_0_6 sky130_rom_krom_rom_base_one_cell_492/D
+ sky130_rom_krom_rom_base_one_cell_723/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_759 wl_0_2 sky130_rom_krom_rom_base_zero_cell_75/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_748 wl_0_2 bl_0_114 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_737 wl_0_2 bl_0_129 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_726 wl_0_2 sky130_rom_krom_rom_base_one_cell_796/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_715 wl_0_2 sky130_rom_krom_rom_base_one_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_704 wl_0_2 sky130_rom_krom_rom_base_one_cell_778/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_589 wl_0_3 sky130_rom_krom_rom_base_one_cell_915/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_578 wl_0_3 sky130_rom_krom_rom_base_one_cell_909/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_567 wl_0_3 sky130_rom_krom_rom_base_one_cell_62/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_556 wl_0_3 bl_0_219 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_545 wl_0_3 sky130_rom_krom_rom_base_one_cell_872/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_534 wl_0_4 sky130_rom_krom_rom_base_one_cell_859/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_523 wl_0_4 sky130_rom_krom_rom_base_one_cell_503/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_512 wl_0_4 sky130_rom_krom_rom_base_one_cell_841/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_501 wl_0_4 sky130_rom_krom_rom_base_one_cell_834/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_14 wl_0_7 sky130_rom_krom_rom_base_one_cell_34/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_25 wl_0_7 sky130_rom_krom_rom_base_one_cell_64/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_36 wl_0_7 sky130_rom_krom_rom_base_one_cell_85/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_47 wl_0_7 sky130_rom_krom_rom_base_zero_cell_47/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_58 wl_0_7 sky130_rom_krom_rom_base_zero_cell_58/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_69 wl_0_7 sky130_rom_krom_rom_base_zero_cell_69/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_320 wl_0_5 sky130_rom_krom_rom_base_zero_cell_47/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1101 wl_0_1 sky130_rom_krom_rom_base_one_cell_973/S
+ bl_0_38 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1112 wl_0_1 sky130_rom_krom_rom_base_one_cell_737/S
+ sky130_rom_krom_rom_base_one_cell_1242/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1123 wl_0_0 sky130_rom_krom_rom_base_one_cell_994/S
+ bl_0_249 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1134 wl_0_0 sky130_rom_krom_rom_base_one_cell_1134/D
+ bl_0_221 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1145 wl_0_0 sky130_rom_krom_rom_base_one_cell_891/S
+ bl_0_199 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1156 wl_0_0 sky130_rom_krom_rom_base_one_cell_423/S
+ bl_0_183 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1167 wl_0_0 sky130_rom_krom_rom_base_one_cell_911/S
+ bl_0_162 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1178 wl_0_0 sky130_rom_krom_rom_base_one_cell_680/S
+ bl_0_138 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_331 wl_0_5 sky130_rom_krom_rom_base_zero_cell_57/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_342 wl_0_5 sky130_rom_krom_rom_base_zero_cell_69/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1189 wl_0_0 sky130_rom_krom_rom_base_one_cell_1189/D
+ bl_0_116 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_397 wl_0_5 sky130_rom_krom_rom_base_one_cell_989/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_386 wl_0_5 sky130_rom_krom_rom_base_one_cell_730/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_375 wl_0_5 sky130_rom_krom_rom_base_one_cell_722/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_364 wl_0_5 sky130_rom_krom_rom_base_zero_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_353 wl_0_5 sky130_rom_krom_rom_base_one_cell_827/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_888 wl_0_2 sky130_rom_krom_rom_base_one_cell_888/D
+ sky130_rom_krom_rom_base_one_cell_888/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_877 wl_0_2 sky130_rom_krom_rom_base_one_cell_877/D
+ bl_0_230 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_866 wl_0_2 sky130_rom_krom_rom_base_one_cell_866/D
+ bl_0_247 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_855 wl_0_3 sky130_rom_krom_rom_base_one_cell_855/D
+ sky130_rom_krom_rom_base_one_cell_983/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_844 wl_0_3 sky130_rom_krom_rom_base_one_cell_844/D
+ sky130_rom_krom_rom_base_one_cell_969/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_833 wl_0_3 sky130_rom_krom_rom_base_one_cell_833/D
+ sky130_rom_krom_rom_base_one_cell_833/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_822 wl_0_3 sky130_rom_krom_rom_base_one_cell_822/D
+ sky130_rom_krom_rom_base_one_cell_942/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_811 wl_0_3 sky130_rom_krom_rom_base_one_cell_811/D
+ sky130_rom_krom_rom_base_one_cell_811/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_800 wl_0_3 sky130_rom_krom_rom_base_one_cell_800/D
+ bl_0_142 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_899 wl_0_2 sky130_rom_krom_rom_base_one_cell_899/D
+ sky130_rom_krom_rom_base_one_cell_899/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_107 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_315/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_118 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_322/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_129 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_327/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_150 wl_0_6 sky130_rom_krom_rom_base_one_cell_771/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_161 wl_0_6 sky130_rom_krom_rom_base_one_cell_662/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_172 wl_0_6 sky130_rom_krom_rom_base_one_cell_98/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_183 wl_0_6 sky130_rom_krom_rom_base_one_cell_561/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_194 wl_0_6 sky130_rom_krom_rom_base_zero_cell_63/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_696 wl_0_4 sky130_rom_krom_rom_base_one_cell_696/D
+ sky130_rom_krom_rom_base_one_cell_937/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_685 wl_0_4 sky130_rom_krom_rom_base_one_cell_685/D
+ sky130_rom_krom_rom_base_one_cell_811/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_674 wl_0_4 sky130_rom_krom_rom_base_one_cell_674/D
+ sky130_rom_krom_rom_base_one_cell_796/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_663 wl_0_4 sky130_rom_krom_rom_base_one_cell_663/D
+ sky130_rom_krom_rom_base_one_cell_663/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_652 wl_0_4 sky130_rom_krom_rom_base_one_cell_652/D
+ sky130_rom_krom_rom_base_one_cell_891/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_641 wl_0_4 sky130_rom_krom_rom_base_one_cell_34/S
+ sky130_rom_krom_rom_base_one_cell_641/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_630 wl_0_4 sky130_rom_krom_rom_base_one_cell_630/D
+ sky130_rom_krom_rom_base_one_cell_748/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_908 wl_0_1 sky130_rom_krom_rom_base_one_cell_974/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_919 wl_0_1 sky130_rom_krom_rom_base_one_cell_982/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_460 wl_0_6 sky130_rom_krom_rom_base_one_cell_460/D
+ sky130_rom_krom_rom_base_one_cell_933/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_471 wl_0_6 sky130_rom_krom_rom_base_zero_cell_76/S
+ sky130_rom_krom_rom_base_one_cell_585/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_482 wl_0_6 sky130_rom_krom_rom_base_zero_cell_88/S
+ sky130_rom_krom_rom_base_one_cell_711/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_493 wl_0_6 sky130_rom_krom_rom_base_one_cell_493/D
+ sky130_rom_krom_rom_base_one_cell_724/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_290 wl_0_7 sky130_rom_krom_rom_base_one_cell_56/S
+ sky130_rom_krom_rom_base_one_cell_417/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_749 wl_0_2 sky130_rom_krom_rom_base_one_cell_457/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_738 wl_0_2 sky130_rom_krom_rom_base_one_cell_563/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_727 wl_0_2 sky130_rom_krom_rom_base_one_cell_441/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_716 wl_0_2 bl_0_165 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_705 wl_0_2 sky130_rom_krom_rom_base_one_cell_423/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_513 wl_0_4 sky130_rom_krom_rom_base_one_cell_844/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_502 wl_0_4 sky130_rom_krom_rom_base_one_cell_480/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_579 wl_0_3 bl_0_165 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_568 wl_0_3 sky130_rom_krom_rom_base_one_cell_897/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_557 wl_0_3 sky130_rom_krom_rom_base_one_cell_644/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_546 wl_0_3 sky130_rom_krom_rom_base_one_cell_874/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_535 wl_0_4 sky130_rom_krom_rom_base_one_cell_860/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_524 wl_0_4 sky130_rom_krom_rom_base_one_cell_852/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_15 wl_0_7 sky130_rom_krom_rom_base_one_cell_36/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_26 wl_0_7 sky130_rom_krom_rom_base_one_cell_66/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_37 wl_0_7 sky130_rom_krom_rom_base_one_cell_86/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_48 wl_0_7 sky130_rom_krom_rom_base_zero_cell_48/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_59 wl_0_7 sky130_rom_krom_rom_base_zero_cell_59/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_310 wl_0_5 sky130_rom_krom_rom_base_one_cell_667/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_321 wl_0_5 sky130_rom_krom_rom_base_one_cell_441/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_332 wl_0_5 sky130_rom_krom_rom_base_one_cell_806/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_343 wl_0_5 sky130_rom_krom_rom_base_one_cell_933/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1102 wl_0_1 sky130_rom_krom_rom_base_one_cell_847/S
+ bl_0_32 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1113 wl_0_1 sky130_rom_krom_rom_base_one_cell_989/S
+ sky130_rom_krom_rom_base_one_cell_1244/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1124 wl_0_0 sky130_rom_krom_rom_base_one_cell_868/S
+ bl_0_244 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1135 wl_0_0 sky130_rom_krom_rom_base_one_cell_1135/D
+ bl_0_220 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1146 wl_0_0 sky130_rom_krom_rom_base_one_cell_1146/D
+ bl_0_198 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1157 wl_0_0 sky130_rom_krom_rom_base_one_cell_1157/D
+ bl_0_182 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1168 wl_0_0 sky130_rom_krom_rom_base_one_cell_1168/D
+ bl_0_160 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1179 wl_0_0 sky130_rom_krom_rom_base_one_cell_1179/D
+ bl_0_137 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_354 wl_0_5 sky130_rom_krom_rom_base_one_cell_707/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_398 wl_0_5 sky130_rom_krom_rom_base_one_cell_739/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_387 wl_0_5 sky130_rom_krom_rom_base_one_cell_851/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_376 wl_0_5 sky130_rom_krom_rom_base_one_cell_723/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_365 wl_0_5 sky130_rom_krom_rom_base_one_cell_711/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_889 wl_0_2 sky130_rom_krom_rom_base_one_cell_889/D
+ sky130_rom_krom_rom_base_one_cell_889/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_878 wl_0_2 sky130_rom_krom_rom_base_one_cell_878/D
+ sky130_rom_krom_rom_base_one_cell_878/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_867 wl_0_2 sky130_rom_krom_rom_base_one_cell_867/D
+ sky130_rom_krom_rom_base_one_cell_996/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_856 wl_0_3 sky130_rom_krom_rom_base_one_cell_856/D
+ sky130_rom_krom_rom_base_one_cell_987/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_845 wl_0_3 sky130_rom_krom_rom_base_one_cell_845/D
+ sky130_rom_krom_rom_base_one_cell_845/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_834 wl_0_3 sky130_rom_krom_rom_base_one_cell_834/D
+ sky130_rom_krom_rom_base_one_cell_955/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_823 wl_0_3 sky130_rom_krom_rom_base_one_cell_823/D
+ sky130_rom_krom_rom_base_one_cell_943/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_812 wl_0_3 sky130_rom_krom_rom_base_one_cell_812/D
+ sky130_rom_krom_rom_base_one_cell_812/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_801 wl_0_3 sky130_rom_krom_rom_base_one_cell_801/D
+ sky130_rom_krom_rom_base_one_cell_801/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_108 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_48/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_119 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_52/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_140 wl_0_6 sky130_rom_krom_rom_base_one_cell_525/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_151 wl_0_6 sky130_rom_krom_rom_base_one_cell_534/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_162 wl_0_6 sky130_rom_krom_rom_base_one_cell_784/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_173 wl_0_6 sky130_rom_krom_rom_base_one_cell_673/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_184 wl_0_6 sky130_rom_krom_rom_base_zero_cell_56/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_195 wl_0_6 sky130_rom_krom_rom_base_one_cell_569/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_620 wl_0_5 sky130_rom_krom_rom_base_one_cell_620/D
+ sky130_rom_krom_rom_base_one_cell_859/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_697 wl_0_4 sky130_rom_krom_rom_base_one_cell_697/D
+ sky130_rom_krom_rom_base_one_cell_939/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_686 wl_0_4 sky130_rom_krom_rom_base_zero_cell_63/S
+ sky130_rom_krom_rom_base_one_cell_812/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_675 wl_0_4 sky130_rom_krom_rom_base_one_cell_675/D
+ sky130_rom_krom_rom_base_one_cell_915/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_664 wl_0_4 sky130_rom_krom_rom_base_one_cell_664/D
+ sky130_rom_krom_rom_base_one_cell_664/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_653 wl_0_4 sky130_rom_krom_rom_base_one_cell_653/D
+ sky130_rom_krom_rom_base_one_cell_893/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_642 wl_0_4 sky130_rom_krom_rom_base_one_cell_642/D
+ sky130_rom_krom_rom_base_one_cell_759/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_631 wl_0_4 sky130_rom_krom_rom_base_one_cell_631/D
+ sky130_rom_krom_rom_base_one_cell_750/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_450 wl_0_6 sky130_rom_krom_rom_base_one_cell_450/D
+ sky130_rom_krom_rom_base_one_cell_681/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_461 wl_0_6 sky130_rom_krom_rom_base_one_cell_461/D
+ sky130_rom_krom_rom_base_one_cell_575/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_472 wl_0_6 sky130_rom_krom_rom_base_one_cell_472/D
+ sky130_rom_krom_rom_base_one_cell_587/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_909 wl_0_1 sky130_rom_krom_rom_base_one_cell_975/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_483 wl_0_6 sky130_rom_krom_rom_base_zero_cell_90/S
+ sky130_rom_krom_rom_base_one_cell_596/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_494 wl_0_6 sky130_rom_krom_rom_base_one_cell_494/D
+ sky130_rom_krom_rom_base_one_cell_494/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_280 wl_0_7 sky130_rom_krom_rom_base_one_cell_42/S
+ sky130_rom_krom_rom_base_one_cell_527/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_291 wl_0_7 sky130_rom_krom_rom_base_one_cell_57/S
+ sky130_rom_krom_rom_base_one_cell_534/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_739 wl_0_2 sky130_rom_krom_rom_base_one_cell_327/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_728 wl_0_2 sky130_rom_krom_rom_base_one_cell_799/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_717 wl_0_2 sky130_rom_krom_rom_base_one_cell_792/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_706 wl_0_2 sky130_rom_krom_rom_base_one_cell_782/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_536 wl_0_4 sky130_rom_krom_rom_base_one_cell_861/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_525 wl_0_4 sky130_rom_krom_rom_base_one_cell_980/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_514 wl_0_4 sky130_rom_krom_rom_base_one_cell_494/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_503 wl_0_4 sky130_rom_krom_rom_base_one_cell_956/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_569 wl_0_3 sky130_rom_krom_rom_base_one_cell_901/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_558 wl_0_3 sky130_rom_krom_rom_base_one_cell_645/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_547 wl_0_3 bl_0_232 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_16 wl_0_7 sky130_rom_krom_rom_base_one_cell_38/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_27 wl_0_7 sky130_rom_krom_rom_base_one_cell_68/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_38 wl_0_7 sky130_rom_krom_rom_base_one_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_49 wl_0_7 sky130_rom_krom_rom_base_zero_cell_49/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_300 wl_0_5 sky130_rom_krom_rom_base_one_cell_423/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_311 wl_0_5 sky130_rom_krom_rom_base_one_cell_668/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_322 wl_0_5 sky130_rom_krom_rom_base_one_cell_798/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_333 wl_0_5 sky130_rom_krom_rom_base_one_cell_327/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_344 wl_0_5 sky130_rom_krom_rom_base_one_cell_693/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1103 wl_0_1 sky130_rom_krom_rom_base_one_cell_979/S
+ sky130_rom_krom_rom_base_one_cell_1231/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1114 wl_0_1 sky130_rom_krom_rom_base_one_cell_739/S
+ sky130_rom_krom_rom_base_one_cell_1245/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1125 wl_0_0 sky130_rom_krom_rom_base_one_cell_998/S
+ bl_0_242 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1136 wl_0_0 sky130_rom_krom_rom_base_one_cell_645/S
+ bl_0_217 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1147 wl_0_0 sky130_rom_krom_rom_base_one_cell_1147/D
+ bl_0_197 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1158 wl_0_0 sky130_rom_krom_rom_base_one_cell_783/S
+ bl_0_180 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1169 wl_0_0 sky130_rom_krom_rom_base_one_cell_1169/D
+ bl_0_159 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_388 wl_0_5 sky130_rom_krom_rom_base_one_cell_503/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_377 wl_0_5 sky130_rom_krom_rom_base_one_cell_724/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_366 wl_0_5 sky130_rom_krom_rom_base_zero_cell_89/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_355 wl_0_5 sky130_rom_krom_rom_base_one_cell_708/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_399 wl_0_4 sky130_rom_krom_rom_base_one_cell_742/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_813 wl_0_3 sky130_rom_krom_rom_base_one_cell_813/D
+ bl_0_114 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_802 wl_0_3 sky130_rom_krom_rom_base_one_cell_802/D
+ sky130_rom_krom_rom_base_one_cell_918/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_879 wl_0_2 sky130_rom_krom_rom_base_one_cell_879/D
+ sky130_rom_krom_rom_base_one_cell_879/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_868 wl_0_2 sky130_rom_krom_rom_base_one_cell_868/D
+ sky130_rom_krom_rom_base_one_cell_868/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_857 wl_0_3 sky130_rom_krom_rom_base_one_cell_857/D
+ sky130_rom_krom_rom_base_one_cell_857/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_846 wl_0_3 sky130_rom_krom_rom_base_one_cell_846/D
+ sky130_rom_krom_rom_base_one_cell_977/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_835 wl_0_3 sky130_rom_krom_rom_base_zero_cell_89/S
+ sky130_rom_krom_rom_base_one_cell_835/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_824 wl_0_3 sky130_rom_krom_rom_base_one_cell_824/D
+ sky130_rom_krom_rom_base_one_cell_944/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_109 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_316/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_130 wl_0_6 sky130_rom_krom_rom_base_zero_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_141 wl_0_6 sky130_rom_krom_rom_base_one_cell_38/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_152 wl_0_6 sky130_rom_krom_rom_base_one_cell_653/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_163 wl_0_6 sky130_rom_krom_rom_base_one_cell_542/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_174 wl_0_6 sky130_rom_krom_rom_base_zero_cell_46/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_185 wl_0_6 sky130_rom_krom_rom_base_zero_cell_57/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_196 wl_0_6 bl_0_115 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_654 wl_0_4 sky130_rom_krom_rom_base_one_cell_61/S
+ sky130_rom_krom_rom_base_one_cell_774/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_643 wl_0_4 sky130_rom_krom_rom_base_one_cell_643/D
+ bl_0_219 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_632 wl_0_4 sky130_rom_krom_rom_base_zero_cell_7/S
+ sky130_rom_krom_rom_base_one_cell_752/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_621 wl_0_5 sky130_rom_krom_rom_base_one_cell_621/D
+ sky130_rom_krom_rom_base_one_cell_860/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_610 wl_0_5 sky130_rom_krom_rom_base_one_cell_610/D
+ bl_0_22 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_698 wl_0_4 sky130_rom_krom_rom_base_one_cell_698/D
+ sky130_rom_krom_rom_base_one_cell_821/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_687 wl_0_4 sky130_rom_krom_rom_base_one_cell_687/D
+ sky130_rom_krom_rom_base_one_cell_687/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_676 wl_0_4 sky130_rom_krom_rom_base_one_cell_676/D
+ sky130_rom_krom_rom_base_one_cell_799/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_665 wl_0_4 sky130_rom_krom_rom_base_one_cell_665/D
+ sky130_rom_krom_rom_base_one_cell_787/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_440 wl_0_6 sky130_rom_krom_rom_base_one_cell_440/D
+ sky130_rom_krom_rom_base_one_cell_551/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_451 wl_0_6 sky130_rom_krom_rom_base_zero_cell_54/S
+ sky130_rom_krom_rom_base_one_cell_804/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_462 wl_0_6 sky130_rom_krom_rom_base_zero_cell_70/S
+ sky130_rom_krom_rom_base_one_cell_576/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_473 wl_0_6 sky130_rom_krom_rom_base_zero_cell_79/S
+ sky130_rom_krom_rom_base_one_cell_588/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_484 wl_0_6 sky130_rom_krom_rom_base_zero_cell_92/S
+ sky130_rom_krom_rom_base_one_cell_714/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_495 wl_0_6 sky130_rom_krom_rom_base_one_cell_495/D
+ sky130_rom_krom_rom_base_one_cell_973/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_729 wl_0_2 bl_0_145 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_718 wl_0_2 sky130_rom_krom_rom_base_one_cell_437/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_707 wl_0_2 bl_0_181 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_270 wl_0_7 sky130_rom_krom_rom_base_one_cell_27/S
+ sky130_rom_krom_rom_base_one_cell_521/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_281 wl_0_7 sky130_rom_krom_rom_base_one_cell_43/S
+ sky130_rom_krom_rom_base_one_cell_411/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_292 wl_0_7 sky130_rom_krom_rom_base_one_cell_58/S
+ sky130_rom_krom_rom_base_one_cell_653/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_559 wl_0_3 sky130_rom_krom_rom_base_one_cell_646/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_548 wl_0_3 sky130_rom_krom_rom_base_one_cell_24/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_537 wl_0_4 sky130_rom_krom_rom_base_one_cell_862/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_526 wl_0_4 bl_0_22 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_515 wl_0_4 sky130_rom_krom_rom_base_one_cell_973/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_504 wl_0_4 sky130_rom_krom_rom_base_one_cell_957/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_17 wl_0_7 sky130_rom_krom_rom_base_one_cell_39/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_28 wl_0_7 sky130_rom_krom_rom_base_one_cell_69/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_39 wl_0_7 sky130_rom_krom_rom_base_one_cell_89/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1104 wl_0_1 sky130_rom_krom_rom_base_one_cell_609/S
+ sky130_rom_krom_rom_base_one_cell_1233/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1115 wl_0_1 sky130_rom_krom_rom_base_one_cell_740/S
+ sky130_rom_krom_rom_base_one_cell_1246/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1126 wl_0_0 sky130_rom_krom_rom_base_one_cell_999/S
+ bl_0_239 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_301 wl_0_5 sky130_rom_krom_rom_base_one_cell_782/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_312 wl_0_5 sky130_rom_krom_rom_base_one_cell_669/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_323 wl_0_5 sky130_rom_krom_rom_base_one_cell_676/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_334 wl_0_5 sky130_rom_krom_rom_base_zero_cell_59/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1137 wl_0_0 sky130_rom_krom_rom_base_one_cell_1137/D
+ bl_0_216 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1148 wl_0_0 sky130_rom_krom_rom_base_one_cell_1148/D
+ bl_0_195 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1159 wl_0_0 sky130_rom_krom_rom_base_one_cell_784/S
+ bl_0_179 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_389 wl_0_5 sky130_rom_krom_rom_base_one_cell_852/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_378 wl_0_5 sky130_rom_krom_rom_base_one_cell_725/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_367 wl_0_5 sky130_rom_krom_rom_base_one_cell_714/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_356 wl_0_5 sky130_rom_krom_rom_base_zero_cell_82/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_345 wl_0_5 sky130_rom_krom_rom_base_one_cell_697/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_836 wl_0_3 sky130_rom_krom_rom_base_one_cell_836/D
+ sky130_rom_krom_rom_base_one_cell_836/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_825 wl_0_3 sky130_rom_krom_rom_base_one_cell_825/D
+ sky130_rom_krom_rom_base_one_cell_946/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_814 wl_0_3 sky130_rom_krom_rom_base_one_cell_814/D
+ sky130_rom_krom_rom_base_one_cell_930/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_803 wl_0_3 sky130_rom_krom_rom_base_one_cell_803/D
+ sky130_rom_krom_rom_base_one_cell_919/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_890 wl_0_1 sky130_rom_krom_rom_base_one_cell_958/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_869 wl_0_2 sky130_rom_krom_rom_base_zero_cell_6/S
+ sky130_rom_krom_rom_base_one_cell_998/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_858 wl_0_3 sky130_rom_krom_rom_base_one_cell_858/D
+ sky130_rom_krom_rom_base_one_cell_858/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_847 wl_0_3 sky130_rom_krom_rom_base_one_cell_847/D
+ sky130_rom_krom_rom_base_one_cell_847/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_120 wl_0_7 sky130_rom_krom_rom_base_one_cell_617/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_131 wl_0_6 sky130_rom_krom_rom_base_zero_cell_8/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_142 wl_0_6 sky130_rom_krom_rom_base_one_cell_646/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_153 wl_0_6 sky130_rom_krom_rom_base_one_cell_61/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_164 wl_0_6 sky130_rom_krom_rom_base_one_cell_663/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_175 wl_0_6 sky130_rom_krom_rom_base_zero_cell_47/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_186 wl_0_6 sky130_rom_krom_rom_base_one_cell_806/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_197 wl_0_6 sky130_rom_krom_rom_base_zero_cell_64/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_688 wl_0_4 sky130_rom_krom_rom_base_one_cell_688/D
+ sky130_rom_krom_rom_base_one_cell_929/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_677 wl_0_4 sky130_rom_krom_rom_base_one_cell_677/D
+ bl_0_145 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_666 wl_0_4 sky130_rom_krom_rom_base_one_cell_666/D
+ sky130_rom_krom_rom_base_one_cell_788/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_655 wl_0_4 sky130_rom_krom_rom_base_one_cell_655/D
+ sky130_rom_krom_rom_base_one_cell_897/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_644 wl_0_4 sky130_rom_krom_rom_base_one_cell_644/D
+ sky130_rom_krom_rom_base_one_cell_644/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_633 wl_0_4 sky130_rom_krom_rom_base_one_cell_633/D
+ sky130_rom_krom_rom_base_one_cell_871/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_622 wl_0_5 sky130_rom_krom_rom_base_one_cell_622/D
+ sky130_rom_krom_rom_base_one_cell_861/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_611 wl_0_5 sky130_rom_krom_rom_base_one_cell_611/D
+ sky130_rom_krom_rom_base_one_cell_733/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_600 wl_0_5 sky130_rom_krom_rom_base_one_cell_600/D
+ sky130_rom_krom_rom_base_one_cell_964/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_699 wl_0_4 sky130_rom_krom_rom_base_one_cell_699/D
+ sky130_rom_krom_rom_base_one_cell_822/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_430 wl_0_6 sky130_rom_krom_rom_base_one_cell_85/S
+ sky130_rom_krom_rom_base_one_cell_666/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_441 wl_0_6 sky130_rom_krom_rom_base_one_cell_441/D
+ sky130_rom_krom_rom_base_one_cell_441/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_452 wl_0_6 sky130_rom_krom_rom_base_zero_cell_55/S
+ sky130_rom_krom_rom_base_one_cell_923/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_463 wl_0_6 sky130_rom_krom_rom_base_one_cell_463/D
+ sky130_rom_krom_rom_base_one_cell_577/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_474 wl_0_6 sky130_rom_krom_rom_base_one_cell_474/D
+ sky130_rom_krom_rom_base_one_cell_827/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_485 wl_0_6 sky130_rom_krom_rom_base_zero_cell_94/S
+ sky130_rom_krom_rom_base_one_cell_715/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_496 wl_0_6 sky130_rom_krom_rom_base_one_cell_496/D
+ sky130_rom_krom_rom_base_one_cell_974/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_719 wl_0_2 sky130_rom_krom_rom_base_one_cell_309/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_708 wl_0_2 sky130_rom_krom_rom_base_one_cell_783/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_260 wl_0_7 sky130_rom_krom_rom_base_one_cell_9/S
+ sky130_rom_krom_rom_base_one_cell_394/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_271 wl_0_7 sky130_rom_krom_rom_base_one_cell_28/S
+ sky130_rom_krom_rom_base_one_cell_880/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_282 wl_0_7 sky130_rom_krom_rom_base_one_cell_46/S
+ sky130_rom_krom_rom_base_one_cell_649/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_293 wl_0_7 sky130_rom_krom_rom_base_one_cell_59/S
+ sky130_rom_krom_rom_base_one_cell_418/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_549 wl_0_3 sky130_rom_krom_rom_base_one_cell_877/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_538 wl_0_4 sky130_rom_krom_rom_base_one_cell_863/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_527 wl_0_4 sky130_rom_krom_rom_base_one_cell_853/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_516 wl_0_4 sky130_rom_krom_rom_base_one_cell_974/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_505 wl_0_4 sky130_rom_krom_rom_base_zero_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_18 wl_0_7 sky130_rom_krom_rom_base_one_cell_44/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_29 wl_0_7 sky130_rom_krom_rom_base_one_cell_71/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_302 wl_0_5 sky130_rom_krom_rom_base_one_cell_662/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1105 wl_0_1 sky130_rom_krom_rom_base_one_cell_850/S
+ bl_0_27 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1116 wl_0_1 sky130_rom_krom_rom_base_one_cell_858/S
+ bl_0_5 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1127 wl_0_0 sky130_rom_krom_rom_base_one_cell_1127/D
+ bl_0_238 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1138 wl_0_0 sky130_rom_krom_rom_base_one_cell_1138/D
+ bl_0_214 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1149 wl_0_0 sky130_rom_krom_rom_base_one_cell_1149/D
+ bl_0_194 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_313 wl_0_5 sky130_rom_krom_rom_base_one_cell_670/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_324 wl_0_5 sky130_rom_krom_rom_base_one_cell_445/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_335 wl_0_5 sky130_rom_krom_rom_base_one_cell_808/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_379 wl_0_5 sky130_rom_krom_rom_base_one_cell_494/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_368 wl_0_5 sky130_rom_krom_rom_base_zero_cell_93/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_357 wl_0_5 bl_0_73 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_346 wl_0_5 sky130_rom_krom_rom_base_one_cell_940/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_859 wl_0_3 sky130_rom_krom_rom_base_one_cell_859/D
+ bl_0_4 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_848 wl_0_3 sky130_rom_krom_rom_base_one_cell_848/D
+ sky130_rom_krom_rom_base_one_cell_978/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_837 wl_0_3 sky130_rom_krom_rom_base_one_cell_837/D
+ sky130_rom_krom_rom_base_one_cell_837/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_826 wl_0_3 sky130_rom_krom_rom_base_one_cell_826/D
+ sky130_rom_krom_rom_base_one_cell_947/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_815 wl_0_3 sky130_rom_krom_rom_base_zero_cell_68/S
+ sky130_rom_krom_rom_base_one_cell_931/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_804 wl_0_3 sky130_rom_krom_rom_base_one_cell_804/D
+ sky130_rom_krom_rom_base_one_cell_922/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_880 wl_0_1 sky130_rom_krom_rom_base_one_cell_948/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_891 wl_0_1 sky130_rom_krom_rom_base_one_cell_835/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_110 wl_0_7 sky130_rom_krom_rom_base_one_cell_502/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_121 wl_0_7 sky130_rom_krom_rom_base_one_cell_623/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_132 wl_0_6 sky130_rom_krom_rom_base_zero_cell_9/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_143 wl_0_6 sky130_rom_krom_rom_base_one_cell_527/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_154 wl_0_6 sky130_rom_krom_rom_base_one_cell_62/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_165 wl_0_6 sky130_rom_krom_rom_base_one_cell_81/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_176 wl_0_6 sky130_rom_krom_rom_base_one_cell_552/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_187 wl_0_6 sky130_rom_krom_rom_base_one_cell_327/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_198 wl_0_6 sky130_rom_krom_rom_base_one_cell_572/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_689 wl_0_4 sky130_rom_krom_rom_base_one_cell_689/D
+ sky130_rom_krom_rom_base_one_cell_814/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_678 wl_0_4 sky130_rom_krom_rom_base_one_cell_678/D
+ sky130_rom_krom_rom_base_one_cell_800/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_667 wl_0_4 sky130_rom_krom_rom_base_one_cell_667/D
+ sky130_rom_krom_rom_base_one_cell_790/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_656 wl_0_4 sky130_rom_krom_rom_base_one_cell_656/D
+ sky130_rom_krom_rom_base_one_cell_776/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_645 wl_0_4 sky130_rom_krom_rom_base_one_cell_38/S
+ sky130_rom_krom_rom_base_one_cell_645/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_634 wl_0_4 sky130_rom_krom_rom_base_zero_cell_9/S
+ sky130_rom_krom_rom_base_one_cell_872/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_623 wl_0_5 sky130_rom_krom_rom_base_one_cell_623/D
+ sky130_rom_krom_rom_base_one_cell_862/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_612 wl_0_5 sky130_rom_krom_rom_base_one_cell_612/D
+ sky130_rom_krom_rom_base_one_cell_734/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_601 wl_0_5 sky130_rom_krom_rom_base_one_cell_601/D
+ sky130_rom_krom_rom_base_one_cell_720/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_420 wl_0_6 sky130_rom_krom_rom_base_one_cell_64/S
+ sky130_rom_krom_rom_base_one_cell_775/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_431 wl_0_6 sky130_rom_krom_rom_base_one_cell_86/S
+ sky130_rom_krom_rom_base_one_cell_545/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_442 wl_0_6 sky130_rom_krom_rom_base_zero_cell_48/S
+ sky130_rom_krom_rom_base_one_cell_798/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_453 wl_0_6 sky130_rom_krom_rom_base_one_cell_453/D
+ sky130_rom_krom_rom_base_one_cell_563/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_464 wl_0_6 sky130_rom_krom_rom_base_zero_cell_71/S
+ sky130_rom_krom_rom_base_one_cell_578/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_475 wl_0_6 sky130_rom_krom_rom_base_zero_cell_81/S
+ sky130_rom_krom_rom_base_one_cell_589/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_486 wl_0_6 sky130_rom_krom_rom_base_one_cell_486/D
+ sky130_rom_krom_rom_base_one_cell_837/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_497 wl_0_6 sky130_rom_krom_rom_base_one_cell_497/D
+ sky130_rom_krom_rom_base_one_cell_975/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_250 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_385/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_261 wl_0_7 sky130_rom_krom_rom_base_one_cell_10/S
+ sky130_rom_krom_rom_base_one_cell_395/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_272 wl_0_7 sky130_rom_krom_rom_base_one_cell_30/S
+ sky130_rom_krom_rom_base_one_cell_405/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_709 wl_0_2 sky130_rom_krom_rom_base_one_cell_784/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_283 wl_0_7 sky130_rom_krom_rom_base_one_cell_47/S
+ sky130_rom_krom_rom_base_one_cell_530/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_294 wl_0_7 sky130_rom_krom_rom_base_one_cell_63/S
+ sky130_rom_krom_rom_base_one_cell_536/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_539 wl_0_3 sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_528 wl_0_4 sky130_rom_krom_rom_base_one_cell_854/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_517 wl_0_4 sky130_rom_krom_rom_base_one_cell_975/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_506 wl_0_4 sky130_rom_krom_rom_base_zero_cell_89/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_19 wl_0_7 sky130_rom_krom_rom_base_one_cell_45/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_303 wl_0_5 sky130_rom_krom_rom_base_one_cell_784/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_314 wl_0_5 sky130_rom_krom_rom_base_one_cell_437/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_325 wl_0_5 sky130_rom_krom_rom_base_one_cell_678/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_336 wl_0_5 sky130_rom_krom_rom_base_one_cell_682/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1106 wl_0_1 sky130_rom_krom_rom_base_one_cell_503/S
+ sky130_rom_krom_rom_base_one_cell_1235/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1117 wl_0_1 sky130_rom_krom_rom_base_one_cell_991/S
+ bl_0_0 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1128 wl_0_0 sky130_rom_krom_rom_base_one_cell_873/S
+ bl_0_235 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1139 wl_0_0 sky130_rom_krom_rom_base_one_cell_1139/D
+ bl_0_213 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_369 wl_0_5 sky130_rom_krom_rom_base_one_cell_715/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_358 wl_0_5 bl_0_72 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_347 wl_0_5 sky130_rom_krom_rom_base_one_cell_698/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_881 wl_0_1 bl_0_80 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_892 wl_0_1 sky130_rom_krom_rom_base_one_cell_959/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_870 wl_0_1 bl_0_98 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_849 wl_0_3 sky130_rom_krom_rom_base_one_cell_849/D
+ sky130_rom_krom_rom_base_one_cell_849/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_838 wl_0_3 sky130_rom_krom_rom_base_zero_cell_96/S
+ sky130_rom_krom_rom_base_one_cell_838/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_827 wl_0_3 sky130_rom_krom_rom_base_one_cell_827/D
+ sky130_rom_krom_rom_base_one_cell_948/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_816 wl_0_3 sky130_rom_krom_rom_base_one_cell_816/D
+ sky130_rom_krom_rom_base_one_cell_816/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_805 wl_0_3 sky130_rom_krom_rom_base_zero_cell_57/S
+ bl_0_129 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_100 wl_0_7 sky130_rom_krom_rom_base_one_cell_601/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_111 wl_0_7 sky130_rom_krom_rom_base_one_cell_851/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_122 wl_0_7 sky130_rom_krom_rom_base_one_cell_624/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_133 wl_0_6 sky130_rom_krom_rom_base_one_cell_755/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_144 wl_0_6 sky130_rom_krom_rom_base_one_cell_45/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_155 wl_0_6 sky130_rom_krom_rom_base_one_cell_536/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_166 wl_0_6 sky130_rom_krom_rom_base_one_cell_544/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_177 wl_0_6 sky130_rom_krom_rom_base_one_cell_553/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_188 wl_0_6 sky130_rom_krom_rom_base_zero_cell_58/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_199 wl_0_6 sky130_rom_krom_rom_base_zero_cell_68/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_602 wl_0_5 sky130_rom_krom_rom_base_one_cell_602/D
+ sky130_rom_krom_rom_base_one_cell_841/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_679 wl_0_4 sky130_rom_krom_rom_base_one_cell_679/D
+ sky130_rom_krom_rom_base_one_cell_679/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_668 wl_0_4 sky130_rom_krom_rom_base_one_cell_668/D
+ sky130_rom_krom_rom_base_one_cell_909/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_657 wl_0_4 sky130_rom_krom_rom_base_one_cell_657/D
+ sky130_rom_krom_rom_base_one_cell_778/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_646 wl_0_4 sky130_rom_krom_rom_base_one_cell_646/D
+ sky130_rom_krom_rom_base_one_cell_646/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_635 wl_0_4 sky130_rom_krom_rom_base_one_cell_635/D
+ sky130_rom_krom_rom_base_one_cell_874/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_624 wl_0_5 sky130_rom_krom_rom_base_one_cell_624/D
+ sky130_rom_krom_rom_base_one_cell_863/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_613 wl_0_5 sky130_rom_krom_rom_base_one_cell_613/D
+ sky130_rom_krom_rom_base_one_cell_986/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_410 wl_0_6 sky130_rom_krom_rom_base_one_cell_410/D
+ sky130_rom_krom_rom_base_one_cell_526/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_421 wl_0_6 sky130_rom_krom_rom_base_one_cell_69/S
+ sky130_rom_krom_rom_base_one_cell_539/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_432 wl_0_6 sky130_rom_krom_rom_base_one_cell_432/D
+ sky130_rom_krom_rom_base_one_cell_667/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_443 wl_0_6 sky130_rom_krom_rom_base_one_cell_443/D
+ sky130_rom_krom_rom_base_one_cell_676/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_454 wl_0_6 sky130_rom_krom_rom_base_one_cell_454/D
+ sky130_rom_krom_rom_base_one_cell_682/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_465 wl_0_6 sky130_rom_krom_rom_base_one_cell_465/D
+ sky130_rom_krom_rom_base_one_cell_693/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_476 wl_0_6 sky130_rom_krom_rom_base_one_cell_476/D
+ sky130_rom_krom_rom_base_one_cell_708/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_487 wl_0_6 sky130_rom_krom_rom_base_zero_cell_95/S
+ sky130_rom_krom_rom_base_one_cell_598/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_498 wl_0_6 sky130_rom_krom_rom_base_one_cell_498/D
+ sky130_rom_krom_rom_base_one_cell_605/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_240 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_380/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_251 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_386/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_262 wl_0_7 sky130_rom_krom_rom_base_one_cell_11/S
+ sky130_rom_krom_rom_base_one_cell_396/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_273 wl_0_7 sky130_rom_krom_rom_base_one_cell_31/S
+ sky130_rom_krom_rom_base_one_cell_273/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_284 wl_0_7 sky130_rom_krom_rom_base_one_cell_48/S
+ sky130_rom_krom_rom_base_one_cell_413/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_295 wl_0_7 sky130_rom_krom_rom_base_one_cell_65/S
+ sky130_rom_krom_rom_base_one_cell_537/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_518 wl_0_4 sky130_rom_krom_rom_base_one_cell_845/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_507 wl_0_4 sky130_rom_krom_rom_base_zero_cell_93/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_529 wl_0_4 sky130_rom_krom_rom_base_one_cell_985/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_304 wl_0_5 sky130_rom_krom_rom_base_one_cell_663/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_315 wl_0_5 sky130_rom_krom_rom_base_one_cell_309/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_326 wl_0_5 bl_0_141 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_337 wl_0_5 sky130_rom_krom_rom_base_zero_cell_63/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1107 wl_0_1 sky130_rom_krom_rom_base_one_cell_852/S
+ bl_0_24 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1118 wl_0_0 sky130_rom_krom_rom_base_one_cell_741/S
+ bl_0_255 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1129 wl_0_0 sky130_rom_krom_rom_base_one_cell_1129/D
+ bl_0_234 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_359 wl_0_5 sky130_rom_krom_rom_base_zero_cell_85/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_348 wl_0_5 sky130_rom_krom_rom_base_zero_cell_75/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_882 wl_0_1 bl_0_79 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_893 wl_0_1 sky130_rom_krom_rom_base_one_cell_960/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_871 wl_0_1 bl_0_97 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_860 wl_0_1 sky130_rom_krom_rom_base_one_cell_327/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_839 wl_0_3 sky130_rom_krom_rom_base_one_cell_839/D
+ bl_0_51 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_828 wl_0_3 sky130_rom_krom_rom_base_one_cell_828/D
+ bl_0_80 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_817 wl_0_3 sky130_rom_krom_rom_base_one_cell_817/D
+ sky130_rom_krom_rom_base_one_cell_934/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_806 wl_0_3 sky130_rom_krom_rom_base_one_cell_806/D
+ sky130_rom_krom_rom_base_one_cell_925/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_101 wl_0_7 sky130_rom_krom_rom_base_one_cell_722/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_112 wl_0_7 sky130_rom_krom_rom_base_one_cell_505/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_123 wl_0_6 sky130_rom_krom_rom_base_one_cell_626/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_134 wl_0_6 sky130_rom_krom_rom_base_one_cell_24/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_145 wl_0_6 sky130_rom_krom_rom_base_one_cell_649/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_156 wl_0_6 sky130_rom_krom_rom_base_one_cell_537/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_167 wl_0_6 sky130_rom_krom_rom_base_one_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_178 wl_0_6 sky130_rom_krom_rom_base_zero_cell_49/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_189 wl_0_6 sky130_rom_krom_rom_base_zero_cell_59/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_636 wl_0_4 sky130_rom_krom_rom_base_one_cell_636/D
+ bl_0_232 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_625 wl_0_4 sky130_rom_krom_rom_base_one_cell_625/D
+ sky130_rom_krom_rom_base_one_cell_741/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_614 wl_0_5 sky130_rom_krom_rom_base_one_cell_614/D
+ sky130_rom_krom_rom_base_one_cell_735/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_603 wl_0_5 sky130_rom_krom_rom_base_one_cell_603/D
+ sky130_rom_krom_rom_base_one_cell_721/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_690 wl_0_2 sky130_rom_krom_rom_base_one_cell_644/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_669 wl_0_4 sky130_rom_krom_rom_base_one_cell_669/D
+ bl_0_165 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_658 wl_0_4 sky130_rom_krom_rom_base_one_cell_658/D
+ sky130_rom_krom_rom_base_one_cell_779/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_647 wl_0_4 sky130_rom_krom_rom_base_one_cell_647/D
+ sky130_rom_krom_rom_base_one_cell_883/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_400 wl_0_6 sky130_rom_krom_rom_base_one_cell_400/D
+ sky130_rom_krom_rom_base_one_cell_635/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_411 wl_0_6 sky130_rom_krom_rom_base_one_cell_411/D
+ sky130_rom_krom_rom_base_one_cell_762/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_422 wl_0_6 sky130_rom_krom_rom_base_one_cell_71/S
+ sky130_rom_krom_rom_base_one_cell_781/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_433 wl_0_6 sky130_rom_krom_rom_base_one_cell_89/S
+ sky130_rom_krom_rom_base_one_cell_668/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_444 wl_0_6 sky130_rom_krom_rom_base_one_cell_444/D
+ sky130_rom_krom_rom_base_one_cell_554/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_455 wl_0_6 sky130_rom_krom_rom_base_zero_cell_61/S
+ sky130_rom_krom_rom_base_one_cell_567/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_466 wl_0_6 sky130_rom_krom_rom_base_one_cell_466/D
+ sky130_rom_krom_rom_base_one_cell_580/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_477 wl_0_6 sky130_rom_krom_rom_base_one_cell_477/D
+ sky130_rom_krom_rom_base_one_cell_592/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_488 wl_0_6 sky130_rom_krom_rom_base_zero_cell_98/S
+ sky130_rom_krom_rom_base_one_cell_600/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_499 wl_0_6 sky130_rom_krom_rom_base_one_cell_499/D
+ sky130_rom_krom_rom_base_one_cell_847/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_230 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_374/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_241 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_510/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_252 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_387/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_263 wl_0_7 sky130_rom_krom_rom_base_one_cell_14/S
+ sky130_rom_krom_rom_base_one_cell_518/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_274 wl_0_7 sky130_rom_krom_rom_base_one_cell_32/S
+ sky130_rom_krom_rom_base_one_cell_406/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_285 wl_0_7 sky130_rom_krom_rom_base_one_cell_49/S
+ sky130_rom_krom_rom_base_one_cell_414/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_296 wl_0_7 sky130_rom_krom_rom_base_one_cell_67/S
+ sky130_rom_krom_rom_base_one_cell_657/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_519 wl_0_4 sky130_rom_krom_rom_base_one_cell_847/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_508 wl_0_4 sky130_rom_krom_rom_base_one_cell_837/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1108 wl_0_1 sky130_rom_krom_rom_base_one_cell_981/S
+ sky130_rom_krom_rom_base_one_cell_1237/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_305 wl_0_5 sky130_rom_krom_rom_base_one_cell_664/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_316 wl_0_5 sky130_rom_krom_rom_base_one_cell_98/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_327 wl_0_5 sky130_rom_krom_rom_base_one_cell_680/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_338 wl_0_5 bl_0_115 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1119 wl_0_0 sky130_rom_krom_rom_base_one_cell_743/S
+ bl_0_253 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_349 wl_0_5 sky130_rom_krom_rom_base_one_cell_945/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_818 wl_0_3 sky130_rom_krom_rom_base_one_cell_818/D
+ sky130_rom_krom_rom_base_one_cell_818/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_807 wl_0_3 sky130_rom_krom_rom_base_one_cell_807/D
+ sky130_rom_krom_rom_base_one_cell_807/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_883 wl_0_1 sky130_rom_krom_rom_base_one_cell_951/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_894 wl_0_1 sky130_rom_krom_rom_base_one_cell_961/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_872 wl_0_1 sky130_rom_krom_rom_base_one_cell_938/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_861 wl_0_1 sky130_rom_krom_rom_base_one_cell_807/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_850 wl_0_1 sky130_rom_krom_rom_base_one_cell_799/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_829 wl_0_3 sky130_rom_krom_rom_base_one_cell_829/D
+ sky130_rom_krom_rom_base_one_cell_829/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_102 wl_0_7 sky130_rom_krom_rom_base_one_cell_493/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_113 wl_0_7 sky130_rom_krom_rom_base_one_cell_506/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_124 wl_0_6 sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_135 wl_0_6 sky130_rom_krom_rom_base_one_cell_521/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_146 wl_0_6 sky130_rom_krom_rom_base_one_cell_530/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_157 wl_0_6 sky130_rom_krom_rom_base_one_cell_66/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_168 wl_0_6 sky130_rom_krom_rom_base_one_cell_547/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_179 wl_0_6 bl_0_141 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_659 wl_0_4 sky130_rom_krom_rom_base_one_cell_659/D
+ sky130_rom_krom_rom_base_one_cell_780/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_648 wl_0_4 sky130_rom_krom_rom_base_one_cell_648/D
+ sky130_rom_krom_rom_base_one_cell_648/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_637 wl_0_4 sky130_rom_krom_rom_base_one_cell_637/D
+ sky130_rom_krom_rom_base_one_cell_877/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_626 wl_0_4 sky130_rom_krom_rom_base_one_cell_626/D
+ sky130_rom_krom_rom_base_one_cell_743/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_615 wl_0_5 sky130_rom_krom_rom_base_one_cell_615/D
+ sky130_rom_krom_rom_base_one_cell_736/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_604 wl_0_5 sky130_rom_krom_rom_base_one_cell_604/D
+ sky130_rom_krom_rom_base_one_cell_844/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_691 wl_0_2 sky130_rom_krom_rom_base_one_cell_645/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_680 wl_0_2 bl_0_240 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_401 wl_0_6 sky130_rom_krom_rom_base_one_cell_401/D
+ sky130_rom_krom_rom_base_one_cell_636/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_412 wl_0_6 sky130_rom_krom_rom_base_one_cell_44/S
+ sky130_rom_krom_rom_base_one_cell_528/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_423 wl_0_6 sky130_rom_krom_rom_base_one_cell_72/S
+ sky130_rom_krom_rom_base_one_cell_423/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_434 wl_0_6 sky130_rom_krom_rom_base_one_cell_434/D
+ sky130_rom_krom_rom_base_one_cell_669/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_445 wl_0_6 sky130_rom_krom_rom_base_one_cell_445/D
+ sky130_rom_krom_rom_base_one_cell_445/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_456 wl_0_6 sky130_rom_krom_rom_base_zero_cell_65/S
+ sky130_rom_krom_rom_base_one_cell_571/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_467 wl_0_6 sky130_rom_krom_rom_base_one_cell_467/D
+ sky130_rom_krom_rom_base_one_cell_940/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_478 wl_0_6 sky130_rom_krom_rom_base_one_cell_478/D
+ sky130_rom_krom_rom_base_one_cell_709/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_489 wl_0_6 sky130_rom_krom_rom_base_zero_cell_99/S
+ sky130_rom_krom_rom_base_one_cell_719/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_990 wl_0_2 sky130_rom_krom_rom_base_one_cell_990/D
+ bl_0_1 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_220 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_370/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_231 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_375/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_242 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_511/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_253 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_388/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_264 wl_0_7 sky130_rom_krom_rom_base_one_cell_15/S
+ sky130_rom_krom_rom_base_one_cell_397/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_275 wl_0_7 sky130_rom_krom_rom_base_one_cell_33/S
+ sky130_rom_krom_rom_base_one_cell_758/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_286 wl_0_7 sky130_rom_krom_rom_base_one_cell_50/S
+ sky130_rom_krom_rom_base_one_cell_415/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_297 wl_0_7 sky130_rom_krom_rom_base_one_cell_70/S
+ sky130_rom_krom_rom_base_one_cell_660/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_509 wl_0_4 sky130_rom_krom_rom_base_zero_cell_96/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1109 wl_0_1 sky130_rom_krom_rom_base_one_cell_854/S
+ sky130_rom_krom_rom_base_one_cell_1239/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_306 wl_0_5 sky130_rom_krom_rom_base_one_cell_905/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_317 wl_0_5 sky130_rom_krom_rom_base_one_cell_673/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_328 wl_0_5 sky130_rom_krom_rom_base_one_cell_681/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_339 wl_0_5 sky130_rom_krom_rom_base_one_cell_457/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_840 wl_0_1 sky130_rom_krom_rom_base_one_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_819 wl_0_3 sky130_rom_krom_rom_base_one_cell_819/D
+ sky130_rom_krom_rom_base_one_cell_936/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_808 wl_0_3 sky130_rom_krom_rom_base_one_cell_808/D
+ sky130_rom_krom_rom_base_one_cell_808/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_873 wl_0_1 sky130_rom_krom_rom_base_one_cell_821/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_884 wl_0_1 bl_0_75 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_895 wl_0_1 bl_0_56 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_862 wl_0_1 bl_0_124 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_851 wl_0_1 bl_0_145 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_103 wl_0_7 sky130_rom_krom_rom_base_one_cell_494/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_114 wl_0_7 sky130_rom_krom_rom_base_one_cell_507/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_125 wl_0_6 sky130_rom_krom_rom_base_one_cell_515/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_136 wl_0_6 sky130_rom_krom_rom_base_one_cell_880/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_147 wl_0_6 sky130_rom_krom_rom_base_one_cell_650/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_158 wl_0_6 sky130_rom_krom_rom_base_one_cell_657/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_169 wl_0_6 sky130_rom_krom_rom_base_one_cell_95/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_692 wl_0_2 sky130_rom_krom_rom_base_one_cell_760/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_681 wl_0_2 sky130_rom_krom_rom_base_one_cell_999/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_670 wl_0_3 sky130_rom_krom_rom_base_one_cell_739/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_649 wl_0_4 sky130_rom_krom_rom_base_one_cell_649/D
+ sky130_rom_krom_rom_base_one_cell_763/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_638 wl_0_4 sky130_rom_krom_rom_base_one_cell_638/D
+ sky130_rom_krom_rom_base_one_cell_878/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_627 wl_0_4 sky130_rom_krom_rom_base_one_cell_627/D
+ sky130_rom_krom_rom_base_one_cell_745/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_616 wl_0_5 sky130_rom_krom_rom_base_one_cell_616/D
+ sky130_rom_krom_rom_base_one_cell_737/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_605 wl_0_5 sky130_rom_krom_rom_base_one_cell_605/D
+ sky130_rom_krom_rom_base_one_cell_727/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_402 wl_0_6 sky130_rom_krom_rom_base_one_cell_25/S
+ sky130_rom_krom_rom_base_one_cell_637/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_413 wl_0_6 sky130_rom_krom_rom_base_one_cell_413/D
+ sky130_rom_krom_rom_base_one_cell_531/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_424 wl_0_6 sky130_rom_krom_rom_base_one_cell_424/D
+ sky130_rom_krom_rom_base_one_cell_782/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_435 wl_0_6 sky130_rom_krom_rom_base_one_cell_435/D
+ sky130_rom_krom_rom_base_one_cell_546/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_446 wl_0_6 sky130_rom_krom_rom_base_zero_cell_50/S
+ sky130_rom_krom_rom_base_one_cell_678/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_457 wl_0_6 sky130_rom_krom_rom_base_zero_cell_66/S
+ sky130_rom_krom_rom_base_one_cell_457/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_468 wl_0_6 sky130_rom_krom_rom_base_one_cell_468/D
+ sky130_rom_krom_rom_base_one_cell_583/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_479 wl_0_6 sky130_rom_krom_rom_base_zero_cell_86/S
+ sky130_rom_krom_rom_base_one_cell_593/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_991 wl_0_2 sky130_rom_krom_rom_base_one_cell_991/D
+ sky130_rom_krom_rom_base_one_cell_991/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_980 wl_0_2 sky130_rom_krom_rom_base_one_cell_980/D
+ sky130_rom_krom_rom_base_one_cell_980/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_210 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_365/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_221 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_726/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_232 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_505/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_243 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_615/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_254 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_623/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_265 wl_0_7 sky130_rom_krom_rom_base_one_cell_17/S
+ sky130_rom_krom_rom_base_one_cell_398/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_276 wl_0_7 sky130_rom_krom_rom_base_one_cell_35/S
+ sky130_rom_krom_rom_base_one_cell_407/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_287 wl_0_7 sky130_rom_krom_rom_base_one_cell_51/S
+ sky130_rom_krom_rom_base_one_cell_650/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_298 wl_0_7 sky130_rom_krom_rom_base_one_cell_73/S
+ sky130_rom_krom_rom_base_one_cell_424/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_307 wl_0_5 sky130_rom_krom_rom_base_one_cell_665/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_318 wl_0_5 sky130_rom_krom_rom_base_one_cell_913/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_329 wl_0_5 sky130_rom_krom_rom_base_one_cell_804/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_874 wl_0_1 sky130_rom_krom_rom_base_one_cell_942/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_863 wl_0_1 sky130_rom_krom_rom_base_one_cell_808/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_852 wl_0_1 bl_0_142 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_841 wl_0_1 sky130_rom_krom_rom_base_one_cell_908/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_830 wl_0_1 bl_0_190 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_809 wl_0_3 sky130_rom_krom_rom_base_one_cell_809/D
+ sky130_rom_krom_rom_base_one_cell_927/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_885 wl_0_1 sky130_rom_krom_rom_base_one_cell_952/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_896 wl_0_1 sky130_rom_krom_rom_base_one_cell_962/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_104 wl_0_7 sky130_rom_krom_rom_base_one_cell_496/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_115 wl_0_7 sky130_rom_krom_rom_base_one_cell_508/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_126 wl_0_6 sky130_rom_krom_rom_base_one_cell_7/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_137 wl_0_6 sky130_rom_krom_rom_base_one_cell_273/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_148 wl_0_6 sky130_rom_krom_rom_base_one_cell_52/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_159 wl_0_6 sky130_rom_krom_rom_base_one_cell_68/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_693 wl_0_2 sky130_rom_krom_rom_base_one_cell_761/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_682 wl_0_2 sky130_rom_krom_rom_base_one_cell_753/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_671 wl_0_3 sky130_rom_krom_rom_base_one_cell_740/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_660 wl_0_3 bl_0_22 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_639 wl_0_4 sky130_rom_krom_rom_base_one_cell_639/D
+ sky130_rom_krom_rom_base_one_cell_756/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_628 wl_0_4 sky130_rom_krom_rom_base_one_cell_628/D
+ sky130_rom_krom_rom_base_one_cell_865/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_617 wl_0_5 sky130_rom_krom_rom_base_one_cell_617/D
+ sky130_rom_krom_rom_base_one_cell_738/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_606 wl_0_5 sky130_rom_krom_rom_base_one_cell_606/D
+ sky130_rom_krom_rom_base_one_cell_728/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_403 wl_0_6 sky130_rom_krom_rom_base_one_cell_403/D
+ sky130_rom_krom_rom_base_one_cell_638/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_414 wl_0_6 sky130_rom_krom_rom_base_one_cell_414/D
+ sky130_rom_krom_rom_base_one_cell_765/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_425 wl_0_6 sky130_rom_krom_rom_base_one_cell_74/S
+ sky130_rom_krom_rom_base_one_cell_540/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_436 wl_0_6 sky130_rom_krom_rom_base_one_cell_92/S
+ sky130_rom_krom_rom_base_one_cell_670/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_447 wl_0_6 sky130_rom_krom_rom_base_one_cell_447/D
+ sky130_rom_krom_rom_base_one_cell_680/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_458 wl_0_6 sky130_rom_krom_rom_base_zero_cell_67/S
+ sky130_rom_krom_rom_base_one_cell_573/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_469 wl_0_6 sky130_rom_krom_rom_base_one_cell_469/D
+ sky130_rom_krom_rom_base_one_cell_584/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_490 wl_0_4 sky130_rom_krom_rom_base_zero_cell_75/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_992 wl_0_1 sky130_rom_krom_rom_base_one_cell_992/D
+ bl_0_254 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_981 wl_0_2 sky130_rom_krom_rom_base_one_cell_981/D
+ sky130_rom_krom_rom_base_one_cell_981/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_970 wl_0_2 sky130_rom_krom_rom_base_one_cell_970/D
+ sky130_rom_krom_rom_base_one_cell_970/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_200 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_361/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_211 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_722/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_222 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_371/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_233 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_376/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_244 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_616/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_255 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_624/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_266 wl_0_7 sky130_rom_krom_rom_base_one_cell_21/S
+ sky130_rom_krom_rom_base_one_cell_400/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_277 wl_0_7 sky130_rom_krom_rom_base_one_cell_37/S
+ sky130_rom_krom_rom_base_one_cell_525/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1090 wl_0_1 sky130_rom_krom_rom_base_one_cell_833/S
+ sky130_rom_krom_rom_base_one_cell_1213/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_288 wl_0_7 sky130_rom_krom_rom_base_one_cell_54/S
+ sky130_rom_krom_rom_base_one_cell_533/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_299 wl_0_7 sky130_rom_krom_rom_base_one_cell_75/S
+ sky130_rom_krom_rom_base_one_cell_662/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_308 wl_0_5 sky130_rom_krom_rom_base_one_cell_666/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_319 wl_0_5 sky130_rom_krom_rom_base_zero_cell_46/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_875 wl_0_1 bl_0_88 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_886 wl_0_1 bl_0_73 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_897 wl_0_1 bl_0_53 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_864 wl_0_1 sky130_rom_krom_rom_base_one_cell_811/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_853 wl_0_1 bl_0_141 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_842 wl_0_1 bl_0_166 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_831 wl_0_1 sky130_rom_krom_rom_base_one_cell_902/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_820 wl_0_1 sky130_rom_krom_rom_base_one_cell_528/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_105 wl_0_7 sky130_rom_krom_rom_base_one_cell_497/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_116 wl_0_7 sky130_rom_krom_rom_base_one_cell_510/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_127 wl_0_6 sky130_rom_krom_rom_base_zero_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_138 wl_0_6 sky130_rom_krom_rom_base_one_cell_758/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_149 wl_0_6 sky130_rom_krom_rom_base_one_cell_533/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_618 wl_0_5 sky130_rom_krom_rom_base_one_cell_618/D
+ sky130_rom_krom_rom_base_one_cell_740/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_607 wl_0_5 sky130_rom_krom_rom_base_one_cell_607/D
+ sky130_rom_krom_rom_base_one_cell_979/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_694 wl_0_2 sky130_rom_krom_rom_base_one_cell_646/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_683 wl_0_2 bl_0_232 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_672 wl_0_2 sky130_rom_krom_rom_base_one_cell_741/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_661 wl_0_3 bl_0_21 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_650 wl_0_3 sky130_rom_krom_rom_base_one_cell_972/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_629 wl_0_4 sky130_rom_krom_rom_base_one_cell_629/D
+ sky130_rom_krom_rom_base_one_cell_995/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_404 wl_0_6 sky130_rom_krom_rom_base_one_cell_29/S
+ sky130_rom_krom_rom_base_one_cell_639/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_415 wl_0_6 sky130_rom_krom_rom_base_one_cell_415/D
+ sky130_rom_krom_rom_base_one_cell_766/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_426 wl_0_6 sky130_rom_krom_rom_base_one_cell_77/S
+ sky130_rom_krom_rom_base_one_cell_541/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_437 wl_0_6 sky130_rom_krom_rom_base_one_cell_94/S
+ sky130_rom_krom_rom_base_one_cell_437/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_448 wl_0_6 sky130_rom_krom_rom_base_one_cell_448/D
+ sky130_rom_krom_rom_base_one_cell_558/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_459 wl_0_6 sky130_rom_krom_rom_base_one_cell_459/D
+ sky130_rom_krom_rom_base_one_cell_459/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_491 wl_0_4 sky130_rom_krom_rom_base_one_cell_945/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_480 wl_0_4 sky130_rom_krom_rom_base_zero_cell_68/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_993 wl_0_1 sky130_rom_krom_rom_base_one_cell_993/D
+ sky130_rom_krom_rom_base_one_cell_993/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_982 wl_0_2 sky130_rom_krom_rom_base_one_cell_982/D
+ sky130_rom_krom_rom_base_one_cell_982/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_971 wl_0_2 sky130_rom_krom_rom_base_one_cell_971/D
+ bl_0_41 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_960 wl_0_2 sky130_rom_krom_rom_base_one_cell_960/D
+ sky130_rom_krom_rom_base_one_cell_960/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_201 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_362/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_212 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_366/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_223 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_499/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_234 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_377/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_245 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_617/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_256 wl_0_7 sky130_rom_krom_rom_base_one_cell_1/S
+ sky130_rom_krom_rom_base_one_cell_390/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_267 wl_0_7 sky130_rom_krom_rom_base_one_cell_22/S
+ sky130_rom_krom_rom_base_one_cell_755/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_278 wl_0_7 sky130_rom_krom_rom_base_one_cell_40/S
+ sky130_rom_krom_rom_base_one_cell_410/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_289 wl_0_7 sky130_rom_krom_rom_base_one_cell_55/S
+ sky130_rom_krom_rom_base_one_cell_771/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1091 wl_0_1 sky130_rom_krom_rom_base_one_cell_955/S
+ bl_0_68 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1080 wl_0_1 sky130_rom_krom_rom_base_one_cell_940/S
+ sky130_rom_krom_rom_base_one_cell_1201/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_790 wl_0_3 sky130_rom_krom_rom_base_one_cell_790/D
+ sky130_rom_krom_rom_base_one_cell_908/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_309 wl_0_5 sky130_rom_krom_rom_base_one_cell_87/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_876 wl_0_1 bl_0_87 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_887 wl_0_1 bl_0_72 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_898 wl_0_1 bl_0_51 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_865 wl_0_1 bl_0_115 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_854 wl_0_1 sky130_rom_krom_rom_base_one_cell_680/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_843 wl_0_1 bl_0_165 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_832 wl_0_1 sky130_rom_krom_rom_base_one_cell_423/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_821 wl_0_1 bl_0_209 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_810 wl_0_1 bl_0_233 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_106 wl_0_7 sky130_rom_krom_rom_base_one_cell_726/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_117 wl_0_7 sky130_rom_krom_rom_base_one_cell_511/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_128 wl_0_6 sky130_rom_krom_rom_base_zero_cell_6/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_139 wl_0_6 sky130_rom_krom_rom_base_one_cell_34/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_640 wl_0_3 sky130_rom_krom_rom_base_one_cell_960/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_619 wl_0_5 sky130_rom_krom_rom_base_one_cell_619/D
+ sky130_rom_krom_rom_base_one_cell_858/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_608 wl_0_5 sky130_rom_krom_rom_base_one_cell_608/D
+ sky130_rom_krom_rom_base_one_cell_729/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_695 wl_0_2 sky130_rom_krom_rom_base_one_cell_528/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_684 wl_0_2 sky130_rom_krom_rom_base_one_cell_756/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_673 wl_0_2 sky130_rom_krom_rom_base_one_cell_992/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_662 wl_0_3 sky130_rom_krom_rom_base_one_cell_981/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_651 wl_0_3 sky130_rom_krom_rom_base_one_cell_494/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_405 wl_0_6 sky130_rom_krom_rom_base_one_cell_405/D
+ sky130_rom_krom_rom_base_one_cell_522/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_416 wl_0_6 sky130_rom_krom_rom_base_one_cell_53/S
+ sky130_rom_krom_rom_base_one_cell_532/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_427 wl_0_6 sky130_rom_krom_rom_base_one_cell_80/S
+ sky130_rom_krom_rom_base_one_cell_664/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_438 wl_0_6 sky130_rom_krom_rom_base_zero_cell_45/S
+ sky130_rom_krom_rom_base_one_cell_550/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_449 wl_0_6 sky130_rom_krom_rom_base_zero_cell_52/S
+ sky130_rom_krom_rom_base_one_cell_559/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1240 wl_0_0 sky130_rom_krom_rom_base_one_cell_983/S
+ bl_0_17 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_481 wl_0_4 sky130_rom_krom_rom_base_one_cell_459/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_470 wl_0_4 sky130_rom_krom_rom_base_one_cell_806/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_492 wl_0_4 sky130_rom_krom_rom_base_one_cell_826/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_994 wl_0_1 sky130_rom_krom_rom_base_one_cell_994/D
+ sky130_rom_krom_rom_base_one_cell_994/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_983 wl_0_2 sky130_rom_krom_rom_base_one_cell_983/D
+ sky130_rom_krom_rom_base_one_cell_983/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_972 wl_0_2 sky130_rom_krom_rom_base_one_cell_972/D
+ bl_0_40 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_961 wl_0_2 sky130_rom_krom_rom_base_zero_cell_93/S
+ sky130_rom_krom_rom_base_one_cell_961/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_950 wl_0_2 sky130_rom_krom_rom_base_one_cell_950/D
+ sky130_rom_krom_rom_base_one_cell_950/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_202 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_95/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_213 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_367/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_224 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_606/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_235 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_506/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_246 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_381/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_257 wl_0_7 sky130_rom_krom_rom_base_one_cell_2/S
+ sky130_rom_krom_rom_base_one_cell_626/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_268 wl_0_7 sky130_rom_krom_rom_base_one_cell_23/S
+ sky130_rom_krom_rom_base_one_cell_401/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_279 wl_0_7 sky130_rom_krom_rom_base_one_cell_41/S
+ sky130_rom_krom_rom_base_one_cell_646/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1081 wl_0_1 sky130_rom_krom_rom_base_one_cell_941/S
+ sky130_rom_krom_rom_base_one_cell_1202/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1092 wl_0_1 sky130_rom_krom_rom_base_one_cell_957/S
+ bl_0_65 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1070 wl_0_1 sky130_rom_krom_rom_base_one_cell_931/S
+ bl_0_109 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_90 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_90/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_791 wl_0_3 sky130_rom_krom_rom_base_one_cell_791/D
+ sky130_rom_krom_rom_base_one_cell_910/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_780 wl_0_3 sky130_rom_krom_rom_base_one_cell_780/D
+ sky130_rom_krom_rom_base_one_cell_900/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_822 wl_0_1 bl_0_208 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_811 wl_0_1 bl_0_232 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_800 wl_0_1 sky130_rom_krom_rom_base_one_cell_741/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_877 wl_0_1 sky130_rom_krom_rom_base_one_cell_945/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_888 wl_0_1 sky130_rom_krom_rom_base_one_cell_480/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_899 wl_0_1 bl_0_50 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_866 wl_0_1 bl_0_114 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_855 wl_0_1 bl_0_136 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_844 wl_0_1 sky130_rom_krom_rom_base_one_cell_911/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_833 wl_0_1 bl_0_181 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_107 wl_0_7 sky130_rom_krom_rom_base_one_cell_499/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_118 wl_0_7 sky130_rom_krom_rom_base_one_cell_615/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_129 wl_0_6 sky130_rom_krom_rom_base_one_cell_518/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_674 wl_0_2 sky130_rom_krom_rom_base_one_cell_743/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_663 wl_0_3 sky130_rom_krom_rom_base_one_cell_984/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_652 wl_0_3 sky130_rom_krom_rom_base_one_cell_973/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_641 wl_0_3 sky130_rom_krom_rom_base_zero_cell_93/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_630 wl_0_3 bl_0_73 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_609 wl_0_5 sky130_rom_krom_rom_base_one_cell_609/D
+ sky130_rom_krom_rom_base_one_cell_609/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_696 wl_0_2 sky130_rom_krom_rom_base_one_cell_648/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_685 wl_0_2 bl_0_225 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_406 wl_0_6 sky130_rom_krom_rom_base_one_cell_406/D
+ sky130_rom_krom_rom_base_one_cell_523/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_417 wl_0_6 sky130_rom_krom_rom_base_one_cell_417/D
+ sky130_rom_krom_rom_base_one_cell_652/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_428 wl_0_6 sky130_rom_krom_rom_base_one_cell_428/D
+ sky130_rom_krom_rom_base_one_cell_905/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_439 wl_0_6 sky130_rom_krom_rom_base_one_cell_439/D
+ sky130_rom_krom_rom_base_one_cell_913/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1241 wl_0_0 sky130_rom_krom_rom_base_one_cell_987/S
+ bl_0_13 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1230 wl_0_0 sky130_rom_krom_rom_base_one_cell_845/S
+ bl_0_35 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_493 wl_0_4 sky130_rom_krom_rom_base_one_cell_827/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_482 wl_0_4 sky130_rom_krom_rom_base_one_cell_932/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_471 wl_0_4 sky130_rom_krom_rom_base_one_cell_327/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_460 wl_0_4 sky130_rom_krom_rom_base_one_cell_801/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_940 wl_0_2 sky130_rom_krom_rom_base_one_cell_940/D
+ sky130_rom_krom_rom_base_one_cell_940/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_995 wl_0_1 sky130_rom_krom_rom_base_one_cell_995/D
+ bl_0_246 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_984 wl_0_2 sky130_rom_krom_rom_base_one_cell_984/D
+ bl_0_16 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_973 wl_0_2 sky130_rom_krom_rom_base_one_cell_973/D
+ sky130_rom_krom_rom_base_one_cell_973/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_962 wl_0_2 sky130_rom_krom_rom_base_one_cell_962/D
+ sky130_rom_krom_rom_base_one_cell_962/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_951 wl_0_2 sky130_rom_krom_rom_base_one_cell_951/D
+ sky130_rom_krom_rom_base_one_cell_951/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_203 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_96/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_214 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_493/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_225 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_372/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1071 wl_0_1 sky130_rom_krom_rom_base_one_cell_459/S
+ sky130_rom_krom_rom_base_one_cell_1194/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1060 wl_0_1 sky130_rom_krom_rom_base_one_cell_925/S
+ bl_0_127 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_236 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_507/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_247 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_382/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_258 wl_0_7 sky130_rom_krom_rom_base_one_cell_6/S
+ sky130_rom_krom_rom_base_one_cell_515/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_269 wl_0_7 sky130_rom_krom_rom_base_one_cell_26/S
+ sky130_rom_krom_rom_base_one_cell_403/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_290 wl_0_5 sky130_rom_krom_rom_base_one_cell_652/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1082 wl_0_1 sky130_rom_krom_rom_base_one_cell_584/S
+ sky130_rom_krom_rom_base_one_cell_1203/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1093 wl_0_1 sky130_rom_krom_rom_base_zero_cell_87/S
+ sky130_rom_krom_rom_base_one_cell_1217/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_80 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_80/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_91 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_91/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_781 wl_0_3 sky130_rom_krom_rom_base_one_cell_781/D
+ sky130_rom_krom_rom_base_one_cell_902/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_770 wl_0_3 sky130_rom_krom_rom_base_one_cell_770/D
+ bl_0_201 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_792 wl_0_3 sky130_rom_krom_rom_base_one_cell_792/D
+ sky130_rom_krom_rom_base_one_cell_792/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_856 wl_0_1 sky130_rom_krom_rom_base_one_cell_921/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_845 wl_0_1 bl_0_158 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_834 wl_0_1 sky130_rom_krom_rom_base_one_cell_783/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_823 wl_0_1 bl_0_206 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_812 wl_0_1 bl_0_231 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_801 wl_0_1 sky130_rom_krom_rom_base_one_cell_743/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_878 wl_0_1 sky130_rom_krom_rom_base_one_cell_946/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_889 wl_0_1 sky130_rom_krom_rom_base_one_cell_956/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_867 wl_0_1 sky130_rom_krom_rom_base_one_cell_457/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_108 wl_0_7 sky130_rom_krom_rom_base_one_cell_606/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_119 wl_0_7 sky130_rom_krom_rom_base_one_cell_616/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_697 wl_0_2 bl_0_209 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_686 wl_0_2 sky130_rom_krom_rom_base_one_cell_273/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_675 wl_0_2 sky130_rom_krom_rom_base_one_cell_993/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_664 wl_0_3 sky130_rom_krom_rom_base_one_cell_985/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_653 wl_0_3 sky130_rom_krom_rom_base_one_cell_974/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_642 wl_0_3 bl_0_56 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_631 wl_0_3 bl_0_72 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_620 wl_0_3 sky130_rom_krom_rom_base_one_cell_940/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_407 wl_0_6 sky130_rom_krom_rom_base_one_cell_407/D
+ sky130_rom_krom_rom_base_one_cell_524/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_418 wl_0_6 sky130_rom_krom_rom_base_one_cell_418/D
+ sky130_rom_krom_rom_base_one_cell_772/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1242 wl_0_0 sky130_rom_krom_rom_base_one_cell_1242/D
+ bl_0_11 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1231 wl_0_0 sky130_rom_krom_rom_base_one_cell_1231/D
+ bl_0_30 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1220 wl_0_0 sky130_rom_krom_rom_base_one_cell_1220/D
+ bl_0_59 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_429 wl_0_6 sky130_rom_krom_rom_base_one_cell_84/S
+ sky130_rom_krom_rom_base_one_cell_665/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_494 wl_0_4 sky130_rom_krom_rom_base_zero_cell_82/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_483 wl_0_4 sky130_rom_krom_rom_base_one_cell_933/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_472 wl_0_4 sky130_rom_krom_rom_base_one_cell_807/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_461 wl_0_4 sky130_rom_krom_rom_base_one_cell_802/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_450 wl_0_4 sky130_rom_krom_rom_base_one_cell_794/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_974 wl_0_2 sky130_rom_krom_rom_base_one_cell_974/D
+ sky130_rom_krom_rom_base_one_cell_974/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_963 wl_0_2 sky130_rom_krom_rom_base_one_cell_963/D
+ bl_0_53 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_952 wl_0_2 sky130_rom_krom_rom_base_one_cell_952/D
+ sky130_rom_krom_rom_base_one_cell_952/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_941 wl_0_2 sky130_rom_krom_rom_base_one_cell_941/D
+ sky130_rom_krom_rom_base_one_cell_941/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_930 wl_0_2 sky130_rom_krom_rom_base_one_cell_930/D
+ sky130_rom_krom_rom_base_one_cell_930/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_996 wl_0_1 sky130_rom_krom_rom_base_one_cell_996/D
+ bl_0_245 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_985 wl_0_2 sky130_rom_krom_rom_base_one_cell_985/D
+ sky130_rom_krom_rom_base_one_cell_985/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_204 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_97/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_215 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_368/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_226 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_608/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_237 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_508/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_248 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_383/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_259 wl_0_7 sky130_rom_krom_rom_base_one_cell_8/S
+ sky130_rom_krom_rom_base_one_cell_393/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1083 wl_0_1 sky130_rom_krom_rom_base_zero_cell_75/S
+ bl_0_90 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1094 wl_0_1 sky130_rom_krom_rom_base_one_cell_711/S
+ bl_0_62 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1072 wl_0_1 sky130_rom_krom_rom_base_one_cell_932/S
+ sky130_rom_krom_rom_base_one_cell_1195/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1061 wl_0_1 sky130_rom_krom_rom_base_one_cell_927/S
+ bl_0_122 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1050 wl_0_1 sky130_rom_krom_rom_base_one_cell_916/S
+ bl_0_147 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_280 wl_0_5 sky130_rom_krom_rom_base_one_cell_38/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_291 wl_0_5 sky130_rom_krom_rom_base_one_cell_653/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_70 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_70/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_81 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_81/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_92 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_92/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_793 wl_0_3 sky130_rom_krom_rom_base_one_cell_98/S
+ sky130_rom_krom_rom_base_one_cell_793/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_782 wl_0_3 sky130_rom_krom_rom_base_one_cell_782/D
+ sky130_rom_krom_rom_base_one_cell_782/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_771 wl_0_3 sky130_rom_krom_rom_base_one_cell_771/D
+ sky130_rom_krom_rom_base_one_cell_890/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_760 wl_0_3 sky130_rom_krom_rom_base_one_cell_760/D
+ sky130_rom_krom_rom_base_one_cell_760/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_590 wl_0_5 sky130_rom_krom_rom_base_one_cell_590/D
+ sky130_rom_krom_rom_base_one_cell_706/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_879 wl_0_1 sky130_rom_krom_rom_base_one_cell_703/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_868 wl_0_1 bl_0_106 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_857 wl_0_1 sky130_rom_krom_rom_base_one_cell_561/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_846 wl_0_1 sky130_rom_krom_rom_base_one_cell_913/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_835 wl_0_1 sky130_rom_krom_rom_base_one_cell_784/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_824 wl_0_1 sky130_rom_krom_rom_base_one_cell_889/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_813 wl_0_1 bl_0_230 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_802 wl_0_1 sky130_rom_krom_rom_base_one_cell_864/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_109 wl_0_7 sky130_rom_krom_rom_base_one_cell_608/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_698 wl_0_2 bl_0_208 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_687 wl_0_2 sky130_rom_krom_rom_base_one_cell_641/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_676 wl_0_2 sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_665 wl_0_3 sky130_rom_krom_rom_base_one_cell_986/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_654 wl_0_3 sky130_rom_krom_rom_base_one_cell_975/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_643 wl_0_3 sky130_rom_krom_rom_base_one_cell_962/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_632 wl_0_3 sky130_rom_krom_rom_base_zero_cell_85/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_621 wl_0_3 sky130_rom_krom_rom_base_one_cell_941/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_610 wl_0_3 sky130_rom_krom_rom_base_one_cell_573/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_408 wl_0_6 sky130_rom_krom_rom_base_one_cell_36/S
+ sky130_rom_krom_rom_base_one_cell_643/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_419 wl_0_6 sky130_rom_krom_rom_base_one_cell_60/S
+ sky130_rom_krom_rom_base_one_cell_535/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1243 wl_0_0 sky130_rom_krom_rom_base_one_cell_988/S
+ bl_0_9 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1232 wl_0_0 sky130_rom_krom_rom_base_one_cell_849/S
+ bl_0_29 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1221 wl_0_0 sky130_rom_krom_rom_base_one_cell_960/S
+ bl_0_58 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1210 wl_0_0 sky130_rom_krom_rom_base_one_cell_1210/D
+ bl_0_77 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_495 wl_0_4 sky130_rom_krom_rom_base_one_cell_831/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_484 wl_0_4 sky130_rom_krom_rom_base_one_cell_817/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_473 wl_0_4 sky130_rom_krom_rom_base_zero_cell_59/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_462 wl_0_4 sky130_rom_krom_rom_base_one_cell_803/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_451 wl_0_4 sky130_rom_krom_rom_base_one_cell_913/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_440 wl_0_4 sky130_rom_krom_rom_base_one_cell_543/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_997 wl_0_1 sky130_rom_krom_rom_base_one_cell_997/D
+ bl_0_243 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_986 wl_0_2 sky130_rom_krom_rom_base_one_cell_986/D
+ bl_0_14 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_975 wl_0_2 sky130_rom_krom_rom_base_one_cell_975/D
+ sky130_rom_krom_rom_base_one_cell_975/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_964 wl_0_2 sky130_rom_krom_rom_base_one_cell_964/D
+ bl_0_50 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_953 wl_0_2 sky130_rom_krom_rom_base_zero_cell_85/S
+ sky130_rom_krom_rom_base_one_cell_953/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_942 wl_0_2 sky130_rom_krom_rom_base_one_cell_942/D
+ sky130_rom_krom_rom_base_one_cell_942/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_931 wl_0_2 sky130_rom_krom_rom_base_one_cell_931/D
+ sky130_rom_krom_rom_base_one_cell_931/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_920 wl_0_2 sky130_rom_krom_rom_base_one_cell_920/D
+ sky130_rom_krom_rom_base_one_cell_920/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_205 precharge gnd_uq0 sky130_rom_krom_rom_base_zero_cell_98/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_216 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_494/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_227 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_373/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_238 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_378/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_249 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_384/D
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_270 wl_0_5 sky130_rom_krom_rom_base_one_cell_636/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_281 wl_0_5 sky130_rom_krom_rom_base_one_cell_760/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_1084 wl_0_1 sky130_rom_krom_rom_base_one_cell_947/S
+ bl_0_84 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1095 wl_0_1 sky130_rom_krom_rom_base_one_cell_836/S
+ sky130_rom_krom_rom_base_one_cell_1220/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1073 wl_0_1 sky130_rom_krom_rom_base_one_cell_816/S
+ bl_0_104 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1062 wl_0_1 sky130_rom_krom_rom_base_one_cell_810/S
+ sky130_rom_krom_rom_base_one_cell_1187/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1051 wl_0_1 sky130_rom_krom_rom_base_one_cell_917/S
+ sky130_rom_krom_rom_base_one_cell_1174/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1040 wl_0_1 sky130_rom_krom_rom_base_one_cell_792/S
+ sky130_rom_krom_rom_base_one_cell_1166/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_292 wl_0_5 sky130_rom_krom_rom_base_one_cell_772/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_60 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_60/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_71 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_71/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_82 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_82/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_93 precharge gnd_uq0 sky130_rom_krom_rom_base_one_cell_93/S
+ gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_794 wl_0_3 sky130_rom_krom_rom_base_one_cell_794/D
+ sky130_rom_krom_rom_base_one_cell_794/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_783 wl_0_3 sky130_rom_krom_rom_base_one_cell_783/D
+ sky130_rom_krom_rom_base_one_cell_783/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_772 wl_0_3 sky130_rom_krom_rom_base_one_cell_772/D
+ bl_0_196 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_761 wl_0_3 sky130_rom_krom_rom_base_one_cell_761/D
+ sky130_rom_krom_rom_base_one_cell_761/S gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_750 wl_0_3 sky130_rom_krom_rom_base_one_cell_750/D
+ sky130_rom_krom_rom_base_one_cell_997/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_1050 wl_0_0 bl_0_10 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_580 wl_0_5 sky130_rom_krom_rom_base_one_cell_580/D
+ sky130_rom_krom_rom_base_one_cell_695/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_591 wl_0_5 sky130_rom_krom_rom_base_one_cell_591/D
+ sky130_rom_krom_rom_base_one_cell_831/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_869 wl_0_1 sky130_rom_krom_rom_base_one_cell_933/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_858 wl_0_1 sky130_rom_krom_rom_base_one_cell_923/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_847 wl_0_1 bl_0_152 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_836 wl_0_1 sky130_rom_krom_rom_base_one_cell_785/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_825 wl_0_1 bl_0_201 gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_814 wl_0_1 sky130_rom_krom_rom_base_one_cell_879/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_803 wl_0_1 sky130_rom_krom_rom_base_one_cell_5/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_622 wl_0_3 sky130_rom_krom_rom_base_one_cell_584/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_611 wl_0_3 sky130_rom_krom_rom_base_one_cell_459/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_600 wl_0_3 sky130_rom_krom_rom_base_one_cell_924/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_699 wl_0_2 sky130_rom_krom_rom_base_one_cell_766/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_688 wl_0_2 sky130_rom_krom_rom_base_one_cell_759/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_677 wl_0_2 sky130_rom_krom_rom_base_one_cell_994/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_666 wl_0_3 sky130_rom_krom_rom_base_one_cell_737/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_655 wl_0_3 sky130_rom_krom_rom_base_one_cell_976/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_644 wl_0_3 sky130_rom_krom_rom_base_one_cell_963/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_633 wl_0_3 sky130_rom_krom_rom_base_one_cell_480/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_one_cell_409 wl_0_6 sky130_rom_krom_rom_base_one_cell_39/S
+ sky130_rom_krom_rom_base_one_cell_760/D gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1200 wl_0_0 sky130_rom_krom_rom_base_one_cell_1200/D
+ bl_0_95 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1244 wl_0_0 sky130_rom_krom_rom_base_one_cell_1244/D
+ bl_0_8 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1233 wl_0_0 sky130_rom_krom_rom_base_one_cell_1233/D
+ bl_0_28 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1222 wl_0_0 sky130_rom_krom_rom_base_one_cell_961/S
+ bl_0_57 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_one_cell_1211 wl_0_0 sky130_rom_krom_rom_base_one_cell_951/S
+ bl_0_76 gnd sky130_rom_krom_rom_base_one_cell
Xsky130_rom_krom_rom_base_zero_cell_463 wl_0_4 sky130_rom_krom_rom_base_one_cell_920/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_452 wl_0_4 sky130_rom_krom_rom_base_zero_cell_46/S
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_441 wl_0_4 sky130_rom_krom_rom_base_one_cell_904/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_430 wl_0_4 sky130_rom_krom_rom_base_one_cell_773/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_496 wl_0_4 sky130_rom_krom_rom_base_one_cell_952/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_485 wl_0_4 sky130_rom_krom_rom_base_one_cell_818/D
+ gnd sky130_rom_krom_rom_base_zero_cell
Xsky130_rom_krom_rom_base_zero_cell_474 wl_0_4 sky130_rom_krom_rom_base_one_cell_808/D
+ gnd sky130_rom_krom_rom_base_zero_cell
.ends

.subckt sky130_rom_krom_pinv_dec_3 A Z vdd w_692_n79# gnd
X0 vdd A Z w_692_n79# sky130_fd_pr__pfet_01v8 ad=1.5p pd=10.6u as=1.5p ps=10.6u w=5u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.504p pd=3.96u as=0.504p ps=3.96u w=1.68u l=0.15u
.ends

.subckt sky130_rom_krom_rom_bitline_inverter in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7
+ in_8 in_9 in_10 in_11 in_12 in_13 in_14 in_16 in_17 in_18 in_19 in_20 in_21 in_22
+ in_23 in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34 in_35 in_36
+ in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45 in_46 in_47 in_48 in_49 in_50
+ in_51 in_52 in_53 in_54 in_55 in_56 in_57 in_58 in_59 in_60 in_61 in_62 in_63 in_64
+ in_65 in_66 in_67 in_68 in_69 in_70 in_71 in_72 in_73 in_74 in_75 in_76 in_77 in_78
+ in_79 in_80 in_81 in_82 in_83 in_84 in_85 in_86 in_87 in_88 in_89 in_90 in_91 in_92
+ in_93 in_94 in_95 in_96 in_97 in_98 in_99 in_100 in_101 in_102 in_103 in_104 in_105
+ in_106 in_107 in_108 in_109 in_110 in_111 in_112 in_113 in_114 in_115 in_116 in_117
+ in_119 in_120 in_121 in_122 in_123 in_124 in_125 in_126 in_127 in_128 in_129 in_130
+ in_131 in_132 in_133 in_134 in_135 in_136 in_137 in_138 in_139 in_140 in_141 in_142
+ in_143 in_144 in_145 in_146 in_147 in_148 in_149 in_150 in_151 in_152 in_153 in_154
+ in_155 in_156 in_157 in_158 in_159 in_160 in_161 in_162 in_163 in_164 in_165 in_167
+ in_168 in_169 in_170 in_171 in_172 in_173 in_174 in_175 in_176 in_177 in_178 in_179
+ in_180 in_181 in_182 in_183 in_184 in_185 in_186 in_187 in_188 in_189 in_190 in_191
+ in_192 in_193 in_194 in_195 in_196 in_197 in_198 in_199 in_200 in_201 in_202 in_203
+ in_204 in_205 in_206 in_207 in_208 in_209 in_210 in_211 in_213 in_214 in_215 in_216
+ in_217 in_218 in_219 in_220 in_221 in_222 in_223 in_224 in_225 in_226 in_227 in_228
+ in_229 in_230 in_231 in_232 in_233 in_234 in_235 in_236 in_237 in_238 in_239 in_240
+ in_241 in_242 in_243 in_244 in_245 in_246 in_247 in_248 in_249 in_250 in_251 in_252
+ in_253 in_254 in_255 out_0 out_1 out_2 out_3 out_4 out_5 out_7 out_8 out_9 out_10
+ out_11 out_12 out_14 out_15 out_16 out_17 out_18 out_19 out_20 out_21 out_22 out_23
+ out_24 out_25 out_26 out_27 out_28 out_29 out_30 out_31 out_32 out_33 out_34 out_35
+ out_36 out_37 out_38 out_39 out_40 out_41 out_42 out_43 out_44 out_45 out_46 out_47
+ out_48 out_49 out_50 out_51 out_52 out_53 out_54 out_55 out_56 out_57 out_58 out_59
+ out_60 out_62 out_63 out_64 out_65 out_66 out_67 out_68 out_69 out_70 out_71 out_72
+ out_73 out_74 out_75 out_76 out_77 out_78 out_79 out_80 out_81 out_82 out_83 out_84
+ out_85 out_86 out_87 out_88 out_89 out_90 out_91 out_92 out_93 out_94 out_95 out_96
+ out_97 out_98 out_99 out_100 out_101 out_102 out_103 out_104 out_105 out_106 out_107
+ out_108 out_109 out_110 out_111 out_112 out_113 out_114 out_115 out_116 out_117
+ out_118 out_119 out_120 out_121 out_122 out_123 out_124 out_125 out_126 out_127
+ out_128 out_129 out_130 out_131 out_132 out_133 out_134 out_135 out_136 out_137
+ out_138 out_139 out_140 out_141 out_142 out_143 out_144 out_145 out_146 out_147
+ out_148 out_149 out_150 out_151 out_152 out_153 out_154 out_155 out_156 out_157
+ out_158 out_159 out_160 out_161 out_162 out_163 out_164 out_165 out_166 out_167
+ out_168 out_169 out_170 out_171 out_172 out_173 out_174 out_175 out_176 out_177
+ out_178 out_179 out_180 out_181 out_182 out_183 out_184 out_185 out_186 out_187
+ out_188 out_189 out_190 out_191 out_192 out_193 out_194 out_195 out_196 out_197
+ out_198 out_199 out_200 out_201 out_202 out_203 out_204 out_205 out_206 out_207
+ out_208 out_209 out_210 out_211 out_213 out_214 out_215 out_216 out_217 out_218
+ out_219 out_220 out_221 out_222 out_223 out_224 out_225 out_226 out_227 out_228
+ out_229 out_230 out_231 out_232 out_233 out_234 out_235 out_236 out_237 out_238
+ out_239 out_240 out_241 out_242 out_243 out_244 out_245 out_246 out_247 out_248
+ out_249 out_250 out_251 out_252 out_253 out_254 out_255 vdd in_15 gnd in_118 in_212
+ out_13 out_6 in_166 out_212 out_61 sky130_rom_krom_pinv_dec_3_9/w_692_n79#
Xsky130_rom_krom_pinv_dec_3_108 in_108 out_108 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_119 in_119 out_119 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_109 in_109 out_109 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_250 in_250 out_250 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_0 in_0 out_0 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_251 in_251 out_251 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_240 in_240 out_240 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_1 in_1 out_1 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_252 in_252 out_252 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_241 in_241 out_241 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_230 in_230 out_230 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_2 in_2 out_2 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_253 in_253 out_253 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_242 in_242 out_242 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_231 in_231 out_231 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_220 in_220 out_220 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_3 in_3 out_3 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_254 in_254 out_254 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_243 in_243 out_243 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_232 in_232 out_232 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_221 in_221 out_221 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_210 in_210 out_210 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_4 in_4 out_4 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_255 in_255 out_255 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_244 in_244 out_244 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_233 in_233 out_233 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_222 in_222 out_222 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_211 in_211 out_211 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_200 in_200 out_200 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_5 in_5 out_5 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_245 in_245 out_245 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_234 in_234 out_234 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_223 in_223 out_223 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_212 in_212 out_212 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_201 in_201 out_201 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_6 in_6 out_6 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_246 in_246 out_246 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_235 in_235 out_235 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_224 in_224 out_224 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_213 in_213 out_213 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_202 in_202 out_202 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_7 in_7 out_7 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_247 in_247 out_247 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_236 in_236 out_236 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_225 in_225 out_225 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_214 in_214 out_214 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_203 in_203 out_203 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_8 in_8 out_8 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_248 in_248 out_248 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_237 in_237 out_237 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_226 in_226 out_226 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_215 in_215 out_215 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_204 in_204 out_204 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_9 in_9 out_9 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_249 in_249 out_249 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_238 in_238 out_238 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_227 in_227 out_227 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_216 in_216 out_216 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_205 in_205 out_205 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_239 in_239 out_239 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_228 in_228 out_228 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_217 in_217 out_217 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_206 in_206 out_206 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_229 in_229 out_229 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_218 in_218 out_218 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_207 in_207 out_207 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_90 in_90 out_90 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_219 in_219 out_219 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_208 in_208 out_208 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_209 in_209 out_209 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_80 in_80 out_80 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_91 in_91 out_91 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_70 in_70 out_70 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_81 in_81 out_81 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_92 in_92 out_92 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_190 in_190 out_190 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_60 in_60 out_60 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_71 in_71 out_71 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_82 in_82 out_82 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_93 in_93 out_93 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_191 in_191 out_191 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_180 in_180 out_180 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_50 in_50 out_50 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_61 in_61 out_61 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_72 in_72 out_72 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_83 in_83 out_83 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_94 in_94 out_94 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_192 in_192 out_192 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_181 in_181 out_181 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_170 in_170 out_170 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_40 in_40 out_40 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_51 in_51 out_51 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_62 in_62 out_62 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_73 in_73 out_73 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_84 in_84 out_84 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_95 in_95 out_95 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_193 in_193 out_193 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_182 in_182 out_182 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_171 in_171 out_171 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_160 in_160 out_160 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_30 in_30 out_30 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_41 in_41 out_41 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_52 in_52 out_52 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_63 in_63 out_63 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_74 in_74 out_74 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_85 in_85 out_85 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_96 in_96 out_96 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_150 in_150 out_150 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_194 in_194 out_194 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_183 in_183 out_183 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_172 in_172 out_172 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_161 in_161 out_161 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_20 in_20 out_20 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_31 in_31 out_31 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_42 in_42 out_42 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_53 in_53 out_53 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_64 in_64 out_64 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_75 in_75 out_75 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_86 in_86 out_86 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_97 in_97 out_97 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_140 in_140 out_140 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_151 in_151 out_151 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_195 in_195 out_195 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_184 in_184 out_184 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_173 in_173 out_173 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_162 in_162 out_162 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_10 in_10 out_10 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_21 in_21 out_21 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_32 in_32 out_32 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_43 in_43 out_43 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_54 in_54 out_54 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_65 in_65 out_65 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_76 in_76 out_76 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_87 in_87 out_87 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_98 in_98 out_98 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_130 in_130 out_130 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_141 in_141 out_141 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_152 in_152 out_152 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_196 in_196 out_196 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_185 in_185 out_185 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_174 in_174 out_174 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_163 in_163 out_163 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_11 in_11 out_11 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_22 in_22 out_22 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_33 in_33 out_33 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_44 in_44 out_44 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_55 in_55 out_55 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_66 in_66 out_66 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_77 in_77 out_77 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_88 in_88 out_88 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_99 in_99 out_99 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_120 in_120 out_120 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_131 in_131 out_131 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_142 in_142 out_142 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_153 in_153 out_153 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_197 in_197 out_197 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_186 in_186 out_186 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_175 in_175 out_175 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_164 in_164 out_164 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_12 in_12 out_12 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_23 in_23 out_23 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_34 in_34 out_34 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_45 in_45 out_45 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_56 in_56 out_56 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_67 in_67 out_67 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_78 in_78 out_78 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_89 in_89 out_89 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_110 in_110 out_110 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_121 in_121 out_121 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_132 in_132 out_132 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_143 in_143 out_143 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_154 in_154 out_154 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_198 in_198 out_198 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_187 in_187 out_187 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_176 in_176 out_176 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_165 in_165 out_165 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_13 in_13 out_13 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_24 in_24 out_24 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_35 in_35 out_35 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_46 in_46 out_46 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_57 in_57 out_57 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_68 in_68 out_68 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_79 in_79 out_79 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_100 in_100 out_100 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_111 in_111 out_111 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_122 in_122 out_122 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_133 in_133 out_133 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_144 in_144 out_144 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_155 in_155 out_155 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_199 in_199 out_199 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_188 in_188 out_188 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_177 in_177 out_177 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_166 in_166 out_166 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_14 in_14 out_14 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_25 in_25 out_25 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_36 in_36 out_36 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_47 in_47 out_47 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_58 in_58 out_58 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_69 in_69 out_69 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_101 in_101 out_101 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_112 in_112 out_112 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_123 in_123 out_123 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_134 in_134 out_134 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_145 in_145 out_145 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_156 in_156 out_156 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_189 in_189 out_189 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_178 in_178 out_178 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_167 in_167 out_167 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_15 in_15 out_15 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_26 in_26 out_26 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_37 in_37 out_37 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_48 in_48 out_48 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_59 in_59 out_59 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_102 in_102 out_102 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_113 in_113 out_113 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_124 in_124 out_124 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_135 in_135 out_135 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_146 in_146 out_146 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_157 in_157 out_157 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_179 in_179 out_179 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_168 in_168 out_168 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_16 in_16 out_16 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_27 in_27 out_27 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_38 in_38 out_38 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_49 in_49 out_49 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_103 in_103 out_103 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_114 in_114 out_114 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_125 in_125 out_125 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_136 in_136 out_136 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_147 in_147 out_147 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_158 in_158 out_158 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_169 in_169 out_169 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_17 in_17 out_17 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_28 in_28 out_28 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_39 in_39 out_39 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_104 in_104 out_104 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_115 in_115 out_115 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_126 in_126 out_126 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_137 in_137 out_137 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_148 in_148 out_148 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_159 in_159 out_159 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_18 in_18 out_18 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_29 in_29 out_29 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_105 in_105 out_105 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_116 in_116 out_116 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_127 in_127 out_127 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_138 in_138 out_138 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_149 in_149 out_149 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_19 in_19 out_19 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_106 in_106 out_106 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_117 in_117 out_117 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_128 in_128 out_128 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_139 in_139 out_139 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_107 in_107 out_107 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_118 in_118 out_118 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
Xsky130_rom_krom_pinv_dec_3_129 in_129 out_129 vdd sky130_rom_krom_pinv_dec_3_9/w_692_n79#
+ gnd sky130_rom_krom_pinv_dec_3
.ends

.subckt sky130_rom_krom_pinv_dec_2 A Z vdd gnd w_504_n45#
X0 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.222p pd=2.08u as=0.222p ps=2.08u w=0.74u l=0.15u
X1 vdd A Z w_504_n45# sky130_fd_pr__pfet_01v8 ad=0.9p pd=6.6u as=0.9p ps=6.6u w=3u l=0.15u
.ends

.subckt sky130_rom_krom_rom_column_decode_wordline_buffer in_0 in_1 in_2 in_3 in_4
+ in_6 in_7 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd in_5
Xsky130_rom_krom_pinv_dec_2_0 in_7 out_7 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_1 in_6 out_6 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_2 in_5 out_5 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_3 in_4 out_4 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_4 in_3 out_3 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_5 in_2 out_2 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_7 in_0 out_0 vdd gnd vdd sky130_rom_krom_pinv_dec_2
Xsky130_rom_krom_pinv_dec_2_6 in_1 out_1 vdd gnd vdd sky130_rom_krom_pinv_dec_2
.ends

.subckt sky130_rom_krom_rom_column_decode A0 A1 A2 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6
+ wl_7 clk vdd_uq0 vdd_uq2 vdd_uq4 vdd precharge vdd_uq1 gnd
Xsky130_rom_krom_rom_row_decode_array_0 sky130_rom_krom_rom_row_decode_array_0/bl_0_0
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_1 sky130_rom_krom_rom_row_decode_array_0/bl_0_2
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_3 sky130_rom_krom_rom_row_decode_array_0/bl_0_4
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_5 sky130_rom_krom_rom_row_decode_array_0/bl_0_6
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_7 sky130_rom_krom_rom_row_decode_array_0/wl_0_1
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_2 sky130_rom_krom_rom_row_decode_array_0/wl_0_3
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_4 sky130_rom_krom_rom_row_decode_array_0/wl_0_5
+ gnd sky130_rom_krom_rom_row_decode_array_0/wl_0_0 vdd_uq0 precharge sky130_rom_krom_rom_row_decode_array
Xsky130_rom_krom_rom_address_control_array_0 A0 A1 A2 sky130_rom_krom_rom_row_decode_array_0/wl_0_5
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_3 sky130_rom_krom_rom_row_decode_array_0/wl_0_1
+ sky130_rom_krom_rom_row_decode_array_0/wl_0_4 sky130_rom_krom_rom_row_decode_array_0/wl_0_2
+ clk vdd_uq1 gnd vdd vdd_uq2 sky130_rom_krom_rom_row_decode_array_0/wl_0_0 sky130_rom_krom_rom_address_control_array
Xsky130_rom_krom_rom_column_decode_wordline_buffer_0 sky130_rom_krom_rom_row_decode_array_0/bl_0_0
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_1 sky130_rom_krom_rom_row_decode_array_0/bl_0_2
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_3 sky130_rom_krom_rom_row_decode_array_0/bl_0_4
+ sky130_rom_krom_rom_row_decode_array_0/bl_0_6 sky130_rom_krom_rom_row_decode_array_0/bl_0_7
+ wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 vdd_uq4 gnd sky130_rom_krom_rom_row_decode_array_0/bl_0_5
+ sky130_rom_krom_rom_column_decode_wordline_buffer
.ends

.subckt sky130_rom_krom clk0 cs0 addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5]
+ dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8]
+ dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17]
+ dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25]
+ dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31] vssd1
Xsky130_rom_krom_rom_row_decode_0 addr0[3] addr0[4] addr0[5] sky130_rom_krom_rom_row_decode_0/wl_0
+ sky130_rom_krom_rom_row_decode_0/wl_1 sky130_rom_krom_rom_row_decode_0/wl_2 sky130_rom_krom_rom_row_decode_0/wl_3
+ sky130_rom_krom_rom_row_decode_0/wl_4 sky130_rom_krom_rom_row_decode_0/wl_5 sky130_rom_krom_rom_row_decode_0/wl_6
+ sky130_rom_krom_rom_row_decode_0/wl_7 sky130_rom_krom_rom_row_decode_0/clk sky130_rom_krom_rom_row_decode_0/vdd_uq0
+ sky130_rom_krom_rom_row_decode_0/vdd_uq2 sky130_rom_krom_rom_row_decode_0/vdd_uq5
+ sky130_rom_krom_rom_row_decode_0/vdd_uq6 sky130_rom_krom_rom_row_decode_0/vdd sky130_rom_krom_rom_row_decode_0/vdd_uq1
+ sky130_rom_krom_rom_row_decode_0/clk gnd sky130_rom_krom_rom_row_decode
Xsky130_rom_krom_rom_output_buffer_0 sky130_rom_krom_rom_output_buffer_0/in_0 sky130_rom_krom_rom_output_buffer_0/in_1
+ sky130_rom_krom_rom_output_buffer_0/in_2 sky130_rom_krom_rom_output_buffer_0/in_3
+ sky130_rom_krom_rom_output_buffer_0/in_4 sky130_rom_krom_rom_output_buffer_0/in_5
+ sky130_rom_krom_rom_output_buffer_0/in_6 sky130_rom_krom_rom_output_buffer_0/in_7
+ sky130_rom_krom_rom_output_buffer_0/in_8 sky130_rom_krom_rom_output_buffer_0/in_9
+ sky130_rom_krom_rom_output_buffer_0/in_10 sky130_rom_krom_rom_output_buffer_0/in_11
+ sky130_rom_krom_rom_output_buffer_0/in_12 sky130_rom_krom_rom_output_buffer_0/in_13
+ sky130_rom_krom_rom_output_buffer_0/in_14 sky130_rom_krom_rom_output_buffer_0/in_15
+ sky130_rom_krom_rom_output_buffer_0/in_16 sky130_rom_krom_rom_output_buffer_0/in_17
+ sky130_rom_krom_rom_output_buffer_0/in_18 sky130_rom_krom_rom_output_buffer_0/in_19
+ sky130_rom_krom_rom_output_buffer_0/in_20 sky130_rom_krom_rom_output_buffer_0/in_21
+ sky130_rom_krom_rom_output_buffer_0/in_22 sky130_rom_krom_rom_output_buffer_0/in_23
+ sky130_rom_krom_rom_output_buffer_0/in_24 sky130_rom_krom_rom_output_buffer_0/in_25
+ sky130_rom_krom_rom_output_buffer_0/in_26 sky130_rom_krom_rom_output_buffer_0/in_27
+ sky130_rom_krom_rom_output_buffer_0/in_28 sky130_rom_krom_rom_output_buffer_0/in_29
+ sky130_rom_krom_rom_output_buffer_0/in_30 sky130_rom_krom_rom_output_buffer_0/in_31
+ dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8]
+ dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17]
+ dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25]
+ dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31] gnd sky130_rom_krom_rom_output_buffer_0/vdd
+ sky130_rom_krom_rom_output_buffer
Xsky130_rom_krom_rom_control_logic_0 clk0 cs0 sky130_rom_krom_rom_column_decode_0/clk
+ sky130_rom_krom_rom_row_decode_0/clk sky130_rom_krom_rom_control_logic_0/vdd gnd
+ sky130_rom_krom_rom_control_logic
Xsky130_rom_krom_rom_column_mux_array_0 sky130_rom_krom_rom_column_mux_array_0/bl_0
+ sky130_rom_krom_rom_column_mux_array_0/bl_1 sky130_rom_krom_rom_column_mux_array_0/bl_3
+ sky130_rom_krom_rom_column_mux_array_0/bl_4 sky130_rom_krom_rom_column_mux_array_0/bl_6
+ sky130_rom_krom_rom_column_mux_array_0/bl_8 sky130_rom_krom_rom_column_mux_array_0/bl_9
+ sky130_rom_krom_rom_column_mux_array_0/bl_11 sky130_rom_krom_rom_column_mux_array_0/bl_15
+ sky130_rom_krom_rom_column_mux_array_0/bl_16 sky130_rom_krom_rom_column_mux_array_0/bl_17
+ sky130_rom_krom_rom_column_mux_array_0/bl_18 sky130_rom_krom_rom_column_mux_array_0/bl_19
+ sky130_rom_krom_rom_column_mux_array_0/bl_26 sky130_rom_krom_rom_column_mux_array_0/bl_27
+ sky130_rom_krom_rom_column_mux_array_0/bl_28 sky130_rom_krom_rom_column_mux_array_0/bl_29
+ sky130_rom_krom_rom_column_mux_array_0/bl_30 sky130_rom_krom_rom_column_mux_array_0/bl_37
+ sky130_rom_krom_rom_column_mux_array_0/bl_38 sky130_rom_krom_rom_column_mux_array_0/bl_39
+ sky130_rom_krom_rom_column_mux_array_0/bl_41 sky130_rom_krom_rom_column_mux_array_0/bl_48
+ sky130_rom_krom_rom_column_mux_array_0/bl_49 sky130_rom_krom_rom_column_mux_array_0/bl_59
+ sky130_rom_krom_rom_column_mux_array_0/bl_71 sky130_rom_krom_rom_column_mux_array_0/bl_74
+ sky130_rom_krom_rom_column_mux_array_0/bl_76 sky130_rom_krom_rom_column_mux_array_0/bl_79
+ sky130_rom_krom_rom_column_mux_array_0/bl_82 sky130_rom_krom_rom_column_mux_array_0/bl_85
+ sky130_rom_krom_rom_column_mux_array_0/bl_87 sky130_rom_krom_rom_column_mux_array_0/bl_90
+ sky130_rom_krom_rom_column_mux_array_0/bl_93 sky130_rom_krom_rom_column_mux_array_0/bl_98
+ sky130_rom_krom_rom_column_mux_array_0/bl_100 sky130_rom_krom_rom_column_mux_array_0/bl_101
+ sky130_rom_krom_rom_column_mux_array_0/bl_102 sky130_rom_krom_rom_column_mux_array_0/bl_104
+ sky130_rom_krom_rom_column_mux_array_0/bl_105 sky130_rom_krom_rom_column_mux_array_0/bl_106
+ sky130_rom_krom_rom_column_mux_array_0/bl_107 sky130_rom_krom_rom_column_mux_array_0/bl_109
+ sky130_rom_krom_rom_column_mux_array_0/bl_110 sky130_rom_krom_rom_column_mux_array_0/bl_112
+ sky130_rom_krom_rom_column_mux_array_0/bl_113 sky130_rom_krom_rom_column_mux_array_0/bl_115
+ sky130_rom_krom_rom_column_mux_array_0/bl_117 sky130_rom_krom_rom_column_mux_array_0/bl_118
+ sky130_rom_krom_rom_column_mux_array_0/bl_120 sky130_rom_krom_rom_column_mux_array_0/bl_121
+ sky130_rom_krom_rom_column_mux_array_0/bl_123 sky130_rom_krom_rom_column_mux_array_0/bl_124
+ sky130_rom_krom_rom_column_mux_array_0/bl_126 sky130_rom_krom_rom_column_mux_array_0/bl_128
+ sky130_rom_krom_rom_column_mux_array_0/bl_129 sky130_rom_krom_rom_column_mux_array_0/bl_130
+ sky130_rom_krom_rom_column_mux_array_0/bl_131 sky130_rom_krom_rom_column_mux_array_0/bl_132
+ sky130_rom_krom_rom_column_mux_array_0/bl_134 sky130_rom_krom_rom_column_mux_array_0/bl_135
+ sky130_rom_krom_rom_column_mux_array_0/bl_136 sky130_rom_krom_rom_column_mux_array_0/bl_137
+ sky130_rom_krom_rom_column_mux_array_0/bl_139 sky130_rom_krom_rom_column_mux_array_0/bl_140
+ sky130_rom_krom_rom_column_mux_array_0/bl_141 sky130_rom_krom_rom_column_mux_array_0/bl_142
+ sky130_rom_krom_rom_column_mux_array_0/bl_143 sky130_rom_krom_rom_column_mux_array_0/bl_145
+ sky130_rom_krom_rom_column_mux_array_0/bl_147 sky130_rom_krom_rom_column_mux_array_0/bl_148
+ sky130_rom_krom_rom_column_mux_array_0/bl_150 sky130_rom_krom_rom_column_mux_array_0/bl_151
+ sky130_rom_krom_rom_column_mux_array_0/bl_153 sky130_rom_krom_rom_column_mux_array_0/bl_154
+ sky130_rom_krom_rom_column_mux_array_0/bl_157 sky130_rom_krom_rom_column_mux_array_0/bl_158
+ sky130_rom_krom_rom_column_mux_array_0/bl_160 sky130_rom_krom_rom_column_mux_array_0/bl_161
+ sky130_rom_krom_rom_column_mux_array_0/bl_163 sky130_rom_krom_rom_column_mux_array_0/bl_164
+ sky130_rom_krom_rom_column_mux_array_0/bl_166 sky130_rom_krom_rom_column_mux_array_0/bl_168
+ sky130_rom_krom_rom_column_mux_array_0/bl_169 sky130_rom_krom_rom_column_mux_array_0/bl_170
+ sky130_rom_krom_rom_column_mux_array_0/bl_171 sky130_rom_krom_rom_column_mux_array_0/bl_172
+ sky130_rom_krom_rom_column_mux_array_0/bl_174 sky130_rom_krom_rom_column_mux_array_0/bl_175
+ sky130_rom_krom_rom_column_mux_array_0/bl_176 sky130_rom_krom_rom_column_mux_array_0/bl_177
+ sky130_rom_krom_rom_column_mux_array_0/bl_179 sky130_rom_krom_rom_column_mux_array_0/bl_182
+ sky130_rom_krom_rom_column_mux_array_0/bl_183 sky130_rom_krom_rom_column_mux_array_0/bl_184
+ sky130_rom_krom_rom_column_mux_array_0/bl_185 sky130_rom_krom_rom_column_mux_array_0/bl_187
+ sky130_rom_krom_rom_column_mux_array_0/bl_188 sky130_rom_krom_rom_column_mux_array_0/bl_189
+ sky130_rom_krom_rom_column_mux_array_0/bl_192 sky130_rom_krom_rom_column_mux_array_0/bl_193
+ sky130_rom_krom_rom_column_mux_array_0/bl_194 sky130_rom_krom_rom_column_mux_array_0/bl_195
+ sky130_rom_krom_rom_column_mux_array_0/bl_196 sky130_rom_krom_rom_column_mux_array_0/bl_197
+ sky130_rom_krom_rom_column_mux_array_0/bl_198 sky130_rom_krom_rom_column_mux_array_0/bl_199
+ sky130_rom_krom_rom_column_mux_array_0/bl_200 sky130_rom_krom_rom_column_mux_array_0/bl_203
+ sky130_rom_krom_rom_column_mux_array_0/bl_208 sky130_rom_krom_rom_column_mux_array_0/bl_211
+ sky130_rom_krom_rom_column_mux_array_0/bl_214 sky130_rom_krom_rom_column_mux_array_0/bl_216
+ sky130_rom_krom_rom_column_mux_array_0/bl_219 sky130_rom_krom_rom_column_mux_array_0/bl_222
+ sky130_rom_krom_rom_column_mux_array_0/bl_225 sky130_rom_krom_rom_column_mux_array_0/bl_227
+ sky130_rom_krom_rom_column_mux_array_0/bl_230 sky130_rom_krom_rom_column_mux_array_0/bl_233
+ sky130_rom_krom_rom_column_mux_array_0/bl_238 sky130_rom_krom_rom_column_mux_array_0/bl_241
+ sky130_rom_krom_rom_column_mux_array_0/bl_244 sky130_rom_krom_rom_column_mux_array_0/bl_248
+ sky130_rom_krom_rom_column_mux_array_0/bl_251 sky130_rom_krom_rom_column_mux_array_0/bl_254
+ sky130_rom_krom_rom_column_decode_0/wl_4 sky130_rom_krom_rom_column_decode_0/wl_5
+ sky130_rom_krom_rom_output_buffer_0/in_0 sky130_rom_krom_rom_output_buffer_0/in_1
+ sky130_rom_krom_rom_output_buffer_0/in_2 sky130_rom_krom_rom_output_buffer_0/in_3
+ sky130_rom_krom_rom_output_buffer_0/in_4 sky130_rom_krom_rom_output_buffer_0/in_5
+ sky130_rom_krom_rom_output_buffer_0/in_6 sky130_rom_krom_rom_output_buffer_0/in_7
+ sky130_rom_krom_rom_output_buffer_0/in_8 sky130_rom_krom_rom_output_buffer_0/in_9
+ sky130_rom_krom_rom_output_buffer_0/in_10 sky130_rom_krom_rom_output_buffer_0/in_11
+ sky130_rom_krom_rom_output_buffer_0/in_12 sky130_rom_krom_rom_output_buffer_0/in_13
+ sky130_rom_krom_rom_output_buffer_0/in_14 sky130_rom_krom_rom_output_buffer_0/in_15
+ sky130_rom_krom_rom_output_buffer_0/in_16 sky130_rom_krom_rom_output_buffer_0/in_17
+ sky130_rom_krom_rom_output_buffer_0/in_18 sky130_rom_krom_rom_output_buffer_0/in_19
+ sky130_rom_krom_rom_output_buffer_0/in_20 sky130_rom_krom_rom_output_buffer_0/in_21
+ sky130_rom_krom_rom_output_buffer_0/in_22 sky130_rom_krom_rom_output_buffer_0/in_23
+ sky130_rom_krom_rom_output_buffer_0/in_24 sky130_rom_krom_rom_output_buffer_0/in_25
+ sky130_rom_krom_rom_output_buffer_0/in_26 sky130_rom_krom_rom_output_buffer_0/in_27
+ sky130_rom_krom_rom_output_buffer_0/in_28 sky130_rom_krom_rom_output_buffer_0/in_29
+ sky130_rom_krom_rom_output_buffer_0/in_30 sky130_rom_krom_rom_output_buffer_0/in_31
+ sky130_rom_krom_rom_column_mux_array_0/bl_14 sky130_rom_krom_rom_column_mux_array_0/bl_22
+ sky130_rom_krom_rom_column_mux_array_0/bl_25 sky130_rom_krom_rom_column_mux_array_0/bl_33
+ sky130_rom_krom_rom_column_mux_array_0/bl_46 sky130_rom_krom_rom_column_mux_array_0/bl_44
+ sky130_rom_krom_rom_column_mux_array_0/bl_52 sky130_rom_krom_rom_column_mux_array_0/bl_55
+ sky130_rom_krom_rom_column_mux_array_0/bl_58 sky130_rom_krom_rom_column_mux_array_0/bl_66
+ sky130_rom_krom_rom_column_mux_array_0/bl_61 sky130_rom_krom_rom_column_mux_array_0/bl_69
+ sky130_rom_krom_rom_column_mux_array_0/bl_64 sky130_rom_krom_rom_column_mux_array_0/bl_190
+ sky130_rom_krom_rom_column_mux_array_0/bl_77 sky130_rom_krom_rom_column_mux_array_0/bl_72
+ sky130_rom_krom_rom_column_mux_array_0/bl_80 sky130_rom_krom_rom_column_mux_array_0/bl_206
+ sky130_rom_krom_rom_column_mux_array_0/bl_75 sky130_rom_krom_rom_column_mux_array_0/bl_201
+ sky130_rom_krom_rom_column_mux_array_0/bl_88 sky130_rom_krom_rom_column_mux_array_0/bl_83
+ sky130_rom_krom_rom_column_mux_array_0/bl_209 sky130_rom_krom_rom_column_mux_array_0/bl_204
+ sky130_rom_krom_rom_column_mux_array_0/bl_96 sky130_rom_krom_rom_column_mux_array_0/bl_91
+ sky130_rom_krom_rom_column_mux_array_0/bl_217 sky130_rom_krom_rom_column_mux_array_0/bl_212
+ sky130_rom_krom_rom_column_mux_array_0/bl_99 sky130_rom_krom_rom_column_mux_array_0/bl_94
+ sky130_rom_krom_rom_column_mux_array_0/bl_220 sky130_rom_krom_rom_column_mux_array_0/bl_215
+ sky130_rom_krom_rom_column_mux_array_0/bl_12 sky130_rom_krom_rom_column_mux_array_0/bl_246
+ sky130_rom_krom_rom_column_mux_array_0/bl_228 sky130_rom_krom_rom_column_mux_array_0/bl_223
+ sky130_rom_krom_rom_column_mux_array_0/bl_20 sky130_rom_krom_rom_column_mux_array_0/bl_236
+ sky130_rom_krom_rom_column_mux_array_0/bl_231 sky130_rom_krom_rom_column_mux_array_0/bl_249
+ sky130_rom_krom_rom_column_mux_array_0/bl_23 sky130_rom_krom_rom_column_mux_array_0/bl_239
+ sky130_rom_krom_rom_column_mux_array_0/bl_36 sky130_rom_krom_rom_column_mux_array_0/bl_252
+ sky130_rom_krom_rom_column_mux_array_0/bl_234 sky130_rom_krom_rom_column_mux_array_0/bl_31
+ sky130_rom_krom_rom_column_mux_array_0/bl_242 sky130_rom_krom_rom_column_mux_array_0/bl_255
+ sky130_rom_krom_rom_column_mux_array_0/bl_34 sky130_rom_krom_rom_column_mux_array_0/bl_245
+ sky130_rom_krom_rom_column_mux_array_0/bl_47 sky130_rom_krom_rom_column_mux_array_0/bl_42
+ sky130_rom_krom_rom_column_mux_array_0/bl_50 sky130_rom_krom_rom_column_mux_array_0/bl_45
+ sky130_rom_krom_rom_column_mux_array_0/bl_53 sky130_rom_krom_rom_column_mux_array_0/bl_56
+ sky130_rom_krom_rom_column_mux_array_0/bl_180 sky130_rom_krom_rom_column_mux_array_0/bl_67
+ sky130_rom_krom_rom_column_mux_array_0/bl_62 sky130_rom_krom_rom_column_mux_array_0/bl_70
+ sky130_rom_krom_rom_column_mux_array_0/bl_65 sky130_rom_krom_rom_column_mux_array_0/bl_191
+ sky130_rom_krom_rom_column_mux_array_0/bl_78 sky130_rom_krom_rom_column_mux_array_0/bl_73
+ sky130_rom_krom_rom_column_mux_array_0/bl_86 sky130_rom_krom_rom_column_mux_array_0/bl_81
+ sky130_rom_krom_rom_column_mux_array_0/bl_207 sky130_rom_krom_rom_column_mux_array_0/bl_202
+ sky130_rom_krom_rom_column_mux_array_0/bl_89 sky130_rom_krom_rom_column_mux_array_0/bl_84
+ sky130_rom_krom_rom_column_mux_array_0/bl_210 sky130_rom_krom_rom_column_mux_array_0/bl_7
+ sky130_rom_krom_rom_column_mux_array_0/bl_205 sky130_rom_krom_rom_column_mux_array_0/bl_97
+ sky130_rom_krom_rom_column_mux_array_0/bl_92 sky130_rom_krom_rom_column_mux_array_0/bl_2
+ sky130_rom_krom_rom_column_mux_array_0/bl_218 sky130_rom_krom_rom_column_mux_array_0/bl_213
+ sky130_rom_krom_rom_column_mux_array_0/bl_10 sky130_rom_krom_rom_column_mux_array_0/bl_95
+ sky130_rom_krom_rom_column_mux_array_0/bl_5 sky130_rom_krom_rom_column_mux_array_0/bl_226
+ sky130_rom_krom_rom_column_mux_array_0/bl_221 sky130_rom_krom_rom_column_mux_array_0/bl_108
+ sky130_rom_krom_rom_column_mux_array_0/bl_103 sky130_rom_krom_rom_column_mux_array_0/bl_13
+ sky130_rom_krom_rom_column_mux_array_0/bl_229 sky130_rom_krom_rom_column_mux_array_0/bl_247
+ sky130_rom_krom_rom_column_mux_array_0/bl_224 sky130_rom_krom_rom_column_mux_array_0/bl_116
+ sky130_rom_krom_rom_column_mux_array_0/bl_111 sky130_rom_krom_rom_column_mux_array_0/bl_21
+ sky130_rom_krom_rom_column_mux_array_0/bl_237 sky130_rom_krom_rom_column_mux_array_0/bl_250
+ sky130_rom_krom_rom_column_mux_array_0/bl_232 sky130_rom_krom_rom_column_mux_array_0/bl_119
+ sky130_rom_krom_rom_column_mux_array_0/bl_114 sky130_rom_krom_rom_column_mux_array_0/bl_24
+ sky130_rom_krom_rom_column_mux_array_0/bl_240 sky130_rom_krom_rom_column_mux_array_0/bl_235
+ sky130_rom_krom_rom_column_mux_array_0/bl_127 sky130_rom_krom_rom_column_mux_array_0/bl_253
+ sky130_rom_krom_rom_column_mux_array_0/bl_32 sky130_rom_krom_rom_column_mux_array_0/bl_122
+ sky130_rom_krom_rom_column_mux_array_0/bl_243 sky130_rom_krom_rom_column_mux_array_0/bl_40
+ sky130_rom_krom_rom_column_mux_array_0/bl_125 sky130_rom_krom_rom_column_mux_array_0/bl_35
+ sky130_rom_krom_rom_column_mux_array_0/bl_138 sky130_rom_krom_rom_column_mux_array_0/bl_133
+ sky130_rom_krom_rom_column_mux_array_0/bl_43 sky130_rom_krom_rom_column_mux_array_0/bl_146
+ sky130_rom_krom_rom_column_mux_array_0/bl_51 sky130_rom_krom_rom_column_mux_array_0/bl_149
+ sky130_rom_krom_rom_column_mux_array_0/bl_144 sky130_rom_krom_rom_column_mux_array_0/bl_54
+ sky130_rom_krom_rom_column_mux_array_0/bl_152 sky130_rom_krom_rom_column_mux_array_0/bl_156
+ sky130_rom_krom_rom_column_mux_array_0/bl_155 sky130_rom_krom_rom_column_mux_array_0/bl_159
+ sky130_rom_krom_rom_column_mux_array_0/bl_167 sky130_rom_krom_rom_column_mux_array_0/bl_162
+ sky130_rom_krom_rom_column_decode_0/wl_0 sky130_rom_krom_rom_column_decode_0/wl_7
+ sky130_rom_krom_rom_column_decode_0/wl_6 sky130_rom_krom_rom_column_mux_array_0/bl_57
+ sky130_rom_krom_rom_column_mux_array_0/bl_165 sky130_rom_krom_rom_column_decode_0/wl_1
+ sky130_rom_krom_rom_column_mux_array_0/bl_178 sky130_rom_krom_rom_column_mux_array_0/bl_173
+ gnd sky130_rom_krom_rom_column_mux_array_0/bl_60 sky130_rom_krom_rom_column_mux_array_0/bl_186
+ sky130_rom_krom_rom_column_mux_array_0/bl_181 sky130_rom_krom_rom_column_mux_array_0/bl_68
+ sky130_rom_krom_rom_column_decode_0/wl_3 sky130_rom_krom_rom_column_mux_array_0/bl_63
+ sky130_rom_krom_rom_column_decode_0/wl_2 sky130_rom_krom_rom_column_mux_array
Xsky130_rom_krom_rom_base_array_0 sky130_rom_krom_rom_base_array_0/bl_0_0 sky130_rom_krom_rom_base_array_0/bl_0_1
+ sky130_rom_krom_rom_base_array_0/bl_0_2 sky130_rom_krom_rom_base_array_0/bl_0_3
+ sky130_rom_krom_rom_base_array_0/bl_0_4 sky130_rom_krom_rom_base_array_0/bl_0_5
+ sky130_rom_krom_rom_base_array_0/bl_0_6 sky130_rom_krom_rom_base_array_0/bl_0_7
+ sky130_rom_krom_rom_base_array_0/bl_0_8 sky130_rom_krom_rom_base_array_0/bl_0_9
+ sky130_rom_krom_rom_base_array_0/bl_0_10 sky130_rom_krom_rom_base_array_0/bl_0_11
+ sky130_rom_krom_rom_base_array_0/bl_0_12 sky130_rom_krom_rom_base_array_0/bl_0_13
+ sky130_rom_krom_rom_base_array_0/bl_0_14 sky130_rom_krom_rom_base_array_0/bl_0_16
+ sky130_rom_krom_rom_base_array_0/bl_0_17 sky130_rom_krom_rom_base_array_0/bl_0_18
+ sky130_rom_krom_rom_base_array_0/bl_0_19 sky130_rom_krom_rom_base_array_0/bl_0_20
+ sky130_rom_krom_rom_base_array_0/bl_0_21 sky130_rom_krom_rom_base_array_0/bl_0_22
+ sky130_rom_krom_rom_base_array_0/bl_0_23 sky130_rom_krom_rom_base_array_0/bl_0_24
+ sky130_rom_krom_rom_base_array_0/bl_0_25 sky130_rom_krom_rom_base_array_0/bl_0_26
+ sky130_rom_krom_rom_base_array_0/bl_0_27 sky130_rom_krom_rom_base_array_0/bl_0_28
+ sky130_rom_krom_rom_base_array_0/bl_0_29 sky130_rom_krom_rom_base_array_0/bl_0_30
+ sky130_rom_krom_rom_base_array_0/bl_0_31 sky130_rom_krom_rom_base_array_0/bl_0_32
+ sky130_rom_krom_rom_base_array_0/bl_0_33 sky130_rom_krom_rom_base_array_0/bl_0_34
+ sky130_rom_krom_rom_base_array_0/bl_0_35 sky130_rom_krom_rom_base_array_0/bl_0_36
+ sky130_rom_krom_rom_base_array_0/bl_0_37 sky130_rom_krom_rom_base_array_0/bl_0_38
+ sky130_rom_krom_rom_base_array_0/bl_0_39 sky130_rom_krom_rom_base_array_0/bl_0_40
+ sky130_rom_krom_rom_base_array_0/bl_0_41 sky130_rom_krom_rom_base_array_0/bl_0_42
+ sky130_rom_krom_rom_base_array_0/bl_0_43 sky130_rom_krom_rom_base_array_0/bl_0_44
+ sky130_rom_krom_rom_base_array_0/bl_0_45 sky130_rom_krom_rom_base_array_0/bl_0_46
+ sky130_rom_krom_rom_base_array_0/bl_0_47 sky130_rom_krom_rom_base_array_0/bl_0_48
+ sky130_rom_krom_rom_base_array_0/bl_0_49 sky130_rom_krom_rom_base_array_0/bl_0_50
+ sky130_rom_krom_rom_base_array_0/bl_0_51 sky130_rom_krom_rom_base_array_0/bl_0_52
+ sky130_rom_krom_rom_base_array_0/bl_0_53 sky130_rom_krom_rom_base_array_0/bl_0_54
+ sky130_rom_krom_rom_base_array_0/bl_0_55 sky130_rom_krom_rom_base_array_0/bl_0_56
+ sky130_rom_krom_rom_base_array_0/bl_0_57 sky130_rom_krom_rom_base_array_0/bl_0_58
+ sky130_rom_krom_rom_base_array_0/bl_0_59 sky130_rom_krom_rom_base_array_0/bl_0_60
+ sky130_rom_krom_rom_base_array_0/bl_0_61 sky130_rom_krom_rom_base_array_0/bl_0_62
+ sky130_rom_krom_rom_base_array_0/bl_0_63 sky130_rom_krom_rom_base_array_0/bl_0_64
+ sky130_rom_krom_rom_base_array_0/bl_0_65 sky130_rom_krom_rom_base_array_0/bl_0_66
+ sky130_rom_krom_rom_base_array_0/bl_0_67 sky130_rom_krom_rom_base_array_0/bl_0_68
+ sky130_rom_krom_rom_base_array_0/bl_0_69 sky130_rom_krom_rom_base_array_0/bl_0_70
+ sky130_rom_krom_rom_base_array_0/bl_0_71 sky130_rom_krom_rom_base_array_0/bl_0_72
+ sky130_rom_krom_rom_base_array_0/bl_0_73 sky130_rom_krom_rom_base_array_0/bl_0_74
+ sky130_rom_krom_rom_base_array_0/bl_0_75 sky130_rom_krom_rom_base_array_0/bl_0_76
+ sky130_rom_krom_rom_base_array_0/bl_0_77 sky130_rom_krom_rom_base_array_0/bl_0_78
+ sky130_rom_krom_rom_base_array_0/bl_0_79 sky130_rom_krom_rom_base_array_0/bl_0_80
+ sky130_rom_krom_rom_base_array_0/bl_0_81 sky130_rom_krom_rom_base_array_0/bl_0_82
+ sky130_rom_krom_rom_base_array_0/bl_0_83 sky130_rom_krom_rom_base_array_0/bl_0_84
+ sky130_rom_krom_rom_base_array_0/bl_0_85 sky130_rom_krom_rom_base_array_0/bl_0_86
+ sky130_rom_krom_rom_base_array_0/bl_0_87 sky130_rom_krom_rom_base_array_0/bl_0_88
+ sky130_rom_krom_rom_base_array_0/bl_0_89 sky130_rom_krom_rom_base_array_0/bl_0_90
+ sky130_rom_krom_rom_base_array_0/bl_0_91 sky130_rom_krom_rom_base_array_0/bl_0_92
+ sky130_rom_krom_rom_base_array_0/bl_0_93 sky130_rom_krom_rom_base_array_0/bl_0_94
+ sky130_rom_krom_rom_base_array_0/bl_0_95 sky130_rom_krom_rom_base_array_0/bl_0_96
+ sky130_rom_krom_rom_base_array_0/bl_0_97 sky130_rom_krom_rom_base_array_0/bl_0_98
+ sky130_rom_krom_rom_base_array_0/bl_0_99 sky130_rom_krom_rom_base_array_0/bl_0_100
+ sky130_rom_krom_rom_base_array_0/bl_0_101 sky130_rom_krom_rom_base_array_0/bl_0_102
+ sky130_rom_krom_rom_base_array_0/bl_0_103 sky130_rom_krom_rom_base_array_0/bl_0_104
+ sky130_rom_krom_rom_base_array_0/bl_0_105 sky130_rom_krom_rom_base_array_0/bl_0_106
+ sky130_rom_krom_rom_base_array_0/bl_0_107 sky130_rom_krom_rom_base_array_0/bl_0_108
+ sky130_rom_krom_rom_base_array_0/bl_0_109 sky130_rom_krom_rom_base_array_0/bl_0_110
+ sky130_rom_krom_rom_base_array_0/bl_0_111 sky130_rom_krom_rom_base_array_0/bl_0_112
+ sky130_rom_krom_rom_base_array_0/bl_0_113 sky130_rom_krom_rom_base_array_0/bl_0_114
+ sky130_rom_krom_rom_base_array_0/bl_0_115 sky130_rom_krom_rom_base_array_0/bl_0_116
+ sky130_rom_krom_rom_base_array_0/bl_0_117 sky130_rom_krom_rom_base_array_0/bl_0_118
+ sky130_rom_krom_rom_base_array_0/bl_0_119 sky130_rom_krom_rom_base_array_0/bl_0_120
+ sky130_rom_krom_rom_base_array_0/bl_0_121 sky130_rom_krom_rom_base_array_0/bl_0_122
+ sky130_rom_krom_rom_base_array_0/bl_0_123 sky130_rom_krom_rom_base_array_0/bl_0_124
+ sky130_rom_krom_rom_base_array_0/bl_0_125 sky130_rom_krom_rom_base_array_0/bl_0_126
+ sky130_rom_krom_rom_base_array_0/bl_0_127 sky130_rom_krom_rom_base_array_0/bl_0_128
+ sky130_rom_krom_rom_base_array_0/bl_0_129 sky130_rom_krom_rom_base_array_0/bl_0_130
+ sky130_rom_krom_rom_base_array_0/bl_0_131 sky130_rom_krom_rom_base_array_0/bl_0_132
+ sky130_rom_krom_rom_base_array_0/bl_0_133 sky130_rom_krom_rom_base_array_0/bl_0_134
+ sky130_rom_krom_rom_base_array_0/bl_0_135 sky130_rom_krom_rom_base_array_0/bl_0_136
+ sky130_rom_krom_rom_base_array_0/bl_0_137 sky130_rom_krom_rom_base_array_0/bl_0_138
+ sky130_rom_krom_rom_base_array_0/bl_0_139 sky130_rom_krom_rom_base_array_0/bl_0_140
+ sky130_rom_krom_rom_base_array_0/bl_0_141 sky130_rom_krom_rom_base_array_0/bl_0_142
+ sky130_rom_krom_rom_base_array_0/bl_0_143 sky130_rom_krom_rom_base_array_0/bl_0_144
+ sky130_rom_krom_rom_base_array_0/bl_0_145 sky130_rom_krom_rom_base_array_0/bl_0_146
+ sky130_rom_krom_rom_base_array_0/bl_0_147 sky130_rom_krom_rom_base_array_0/bl_0_148
+ sky130_rom_krom_rom_base_array_0/bl_0_149 sky130_rom_krom_rom_base_array_0/bl_0_150
+ sky130_rom_krom_rom_base_array_0/bl_0_151 sky130_rom_krom_rom_base_array_0/bl_0_152
+ sky130_rom_krom_rom_base_array_0/bl_0_153 sky130_rom_krom_rom_base_array_0/bl_0_154
+ sky130_rom_krom_rom_base_array_0/bl_0_155 sky130_rom_krom_rom_base_array_0/bl_0_156
+ sky130_rom_krom_rom_base_array_0/bl_0_157 sky130_rom_krom_rom_base_array_0/bl_0_158
+ sky130_rom_krom_rom_base_array_0/bl_0_159 sky130_rom_krom_rom_base_array_0/bl_0_160
+ sky130_rom_krom_rom_base_array_0/bl_0_161 sky130_rom_krom_rom_base_array_0/bl_0_162
+ sky130_rom_krom_rom_base_array_0/bl_0_163 sky130_rom_krom_rom_base_array_0/bl_0_164
+ sky130_rom_krom_rom_base_array_0/bl_0_165 sky130_rom_krom_rom_base_array_0/bl_0_166
+ sky130_rom_krom_rom_base_array_0/bl_0_167 sky130_rom_krom_rom_base_array_0/bl_0_168
+ sky130_rom_krom_rom_base_array_0/bl_0_169 sky130_rom_krom_rom_base_array_0/bl_0_170
+ sky130_rom_krom_rom_base_array_0/bl_0_171 sky130_rom_krom_rom_base_array_0/bl_0_172
+ sky130_rom_krom_rom_base_array_0/bl_0_173 sky130_rom_krom_rom_base_array_0/bl_0_174
+ sky130_rom_krom_rom_base_array_0/bl_0_175 sky130_rom_krom_rom_base_array_0/bl_0_176
+ sky130_rom_krom_rom_base_array_0/bl_0_177 sky130_rom_krom_rom_base_array_0/bl_0_178
+ sky130_rom_krom_rom_base_array_0/bl_0_179 sky130_rom_krom_rom_base_array_0/bl_0_180
+ sky130_rom_krom_rom_base_array_0/bl_0_181 sky130_rom_krom_rom_base_array_0/bl_0_182
+ sky130_rom_krom_rom_base_array_0/bl_0_183 sky130_rom_krom_rom_base_array_0/bl_0_184
+ sky130_rom_krom_rom_base_array_0/bl_0_185 sky130_rom_krom_rom_base_array_0/bl_0_186
+ sky130_rom_krom_rom_base_array_0/bl_0_187 sky130_rom_krom_rom_base_array_0/bl_0_188
+ sky130_rom_krom_rom_base_array_0/bl_0_189 sky130_rom_krom_rom_base_array_0/bl_0_190
+ sky130_rom_krom_rom_base_array_0/bl_0_191 sky130_rom_krom_rom_base_array_0/bl_0_192
+ sky130_rom_krom_rom_base_array_0/bl_0_193 sky130_rom_krom_rom_base_array_0/bl_0_194
+ sky130_rom_krom_rom_base_array_0/bl_0_195 sky130_rom_krom_rom_base_array_0/bl_0_196
+ sky130_rom_krom_rom_base_array_0/bl_0_197 sky130_rom_krom_rom_base_array_0/bl_0_198
+ sky130_rom_krom_rom_base_array_0/bl_0_199 sky130_rom_krom_rom_base_array_0/bl_0_200
+ sky130_rom_krom_rom_base_array_0/bl_0_201 sky130_rom_krom_rom_base_array_0/bl_0_202
+ sky130_rom_krom_rom_base_array_0/bl_0_203 sky130_rom_krom_rom_base_array_0/bl_0_204
+ sky130_rom_krom_rom_base_array_0/bl_0_205 sky130_rom_krom_rom_base_array_0/bl_0_206
+ sky130_rom_krom_rom_base_array_0/bl_0_207 sky130_rom_krom_rom_base_array_0/bl_0_208
+ sky130_rom_krom_rom_base_array_0/bl_0_209 sky130_rom_krom_rom_base_array_0/bl_0_210
+ sky130_rom_krom_rom_base_array_0/bl_0_211 sky130_rom_krom_rom_base_array_0/bl_0_212
+ sky130_rom_krom_rom_base_array_0/bl_0_213 sky130_rom_krom_rom_base_array_0/bl_0_214
+ sky130_rom_krom_rom_base_array_0/bl_0_215 sky130_rom_krom_rom_base_array_0/bl_0_216
+ sky130_rom_krom_rom_base_array_0/bl_0_217 sky130_rom_krom_rom_base_array_0/bl_0_218
+ sky130_rom_krom_rom_base_array_0/bl_0_219 sky130_rom_krom_rom_base_array_0/bl_0_220
+ sky130_rom_krom_rom_base_array_0/bl_0_221 sky130_rom_krom_rom_base_array_0/bl_0_222
+ sky130_rom_krom_rom_base_array_0/bl_0_223 sky130_rom_krom_rom_base_array_0/bl_0_224
+ sky130_rom_krom_rom_base_array_0/bl_0_225 sky130_rom_krom_rom_base_array_0/bl_0_226
+ sky130_rom_krom_rom_base_array_0/bl_0_227 sky130_rom_krom_rom_base_array_0/bl_0_228
+ sky130_rom_krom_rom_base_array_0/bl_0_229 sky130_rom_krom_rom_base_array_0/bl_0_230
+ sky130_rom_krom_rom_base_array_0/bl_0_231 sky130_rom_krom_rom_base_array_0/bl_0_232
+ sky130_rom_krom_rom_base_array_0/bl_0_233 sky130_rom_krom_rom_base_array_0/bl_0_234
+ sky130_rom_krom_rom_base_array_0/bl_0_235 sky130_rom_krom_rom_base_array_0/bl_0_236
+ sky130_rom_krom_rom_base_array_0/bl_0_237 sky130_rom_krom_rom_base_array_0/bl_0_238
+ sky130_rom_krom_rom_base_array_0/bl_0_239 sky130_rom_krom_rom_base_array_0/bl_0_240
+ sky130_rom_krom_rom_base_array_0/bl_0_241 sky130_rom_krom_rom_base_array_0/bl_0_242
+ sky130_rom_krom_rom_base_array_0/bl_0_243 sky130_rom_krom_rom_base_array_0/bl_0_244
+ sky130_rom_krom_rom_base_array_0/bl_0_245 sky130_rom_krom_rom_base_array_0/bl_0_246
+ sky130_rom_krom_rom_base_array_0/bl_0_247 sky130_rom_krom_rom_base_array_0/bl_0_248
+ sky130_rom_krom_rom_base_array_0/bl_0_249 sky130_rom_krom_rom_base_array_0/bl_0_250
+ sky130_rom_krom_rom_base_array_0/bl_0_251 sky130_rom_krom_rom_base_array_0/bl_0_252
+ sky130_rom_krom_rom_base_array_0/bl_0_253 sky130_rom_krom_rom_base_array_0/bl_0_254
+ sky130_rom_krom_rom_base_array_0/bl_0_255 sky130_rom_krom_rom_row_decode_0/wl_1
+ sky130_rom_krom_rom_row_decode_0/wl_2 sky130_rom_krom_rom_row_decode_0/wl_4 sky130_rom_krom_rom_row_decode_0/wl_5
+ sky130_rom_krom_rom_row_decode_0/wl_6 sky130_rom_krom_rom_row_decode_0/wl_7 gnd
+ sky130_rom_krom_rom_base_array_0/gnd_uq0 sky130_rom_krom_rom_base_array_0/bl_0_15
+ sky130_rom_krom_rom_row_decode_0/wl_0 sky130_rom_krom_rom_column_decode_0/clk sky130_rom_krom_rom_row_decode_0/wl_3
+ sky130_rom_krom_rom_base_array_0/vdd sky130_rom_krom_rom_base_array
Xsky130_rom_krom_rom_bitline_inverter_0 sky130_rom_krom_rom_base_array_0/bl_0_0 sky130_rom_krom_rom_base_array_0/bl_0_1
+ sky130_rom_krom_rom_base_array_0/bl_0_2 sky130_rom_krom_rom_base_array_0/bl_0_3
+ sky130_rom_krom_rom_base_array_0/bl_0_4 sky130_rom_krom_rom_base_array_0/bl_0_5
+ sky130_rom_krom_rom_base_array_0/bl_0_6 sky130_rom_krom_rom_base_array_0/bl_0_7
+ sky130_rom_krom_rom_base_array_0/bl_0_8 sky130_rom_krom_rom_base_array_0/bl_0_9
+ sky130_rom_krom_rom_base_array_0/bl_0_10 sky130_rom_krom_rom_base_array_0/bl_0_11
+ sky130_rom_krom_rom_base_array_0/bl_0_12 sky130_rom_krom_rom_base_array_0/bl_0_13
+ sky130_rom_krom_rom_base_array_0/bl_0_14 sky130_rom_krom_rom_base_array_0/bl_0_16
+ sky130_rom_krom_rom_base_array_0/bl_0_17 sky130_rom_krom_rom_base_array_0/bl_0_18
+ sky130_rom_krom_rom_base_array_0/bl_0_19 sky130_rom_krom_rom_base_array_0/bl_0_20
+ sky130_rom_krom_rom_base_array_0/bl_0_21 sky130_rom_krom_rom_base_array_0/bl_0_22
+ sky130_rom_krom_rom_base_array_0/bl_0_23 sky130_rom_krom_rom_base_array_0/bl_0_24
+ sky130_rom_krom_rom_base_array_0/bl_0_25 sky130_rom_krom_rom_base_array_0/bl_0_26
+ sky130_rom_krom_rom_base_array_0/bl_0_27 sky130_rom_krom_rom_base_array_0/bl_0_28
+ sky130_rom_krom_rom_base_array_0/bl_0_29 sky130_rom_krom_rom_base_array_0/bl_0_30
+ sky130_rom_krom_rom_base_array_0/bl_0_31 sky130_rom_krom_rom_base_array_0/bl_0_32
+ sky130_rom_krom_rom_base_array_0/bl_0_33 sky130_rom_krom_rom_base_array_0/bl_0_34
+ sky130_rom_krom_rom_base_array_0/bl_0_35 sky130_rom_krom_rom_base_array_0/bl_0_36
+ sky130_rom_krom_rom_base_array_0/bl_0_37 sky130_rom_krom_rom_base_array_0/bl_0_38
+ sky130_rom_krom_rom_base_array_0/bl_0_39 sky130_rom_krom_rom_base_array_0/bl_0_40
+ sky130_rom_krom_rom_base_array_0/bl_0_41 sky130_rom_krom_rom_base_array_0/bl_0_42
+ sky130_rom_krom_rom_base_array_0/bl_0_43 sky130_rom_krom_rom_base_array_0/bl_0_44
+ sky130_rom_krom_rom_base_array_0/bl_0_45 sky130_rom_krom_rom_base_array_0/bl_0_46
+ sky130_rom_krom_rom_base_array_0/bl_0_47 sky130_rom_krom_rom_base_array_0/bl_0_48
+ sky130_rom_krom_rom_base_array_0/bl_0_49 sky130_rom_krom_rom_base_array_0/bl_0_50
+ sky130_rom_krom_rom_base_array_0/bl_0_51 sky130_rom_krom_rom_base_array_0/bl_0_52
+ sky130_rom_krom_rom_base_array_0/bl_0_53 sky130_rom_krom_rom_base_array_0/bl_0_54
+ sky130_rom_krom_rom_base_array_0/bl_0_55 sky130_rom_krom_rom_base_array_0/bl_0_56
+ sky130_rom_krom_rom_base_array_0/bl_0_57 sky130_rom_krom_rom_base_array_0/bl_0_58
+ sky130_rom_krom_rom_base_array_0/bl_0_59 sky130_rom_krom_rom_base_array_0/bl_0_60
+ sky130_rom_krom_rom_base_array_0/bl_0_61 sky130_rom_krom_rom_base_array_0/bl_0_62
+ sky130_rom_krom_rom_base_array_0/bl_0_63 sky130_rom_krom_rom_base_array_0/bl_0_64
+ sky130_rom_krom_rom_base_array_0/bl_0_65 sky130_rom_krom_rom_base_array_0/bl_0_66
+ sky130_rom_krom_rom_base_array_0/bl_0_67 sky130_rom_krom_rom_base_array_0/bl_0_68
+ sky130_rom_krom_rom_base_array_0/bl_0_69 sky130_rom_krom_rom_base_array_0/bl_0_70
+ sky130_rom_krom_rom_base_array_0/bl_0_71 sky130_rom_krom_rom_base_array_0/bl_0_72
+ sky130_rom_krom_rom_base_array_0/bl_0_73 sky130_rom_krom_rom_base_array_0/bl_0_74
+ sky130_rom_krom_rom_base_array_0/bl_0_75 sky130_rom_krom_rom_base_array_0/bl_0_76
+ sky130_rom_krom_rom_base_array_0/bl_0_77 sky130_rom_krom_rom_base_array_0/bl_0_78
+ sky130_rom_krom_rom_base_array_0/bl_0_79 sky130_rom_krom_rom_base_array_0/bl_0_80
+ sky130_rom_krom_rom_base_array_0/bl_0_81 sky130_rom_krom_rom_base_array_0/bl_0_82
+ sky130_rom_krom_rom_base_array_0/bl_0_83 sky130_rom_krom_rom_base_array_0/bl_0_84
+ sky130_rom_krom_rom_base_array_0/bl_0_85 sky130_rom_krom_rom_base_array_0/bl_0_86
+ sky130_rom_krom_rom_base_array_0/bl_0_87 sky130_rom_krom_rom_base_array_0/bl_0_88
+ sky130_rom_krom_rom_base_array_0/bl_0_89 sky130_rom_krom_rom_base_array_0/bl_0_90
+ sky130_rom_krom_rom_base_array_0/bl_0_91 sky130_rom_krom_rom_base_array_0/bl_0_92
+ sky130_rom_krom_rom_base_array_0/bl_0_93 sky130_rom_krom_rom_base_array_0/bl_0_94
+ sky130_rom_krom_rom_base_array_0/bl_0_95 sky130_rom_krom_rom_base_array_0/bl_0_96
+ sky130_rom_krom_rom_base_array_0/bl_0_97 sky130_rom_krom_rom_base_array_0/bl_0_98
+ sky130_rom_krom_rom_base_array_0/bl_0_99 sky130_rom_krom_rom_base_array_0/bl_0_100
+ sky130_rom_krom_rom_base_array_0/bl_0_101 sky130_rom_krom_rom_base_array_0/bl_0_102
+ sky130_rom_krom_rom_base_array_0/bl_0_103 sky130_rom_krom_rom_base_array_0/bl_0_104
+ sky130_rom_krom_rom_base_array_0/bl_0_105 sky130_rom_krom_rom_base_array_0/bl_0_106
+ sky130_rom_krom_rom_base_array_0/bl_0_107 sky130_rom_krom_rom_base_array_0/bl_0_108
+ sky130_rom_krom_rom_base_array_0/bl_0_109 sky130_rom_krom_rom_base_array_0/bl_0_110
+ sky130_rom_krom_rom_base_array_0/bl_0_111 sky130_rom_krom_rom_base_array_0/bl_0_112
+ sky130_rom_krom_rom_base_array_0/bl_0_113 sky130_rom_krom_rom_base_array_0/bl_0_114
+ sky130_rom_krom_rom_base_array_0/bl_0_115 sky130_rom_krom_rom_base_array_0/bl_0_116
+ sky130_rom_krom_rom_base_array_0/bl_0_117 sky130_rom_krom_rom_base_array_0/bl_0_119
+ sky130_rom_krom_rom_base_array_0/bl_0_120 sky130_rom_krom_rom_base_array_0/bl_0_121
+ sky130_rom_krom_rom_base_array_0/bl_0_122 sky130_rom_krom_rom_base_array_0/bl_0_123
+ sky130_rom_krom_rom_base_array_0/bl_0_124 sky130_rom_krom_rom_base_array_0/bl_0_125
+ sky130_rom_krom_rom_base_array_0/bl_0_126 sky130_rom_krom_rom_base_array_0/bl_0_127
+ sky130_rom_krom_rom_base_array_0/bl_0_128 sky130_rom_krom_rom_base_array_0/bl_0_129
+ sky130_rom_krom_rom_base_array_0/bl_0_130 sky130_rom_krom_rom_base_array_0/bl_0_131
+ sky130_rom_krom_rom_base_array_0/bl_0_132 sky130_rom_krom_rom_base_array_0/bl_0_133
+ sky130_rom_krom_rom_base_array_0/bl_0_134 sky130_rom_krom_rom_base_array_0/bl_0_135
+ sky130_rom_krom_rom_base_array_0/bl_0_136 sky130_rom_krom_rom_base_array_0/bl_0_137
+ sky130_rom_krom_rom_base_array_0/bl_0_138 sky130_rom_krom_rom_base_array_0/bl_0_139
+ sky130_rom_krom_rom_base_array_0/bl_0_140 sky130_rom_krom_rom_base_array_0/bl_0_141
+ sky130_rom_krom_rom_base_array_0/bl_0_142 sky130_rom_krom_rom_base_array_0/bl_0_143
+ sky130_rom_krom_rom_base_array_0/bl_0_144 sky130_rom_krom_rom_base_array_0/bl_0_145
+ sky130_rom_krom_rom_base_array_0/bl_0_146 sky130_rom_krom_rom_base_array_0/bl_0_147
+ sky130_rom_krom_rom_base_array_0/bl_0_148 sky130_rom_krom_rom_base_array_0/bl_0_149
+ sky130_rom_krom_rom_base_array_0/bl_0_150 sky130_rom_krom_rom_base_array_0/bl_0_151
+ sky130_rom_krom_rom_base_array_0/bl_0_152 sky130_rom_krom_rom_base_array_0/bl_0_153
+ sky130_rom_krom_rom_base_array_0/bl_0_154 sky130_rom_krom_rom_base_array_0/bl_0_155
+ sky130_rom_krom_rom_base_array_0/bl_0_156 sky130_rom_krom_rom_base_array_0/bl_0_157
+ sky130_rom_krom_rom_base_array_0/bl_0_158 sky130_rom_krom_rom_base_array_0/bl_0_159
+ sky130_rom_krom_rom_base_array_0/bl_0_160 sky130_rom_krom_rom_base_array_0/bl_0_161
+ sky130_rom_krom_rom_base_array_0/bl_0_162 sky130_rom_krom_rom_base_array_0/bl_0_163
+ sky130_rom_krom_rom_base_array_0/bl_0_164 sky130_rom_krom_rom_base_array_0/bl_0_165
+ sky130_rom_krom_rom_base_array_0/bl_0_167 sky130_rom_krom_rom_base_array_0/bl_0_168
+ sky130_rom_krom_rom_base_array_0/bl_0_169 sky130_rom_krom_rom_base_array_0/bl_0_170
+ sky130_rom_krom_rom_base_array_0/bl_0_171 sky130_rom_krom_rom_base_array_0/bl_0_172
+ sky130_rom_krom_rom_base_array_0/bl_0_173 sky130_rom_krom_rom_base_array_0/bl_0_174
+ sky130_rom_krom_rom_base_array_0/bl_0_175 sky130_rom_krom_rom_base_array_0/bl_0_176
+ sky130_rom_krom_rom_base_array_0/bl_0_177 sky130_rom_krom_rom_base_array_0/bl_0_178
+ sky130_rom_krom_rom_base_array_0/bl_0_179 sky130_rom_krom_rom_base_array_0/bl_0_180
+ sky130_rom_krom_rom_base_array_0/bl_0_181 sky130_rom_krom_rom_base_array_0/bl_0_182
+ sky130_rom_krom_rom_base_array_0/bl_0_183 sky130_rom_krom_rom_base_array_0/bl_0_184
+ sky130_rom_krom_rom_base_array_0/bl_0_185 sky130_rom_krom_rom_base_array_0/bl_0_186
+ sky130_rom_krom_rom_base_array_0/bl_0_187 sky130_rom_krom_rom_base_array_0/bl_0_188
+ sky130_rom_krom_rom_base_array_0/bl_0_189 sky130_rom_krom_rom_base_array_0/bl_0_190
+ sky130_rom_krom_rom_base_array_0/bl_0_191 sky130_rom_krom_rom_base_array_0/bl_0_192
+ sky130_rom_krom_rom_base_array_0/bl_0_193 sky130_rom_krom_rom_base_array_0/bl_0_194
+ sky130_rom_krom_rom_base_array_0/bl_0_195 sky130_rom_krom_rom_base_array_0/bl_0_196
+ sky130_rom_krom_rom_base_array_0/bl_0_197 sky130_rom_krom_rom_base_array_0/bl_0_198
+ sky130_rom_krom_rom_base_array_0/bl_0_199 sky130_rom_krom_rom_base_array_0/bl_0_200
+ sky130_rom_krom_rom_base_array_0/bl_0_201 sky130_rom_krom_rom_base_array_0/bl_0_202
+ sky130_rom_krom_rom_base_array_0/bl_0_203 sky130_rom_krom_rom_base_array_0/bl_0_204
+ sky130_rom_krom_rom_base_array_0/bl_0_205 sky130_rom_krom_rom_base_array_0/bl_0_206
+ sky130_rom_krom_rom_base_array_0/bl_0_207 sky130_rom_krom_rom_base_array_0/bl_0_208
+ sky130_rom_krom_rom_base_array_0/bl_0_209 sky130_rom_krom_rom_base_array_0/bl_0_210
+ sky130_rom_krom_rom_base_array_0/bl_0_211 sky130_rom_krom_rom_base_array_0/bl_0_213
+ sky130_rom_krom_rom_base_array_0/bl_0_214 sky130_rom_krom_rom_base_array_0/bl_0_215
+ sky130_rom_krom_rom_base_array_0/bl_0_216 sky130_rom_krom_rom_base_array_0/bl_0_217
+ sky130_rom_krom_rom_base_array_0/bl_0_218 sky130_rom_krom_rom_base_array_0/bl_0_219
+ sky130_rom_krom_rom_base_array_0/bl_0_220 sky130_rom_krom_rom_base_array_0/bl_0_221
+ sky130_rom_krom_rom_base_array_0/bl_0_222 sky130_rom_krom_rom_base_array_0/bl_0_223
+ sky130_rom_krom_rom_base_array_0/bl_0_224 sky130_rom_krom_rom_base_array_0/bl_0_225
+ sky130_rom_krom_rom_base_array_0/bl_0_226 sky130_rom_krom_rom_base_array_0/bl_0_227
+ sky130_rom_krom_rom_base_array_0/bl_0_228 sky130_rom_krom_rom_base_array_0/bl_0_229
+ sky130_rom_krom_rom_base_array_0/bl_0_230 sky130_rom_krom_rom_base_array_0/bl_0_231
+ sky130_rom_krom_rom_base_array_0/bl_0_232 sky130_rom_krom_rom_base_array_0/bl_0_233
+ sky130_rom_krom_rom_base_array_0/bl_0_234 sky130_rom_krom_rom_base_array_0/bl_0_235
+ sky130_rom_krom_rom_base_array_0/bl_0_236 sky130_rom_krom_rom_base_array_0/bl_0_237
+ sky130_rom_krom_rom_base_array_0/bl_0_238 sky130_rom_krom_rom_base_array_0/bl_0_239
+ sky130_rom_krom_rom_base_array_0/bl_0_240 sky130_rom_krom_rom_base_array_0/bl_0_241
+ sky130_rom_krom_rom_base_array_0/bl_0_242 sky130_rom_krom_rom_base_array_0/bl_0_243
+ sky130_rom_krom_rom_base_array_0/bl_0_244 sky130_rom_krom_rom_base_array_0/bl_0_245
+ sky130_rom_krom_rom_base_array_0/bl_0_246 sky130_rom_krom_rom_base_array_0/bl_0_247
+ sky130_rom_krom_rom_base_array_0/bl_0_248 sky130_rom_krom_rom_base_array_0/bl_0_249
+ sky130_rom_krom_rom_base_array_0/bl_0_250 sky130_rom_krom_rom_base_array_0/bl_0_251
+ sky130_rom_krom_rom_base_array_0/bl_0_252 sky130_rom_krom_rom_base_array_0/bl_0_253
+ sky130_rom_krom_rom_base_array_0/bl_0_254 sky130_rom_krom_rom_base_array_0/bl_0_255
+ sky130_rom_krom_rom_column_mux_array_0/bl_0 sky130_rom_krom_rom_column_mux_array_0/bl_1
+ sky130_rom_krom_rom_column_mux_array_0/bl_2 sky130_rom_krom_rom_column_mux_array_0/bl_3
+ sky130_rom_krom_rom_column_mux_array_0/bl_4 sky130_rom_krom_rom_column_mux_array_0/bl_5
+ sky130_rom_krom_rom_column_mux_array_0/bl_7 sky130_rom_krom_rom_column_mux_array_0/bl_8
+ sky130_rom_krom_rom_column_mux_array_0/bl_9 sky130_rom_krom_rom_column_mux_array_0/bl_10
+ sky130_rom_krom_rom_column_mux_array_0/bl_11 sky130_rom_krom_rom_column_mux_array_0/bl_12
+ sky130_rom_krom_rom_column_mux_array_0/bl_14 sky130_rom_krom_rom_column_mux_array_0/bl_15
+ sky130_rom_krom_rom_column_mux_array_0/bl_16 sky130_rom_krom_rom_column_mux_array_0/bl_17
+ sky130_rom_krom_rom_column_mux_array_0/bl_18 sky130_rom_krom_rom_column_mux_array_0/bl_19
+ sky130_rom_krom_rom_column_mux_array_0/bl_20 sky130_rom_krom_rom_column_mux_array_0/bl_21
+ sky130_rom_krom_rom_column_mux_array_0/bl_22 sky130_rom_krom_rom_column_mux_array_0/bl_23
+ sky130_rom_krom_rom_column_mux_array_0/bl_24 sky130_rom_krom_rom_column_mux_array_0/bl_25
+ sky130_rom_krom_rom_column_mux_array_0/bl_26 sky130_rom_krom_rom_column_mux_array_0/bl_27
+ sky130_rom_krom_rom_column_mux_array_0/bl_28 sky130_rom_krom_rom_column_mux_array_0/bl_29
+ sky130_rom_krom_rom_column_mux_array_0/bl_30 sky130_rom_krom_rom_column_mux_array_0/bl_31
+ sky130_rom_krom_rom_column_mux_array_0/bl_32 sky130_rom_krom_rom_column_mux_array_0/bl_33
+ sky130_rom_krom_rom_column_mux_array_0/bl_34 sky130_rom_krom_rom_column_mux_array_0/bl_35
+ sky130_rom_krom_rom_column_mux_array_0/bl_36 sky130_rom_krom_rom_column_mux_array_0/bl_37
+ sky130_rom_krom_rom_column_mux_array_0/bl_38 sky130_rom_krom_rom_column_mux_array_0/bl_39
+ sky130_rom_krom_rom_column_mux_array_0/bl_40 sky130_rom_krom_rom_column_mux_array_0/bl_41
+ sky130_rom_krom_rom_column_mux_array_0/bl_42 sky130_rom_krom_rom_column_mux_array_0/bl_43
+ sky130_rom_krom_rom_column_mux_array_0/bl_44 sky130_rom_krom_rom_column_mux_array_0/bl_45
+ sky130_rom_krom_rom_column_mux_array_0/bl_46 sky130_rom_krom_rom_column_mux_array_0/bl_47
+ sky130_rom_krom_rom_column_mux_array_0/bl_48 sky130_rom_krom_rom_column_mux_array_0/bl_49
+ sky130_rom_krom_rom_column_mux_array_0/bl_50 sky130_rom_krom_rom_column_mux_array_0/bl_51
+ sky130_rom_krom_rom_column_mux_array_0/bl_52 sky130_rom_krom_rom_column_mux_array_0/bl_53
+ sky130_rom_krom_rom_column_mux_array_0/bl_54 sky130_rom_krom_rom_column_mux_array_0/bl_55
+ sky130_rom_krom_rom_column_mux_array_0/bl_56 sky130_rom_krom_rom_column_mux_array_0/bl_57
+ sky130_rom_krom_rom_column_mux_array_0/bl_58 sky130_rom_krom_rom_column_mux_array_0/bl_59
+ sky130_rom_krom_rom_column_mux_array_0/bl_60 sky130_rom_krom_rom_column_mux_array_0/bl_62
+ sky130_rom_krom_rom_column_mux_array_0/bl_63 sky130_rom_krom_rom_column_mux_array_0/bl_64
+ sky130_rom_krom_rom_column_mux_array_0/bl_65 sky130_rom_krom_rom_column_mux_array_0/bl_66
+ sky130_rom_krom_rom_column_mux_array_0/bl_67 sky130_rom_krom_rom_column_mux_array_0/bl_68
+ sky130_rom_krom_rom_column_mux_array_0/bl_69 sky130_rom_krom_rom_column_mux_array_0/bl_70
+ sky130_rom_krom_rom_column_mux_array_0/bl_71 sky130_rom_krom_rom_column_mux_array_0/bl_72
+ sky130_rom_krom_rom_column_mux_array_0/bl_73 sky130_rom_krom_rom_column_mux_array_0/bl_74
+ sky130_rom_krom_rom_column_mux_array_0/bl_75 sky130_rom_krom_rom_column_mux_array_0/bl_76
+ sky130_rom_krom_rom_column_mux_array_0/bl_77 sky130_rom_krom_rom_column_mux_array_0/bl_78
+ sky130_rom_krom_rom_column_mux_array_0/bl_79 sky130_rom_krom_rom_column_mux_array_0/bl_80
+ sky130_rom_krom_rom_column_mux_array_0/bl_81 sky130_rom_krom_rom_column_mux_array_0/bl_82
+ sky130_rom_krom_rom_column_mux_array_0/bl_83 sky130_rom_krom_rom_column_mux_array_0/bl_84
+ sky130_rom_krom_rom_column_mux_array_0/bl_85 sky130_rom_krom_rom_column_mux_array_0/bl_86
+ sky130_rom_krom_rom_column_mux_array_0/bl_87 sky130_rom_krom_rom_column_mux_array_0/bl_88
+ sky130_rom_krom_rom_column_mux_array_0/bl_89 sky130_rom_krom_rom_column_mux_array_0/bl_90
+ sky130_rom_krom_rom_column_mux_array_0/bl_91 sky130_rom_krom_rom_column_mux_array_0/bl_92
+ sky130_rom_krom_rom_column_mux_array_0/bl_93 sky130_rom_krom_rom_column_mux_array_0/bl_94
+ sky130_rom_krom_rom_column_mux_array_0/bl_95 sky130_rom_krom_rom_column_mux_array_0/bl_96
+ sky130_rom_krom_rom_column_mux_array_0/bl_97 sky130_rom_krom_rom_column_mux_array_0/bl_98
+ sky130_rom_krom_rom_column_mux_array_0/bl_99 sky130_rom_krom_rom_column_mux_array_0/bl_100
+ sky130_rom_krom_rom_column_mux_array_0/bl_101 sky130_rom_krom_rom_column_mux_array_0/bl_102
+ sky130_rom_krom_rom_column_mux_array_0/bl_103 sky130_rom_krom_rom_column_mux_array_0/bl_104
+ sky130_rom_krom_rom_column_mux_array_0/bl_105 sky130_rom_krom_rom_column_mux_array_0/bl_106
+ sky130_rom_krom_rom_column_mux_array_0/bl_107 sky130_rom_krom_rom_column_mux_array_0/bl_108
+ sky130_rom_krom_rom_column_mux_array_0/bl_109 sky130_rom_krom_rom_column_mux_array_0/bl_110
+ sky130_rom_krom_rom_column_mux_array_0/bl_111 sky130_rom_krom_rom_column_mux_array_0/bl_112
+ sky130_rom_krom_rom_column_mux_array_0/bl_113 sky130_rom_krom_rom_column_mux_array_0/bl_114
+ sky130_rom_krom_rom_column_mux_array_0/bl_115 sky130_rom_krom_rom_column_mux_array_0/bl_116
+ sky130_rom_krom_rom_column_mux_array_0/bl_117 sky130_rom_krom_rom_column_mux_array_0/bl_118
+ sky130_rom_krom_rom_column_mux_array_0/bl_119 sky130_rom_krom_rom_column_mux_array_0/bl_120
+ sky130_rom_krom_rom_column_mux_array_0/bl_121 sky130_rom_krom_rom_column_mux_array_0/bl_122
+ sky130_rom_krom_rom_column_mux_array_0/bl_123 sky130_rom_krom_rom_column_mux_array_0/bl_124
+ sky130_rom_krom_rom_column_mux_array_0/bl_125 sky130_rom_krom_rom_column_mux_array_0/bl_126
+ sky130_rom_krom_rom_column_mux_array_0/bl_127 sky130_rom_krom_rom_column_mux_array_0/bl_128
+ sky130_rom_krom_rom_column_mux_array_0/bl_129 sky130_rom_krom_rom_column_mux_array_0/bl_130
+ sky130_rom_krom_rom_column_mux_array_0/bl_131 sky130_rom_krom_rom_column_mux_array_0/bl_132
+ sky130_rom_krom_rom_column_mux_array_0/bl_133 sky130_rom_krom_rom_column_mux_array_0/bl_134
+ sky130_rom_krom_rom_column_mux_array_0/bl_135 sky130_rom_krom_rom_column_mux_array_0/bl_136
+ sky130_rom_krom_rom_column_mux_array_0/bl_137 sky130_rom_krom_rom_column_mux_array_0/bl_138
+ sky130_rom_krom_rom_column_mux_array_0/bl_139 sky130_rom_krom_rom_column_mux_array_0/bl_140
+ sky130_rom_krom_rom_column_mux_array_0/bl_141 sky130_rom_krom_rom_column_mux_array_0/bl_142
+ sky130_rom_krom_rom_column_mux_array_0/bl_143 sky130_rom_krom_rom_column_mux_array_0/bl_144
+ sky130_rom_krom_rom_column_mux_array_0/bl_145 sky130_rom_krom_rom_column_mux_array_0/bl_146
+ sky130_rom_krom_rom_column_mux_array_0/bl_147 sky130_rom_krom_rom_column_mux_array_0/bl_148
+ sky130_rom_krom_rom_column_mux_array_0/bl_149 sky130_rom_krom_rom_column_mux_array_0/bl_150
+ sky130_rom_krom_rom_column_mux_array_0/bl_151 sky130_rom_krom_rom_column_mux_array_0/bl_152
+ sky130_rom_krom_rom_column_mux_array_0/bl_153 sky130_rom_krom_rom_column_mux_array_0/bl_154
+ sky130_rom_krom_rom_column_mux_array_0/bl_155 sky130_rom_krom_rom_column_mux_array_0/bl_156
+ sky130_rom_krom_rom_column_mux_array_0/bl_157 sky130_rom_krom_rom_column_mux_array_0/bl_158
+ sky130_rom_krom_rom_column_mux_array_0/bl_159 sky130_rom_krom_rom_column_mux_array_0/bl_160
+ sky130_rom_krom_rom_column_mux_array_0/bl_161 sky130_rom_krom_rom_column_mux_array_0/bl_162
+ sky130_rom_krom_rom_column_mux_array_0/bl_163 sky130_rom_krom_rom_column_mux_array_0/bl_164
+ sky130_rom_krom_rom_column_mux_array_0/bl_165 sky130_rom_krom_rom_column_mux_array_0/bl_166
+ sky130_rom_krom_rom_column_mux_array_0/bl_167 sky130_rom_krom_rom_column_mux_array_0/bl_168
+ sky130_rom_krom_rom_column_mux_array_0/bl_169 sky130_rom_krom_rom_column_mux_array_0/bl_170
+ sky130_rom_krom_rom_column_mux_array_0/bl_171 sky130_rom_krom_rom_column_mux_array_0/bl_172
+ sky130_rom_krom_rom_column_mux_array_0/bl_173 sky130_rom_krom_rom_column_mux_array_0/bl_174
+ sky130_rom_krom_rom_column_mux_array_0/bl_175 sky130_rom_krom_rom_column_mux_array_0/bl_176
+ sky130_rom_krom_rom_column_mux_array_0/bl_177 sky130_rom_krom_rom_column_mux_array_0/bl_178
+ sky130_rom_krom_rom_column_mux_array_0/bl_179 sky130_rom_krom_rom_column_mux_array_0/bl_180
+ sky130_rom_krom_rom_column_mux_array_0/bl_181 sky130_rom_krom_rom_column_mux_array_0/bl_182
+ sky130_rom_krom_rom_column_mux_array_0/bl_183 sky130_rom_krom_rom_column_mux_array_0/bl_184
+ sky130_rom_krom_rom_column_mux_array_0/bl_185 sky130_rom_krom_rom_column_mux_array_0/bl_186
+ sky130_rom_krom_rom_column_mux_array_0/bl_187 sky130_rom_krom_rom_column_mux_array_0/bl_188
+ sky130_rom_krom_rom_column_mux_array_0/bl_189 sky130_rom_krom_rom_column_mux_array_0/bl_190
+ sky130_rom_krom_rom_column_mux_array_0/bl_191 sky130_rom_krom_rom_column_mux_array_0/bl_192
+ sky130_rom_krom_rom_column_mux_array_0/bl_193 sky130_rom_krom_rom_column_mux_array_0/bl_194
+ sky130_rom_krom_rom_column_mux_array_0/bl_195 sky130_rom_krom_rom_column_mux_array_0/bl_196
+ sky130_rom_krom_rom_column_mux_array_0/bl_197 sky130_rom_krom_rom_column_mux_array_0/bl_198
+ sky130_rom_krom_rom_column_mux_array_0/bl_199 sky130_rom_krom_rom_column_mux_array_0/bl_200
+ sky130_rom_krom_rom_column_mux_array_0/bl_201 sky130_rom_krom_rom_column_mux_array_0/bl_202
+ sky130_rom_krom_rom_column_mux_array_0/bl_203 sky130_rom_krom_rom_column_mux_array_0/bl_204
+ sky130_rom_krom_rom_column_mux_array_0/bl_205 sky130_rom_krom_rom_column_mux_array_0/bl_206
+ sky130_rom_krom_rom_column_mux_array_0/bl_207 sky130_rom_krom_rom_column_mux_array_0/bl_208
+ sky130_rom_krom_rom_column_mux_array_0/bl_209 sky130_rom_krom_rom_column_mux_array_0/bl_210
+ sky130_rom_krom_rom_column_mux_array_0/bl_211 sky130_rom_krom_rom_column_mux_array_0/bl_213
+ sky130_rom_krom_rom_column_mux_array_0/bl_214 sky130_rom_krom_rom_column_mux_array_0/bl_215
+ sky130_rom_krom_rom_column_mux_array_0/bl_216 sky130_rom_krom_rom_column_mux_array_0/bl_217
+ sky130_rom_krom_rom_column_mux_array_0/bl_218 sky130_rom_krom_rom_column_mux_array_0/bl_219
+ sky130_rom_krom_rom_column_mux_array_0/bl_220 sky130_rom_krom_rom_column_mux_array_0/bl_221
+ sky130_rom_krom_rom_column_mux_array_0/bl_222 sky130_rom_krom_rom_column_mux_array_0/bl_223
+ sky130_rom_krom_rom_column_mux_array_0/bl_224 sky130_rom_krom_rom_column_mux_array_0/bl_225
+ sky130_rom_krom_rom_column_mux_array_0/bl_226 sky130_rom_krom_rom_column_mux_array_0/bl_227
+ sky130_rom_krom_rom_column_mux_array_0/bl_228 sky130_rom_krom_rom_column_mux_array_0/bl_229
+ sky130_rom_krom_rom_column_mux_array_0/bl_230 sky130_rom_krom_rom_column_mux_array_0/bl_231
+ sky130_rom_krom_rom_column_mux_array_0/bl_232 sky130_rom_krom_rom_column_mux_array_0/bl_233
+ sky130_rom_krom_rom_column_mux_array_0/bl_234 sky130_rom_krom_rom_column_mux_array_0/bl_235
+ sky130_rom_krom_rom_column_mux_array_0/bl_236 sky130_rom_krom_rom_column_mux_array_0/bl_237
+ sky130_rom_krom_rom_column_mux_array_0/bl_238 sky130_rom_krom_rom_column_mux_array_0/bl_239
+ sky130_rom_krom_rom_column_mux_array_0/bl_240 sky130_rom_krom_rom_column_mux_array_0/bl_241
+ sky130_rom_krom_rom_column_mux_array_0/bl_242 sky130_rom_krom_rom_column_mux_array_0/bl_243
+ sky130_rom_krom_rom_column_mux_array_0/bl_244 sky130_rom_krom_rom_column_mux_array_0/bl_245
+ sky130_rom_krom_rom_column_mux_array_0/bl_246 sky130_rom_krom_rom_column_mux_array_0/bl_247
+ sky130_rom_krom_rom_column_mux_array_0/bl_248 sky130_rom_krom_rom_column_mux_array_0/bl_249
+ sky130_rom_krom_rom_column_mux_array_0/bl_250 sky130_rom_krom_rom_column_mux_array_0/bl_251
+ sky130_rom_krom_rom_column_mux_array_0/bl_252 sky130_rom_krom_rom_column_mux_array_0/bl_253
+ sky130_rom_krom_rom_column_mux_array_0/bl_254 sky130_rom_krom_rom_column_mux_array_0/bl_255
+ sky130_rom_krom_rom_bitline_inverter_0/vdd sky130_rom_krom_rom_base_array_0/bl_0_15
+ gnd sky130_rom_krom_rom_base_array_0/bl_0_118 sky130_rom_krom_rom_base_array_0/bl_0_212
+ sky130_rom_krom_rom_column_mux_array_0/bl_13 sky130_rom_krom_rom_column_mux_array_0/bl_6
+ sky130_rom_krom_rom_base_array_0/bl_0_166 sky130_rom_krom_rom_column_mux_array_0/bl_212
+ sky130_rom_krom_rom_column_mux_array_0/bl_61 sky130_rom_krom_rom_base_array_0/vdd
+ sky130_rom_krom_rom_bitline_inverter
Xsky130_rom_krom_rom_column_decode_0 addr0[0] addr0[1] addr0[2] sky130_rom_krom_rom_column_decode_0/wl_0
+ sky130_rom_krom_rom_column_decode_0/wl_1 sky130_rom_krom_rom_column_decode_0/wl_2
+ sky130_rom_krom_rom_column_decode_0/wl_3 sky130_rom_krom_rom_column_decode_0/wl_4
+ sky130_rom_krom_rom_column_decode_0/wl_5 sky130_rom_krom_rom_column_decode_0/wl_6
+ sky130_rom_krom_rom_column_decode_0/wl_7 sky130_rom_krom_rom_column_decode_0/clk
+ sky130_rom_krom_rom_column_decode_0/vdd_uq0 sky130_rom_krom_rom_column_decode_0/vdd_uq2
+ sky130_rom_krom_rom_column_decode_0/vdd_uq4 sky130_rom_krom_rom_column_decode_0/vdd
+ sky130_rom_krom_rom_column_decode_0/clk sky130_rom_krom_rom_column_decode_0/vdd_uq1
+ gnd sky130_rom_krom_rom_column_decode
.ends

