magic
tech sky130A
magscale 1 2
timestamp 1581320207
<< checkpaint >>
rect -1296 -1309 3892 6566
<< locali >>
rect 1265 5240 1281 5274
rect 1315 5240 1331 5274
rect 64 3997 98 4013
rect 64 3947 98 3963
rect 2087 3925 2121 3959
rect 973 2611 989 2645
rect 1023 2611 1039 2645
rect 2342 2383 2376 2399
rect 2342 2333 2376 2349
rect 64 1244 98 1310
rect 1611 1232 1645 1248
rect 1611 1182 1645 1198
rect 2224 535 2258 551
rect 2224 485 2258 501
rect 2124 237 2158 303
rect 973 -17 989 17
rect 1023 -17 1039 17
<< viali >>
rect 1281 5240 1315 5274
rect 64 3963 98 3997
rect 989 2611 1023 2645
rect 2342 2349 2376 2383
rect 1611 1198 1645 1232
rect 2224 501 2258 535
rect 989 -17 1023 17
<< metal1 >>
rect 1272 5283 1324 5289
rect 1272 5225 1324 5231
rect 52 3997 110 4003
rect 52 3963 64 3997
rect 98 3963 110 3997
rect 52 3957 110 3963
rect 67 3882 95 3957
rect 67 3854 2373 3882
rect 980 2654 1032 2660
rect 980 2596 1032 2602
rect 2345 2389 2373 3854
rect 2330 2383 2388 2389
rect 2330 2349 2342 2383
rect 2376 2349 2388 2383
rect 2330 2343 2388 2349
rect 1599 1232 1657 1238
rect 1599 1198 1611 1232
rect 1645 1198 1657 1232
rect 1599 1192 1657 1198
rect 1614 532 1642 1192
rect 2212 535 2270 541
rect 2212 532 2224 535
rect 1614 504 2224 532
rect 2212 501 2224 504
rect 2258 501 2270 535
rect 2212 495 2270 501
rect 980 26 1032 32
rect 980 -32 1032 -26
<< via1 >>
rect 1272 5274 1324 5283
rect 1272 5240 1281 5274
rect 1281 5240 1315 5274
rect 1315 5240 1324 5274
rect 1272 5231 1324 5240
rect 980 2645 1032 2654
rect 980 2611 989 2645
rect 989 2611 1023 2645
rect 1023 2611 1032 2645
rect 980 2602 1032 2611
rect 980 17 1032 26
rect 980 -17 989 17
rect 989 -17 1023 17
rect 1023 -17 1032 17
rect 980 -26 1032 -17
<< metal2 >>
rect 1261 5229 1270 5285
rect 1326 5229 1335 5285
rect 969 2600 978 2656
rect 1034 2600 1043 2656
rect 969 -28 978 28
rect 1034 -28 1043 28
<< via2 >>
rect 1270 5283 1326 5285
rect 1270 5231 1272 5283
rect 1272 5231 1324 5283
rect 1324 5231 1326 5283
rect 1270 5229 1326 5231
rect 978 2654 1034 2656
rect 978 2602 980 2654
rect 980 2602 1032 2654
rect 1032 2602 1034 2654
rect 978 2600 1034 2602
rect 978 26 1034 28
rect 978 -26 980 26
rect 980 -26 1032 26
rect 1032 -26 1034 26
rect 978 -28 1034 -26
<< metal3 >>
rect 1249 5285 1347 5306
rect 1249 5229 1270 5285
rect 1326 5229 1347 5285
rect 1249 5208 1347 5229
rect 957 2656 1055 2677
rect 957 2600 978 2656
rect 1034 2600 1055 2656
rect 957 2579 1055 2600
rect 957 28 1055 49
rect 957 -28 978 28
rect 1034 -28 1055 28
rect 957 -49 1055 -28
use sky130_rom_krom_rom_clock_driver  sky130_rom_krom_rom_clock_driver_0
timestamp 1581320207
transform 1 0 0 0 1 0
box -36 -17 2048 2686
use sky130_rom_krom_rom_control_nand  sky130_rom_krom_rom_control_nand_0
timestamp 1581320207
transform 1 0 2012 0 1 0
box -36 -17 414 2686
use sky130_rom_krom_rom_precharge_driver  sky130_rom_krom_rom_precharge_driver_0
timestamp 1581320207
transform 1 0 0 0 -1 5257
box -36 -17 2632 2686
<< labels >>
rlabel locali s 81 1277 81 1277 4 clk_in
port 2 nsew
rlabel locali s 1628 1215 1628 1215 4 clk_out
port 3 nsew
rlabel locali s 2104 3942 2104 3942 4 prechrg
port 4 nsew
rlabel locali s 2141 270 2141 270 4 CS
port 5 nsew
rlabel metal3 s 1249 5208 1347 5306 4 gnd
port 7 nsew
rlabel metal3 s 957 -49 1055 49 4 gnd
port 7 nsew
rlabel metal3 s 957 2579 1055 2677 4 vdd
port 9 nsew
<< properties >>
string FIXED_BBOX 969 -33 1043 0
<< end >>
