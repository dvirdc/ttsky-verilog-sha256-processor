magic
tech sky130A
magscale 1 2
timestamp 1581320221
<< checkpaint >>
rect -2756 -2756 22930 18690
<< locali >>
rect 6723 15560 6757 15576
rect 6723 15510 6757 15526
rect 6723 15356 6757 15372
rect 6723 15306 6757 15322
rect 6723 15152 6757 15168
rect 6723 15102 6757 15118
rect 6723 14948 6757 14964
rect 6723 14898 6757 14914
rect 6723 14744 6757 14760
rect 6723 14694 6757 14710
rect 6723 14540 6757 14556
rect 6723 14490 6757 14506
rect 6723 14336 6757 14352
rect 6723 14286 6757 14302
rect 6723 14132 6757 14148
rect 6723 14082 6757 14098
rect 6723 13824 6757 13840
rect 6723 13774 6757 13790
rect 6723 13620 6757 13636
rect 6723 13570 6757 13586
rect 6723 13416 6757 13432
rect 6723 13366 6757 13382
rect 6723 13212 6757 13228
rect 6723 13162 6757 13178
rect 6723 13008 6757 13024
rect 6723 12958 6757 12974
rect 6723 12804 6757 12820
rect 6723 12754 6757 12770
rect 6723 12600 6757 12616
rect 6723 12550 6757 12566
rect 6723 12396 6757 12412
rect 6723 12346 6757 12362
rect 6723 12088 6757 12104
rect 6723 12038 6757 12054
rect 6723 11884 6757 11900
rect 6723 11834 6757 11850
rect 6723 11680 6757 11696
rect 6723 11630 6757 11646
rect 6723 11476 6757 11492
rect 6723 11426 6757 11442
rect 6723 11272 6757 11288
rect 6723 11222 6757 11238
rect 6723 11068 6757 11084
rect 6723 11018 6757 11034
rect 6723 10864 6757 10880
rect 6723 10814 6757 10830
rect 6723 10660 6757 10676
rect 6723 10610 6757 10626
rect 6723 10352 6757 10368
rect 6723 10302 6757 10318
rect 6723 10148 6757 10164
rect 6723 10098 6757 10114
rect 6723 9944 6757 9960
rect 6723 9894 6757 9910
rect 6723 9740 6757 9756
rect 6723 9690 6757 9706
rect 6723 9536 6757 9552
rect 6723 9486 6757 9502
rect 6723 9332 6757 9348
rect 6723 9282 6757 9298
rect 6723 9128 6757 9144
rect 6723 9078 6757 9094
rect 6723 8924 6757 8940
rect 6723 8874 6757 8890
rect 6978 7799 6994 7833
rect 7028 7799 7044 7833
rect 7182 7799 7198 7833
rect 7232 7799 7248 7833
rect 7386 7799 7402 7833
rect 7436 7799 7452 7833
rect 7590 7799 7606 7833
rect 7640 7799 7656 7833
rect 7794 7799 7810 7833
rect 7844 7799 7860 7833
rect 7998 7799 8014 7833
rect 8048 7799 8064 7833
rect 8202 7799 8218 7833
rect 8252 7799 8268 7833
rect 8406 7799 8422 7833
rect 8456 7799 8472 7833
rect 8610 7799 8626 7833
rect 8660 7799 8676 7833
rect 8814 7799 8830 7833
rect 8864 7799 8880 7833
rect 9018 7799 9034 7833
rect 9068 7799 9084 7833
rect 9222 7799 9238 7833
rect 9272 7799 9288 7833
rect 9426 7799 9442 7833
rect 9476 7799 9492 7833
rect 9630 7799 9646 7833
rect 9680 7799 9696 7833
rect 9834 7799 9850 7833
rect 9884 7799 9900 7833
rect 10038 7799 10054 7833
rect 10088 7799 10104 7833
rect 10242 7799 10258 7833
rect 10292 7799 10308 7833
rect 10446 7799 10462 7833
rect 10496 7799 10512 7833
rect 10650 7799 10666 7833
rect 10700 7799 10716 7833
rect 10854 7799 10870 7833
rect 10904 7799 10920 7833
rect 11058 7799 11074 7833
rect 11108 7799 11124 7833
rect 11262 7799 11278 7833
rect 11312 7799 11328 7833
rect 11466 7799 11482 7833
rect 11516 7799 11532 7833
rect 11670 7799 11686 7833
rect 11720 7799 11736 7833
rect 11874 7799 11890 7833
rect 11924 7799 11940 7833
rect 12078 7799 12094 7833
rect 12128 7799 12144 7833
rect 12282 7799 12298 7833
rect 12332 7799 12348 7833
rect 12486 7799 12502 7833
rect 12536 7799 12552 7833
rect 12690 7799 12706 7833
rect 12740 7799 12756 7833
rect 12894 7799 12910 7833
rect 12944 7799 12960 7833
rect 13098 7799 13114 7833
rect 13148 7799 13164 7833
rect 13302 7799 13318 7833
rect 13352 7799 13368 7833
rect 13506 7799 13522 7833
rect 13556 7799 13572 7833
rect 13710 7799 13726 7833
rect 13760 7799 13776 7833
rect 13914 7799 13930 7833
rect 13964 7799 13980 7833
rect 14118 7799 14134 7833
rect 14168 7799 14184 7833
rect 14322 7799 14338 7833
rect 14372 7799 14388 7833
rect 14526 7799 14542 7833
rect 14576 7799 14592 7833
rect 14730 7799 14746 7833
rect 14780 7799 14796 7833
rect 14934 7799 14950 7833
rect 14984 7799 15000 7833
rect 15138 7799 15154 7833
rect 15188 7799 15204 7833
rect 15342 7799 15358 7833
rect 15392 7799 15408 7833
rect 15546 7799 15562 7833
rect 15596 7799 15612 7833
rect 15750 7799 15766 7833
rect 15800 7799 15816 7833
rect 15954 7799 15970 7833
rect 16004 7799 16020 7833
rect 16158 7799 16174 7833
rect 16208 7799 16224 7833
rect 16362 7799 16378 7833
rect 16412 7799 16428 7833
rect 16566 7799 16582 7833
rect 16616 7799 16632 7833
rect 16770 7799 16786 7833
rect 16820 7799 16836 7833
rect 16974 7799 16990 7833
rect 17024 7799 17040 7833
rect 17178 7799 17194 7833
rect 17228 7799 17244 7833
rect 17382 7799 17398 7833
rect 17432 7799 17448 7833
rect 17586 7799 17602 7833
rect 17636 7799 17652 7833
rect 17790 7799 17806 7833
rect 17840 7799 17856 7833
rect 17994 7799 18010 7833
rect 18044 7799 18060 7833
rect 18198 7799 18214 7833
rect 18248 7799 18264 7833
rect 18402 7799 18418 7833
rect 18452 7799 18468 7833
rect 18606 7799 18622 7833
rect 18656 7799 18672 7833
rect 18810 7799 18826 7833
rect 18860 7799 18876 7833
rect 19014 7799 19030 7833
rect 19064 7799 19080 7833
rect 19218 7799 19234 7833
rect 19268 7799 19284 7833
rect 19422 7799 19438 7833
rect 19472 7799 19488 7833
rect 19626 7799 19642 7833
rect 19676 7799 19692 7833
rect 19830 7799 19846 7833
rect 19880 7799 19896 7833
rect 6978 6204 6994 6238
rect 7028 6204 7044 6238
rect 7182 6204 7198 6238
rect 7232 6204 7248 6238
rect 7386 6204 7402 6238
rect 7436 6204 7452 6238
rect 7590 6204 7606 6238
rect 7640 6204 7656 6238
rect 7794 6204 7810 6238
rect 7844 6204 7860 6238
rect 7998 6204 8014 6238
rect 8048 6204 8064 6238
rect 8202 6204 8218 6238
rect 8252 6204 8268 6238
rect 8406 6204 8422 6238
rect 8456 6204 8472 6238
rect 8610 6204 8626 6238
rect 8660 6204 8676 6238
rect 8814 6204 8830 6238
rect 8864 6204 8880 6238
rect 9018 6204 9034 6238
rect 9068 6204 9084 6238
rect 9222 6204 9238 6238
rect 9272 6204 9288 6238
rect 9426 6204 9442 6238
rect 9476 6204 9492 6238
rect 9630 6204 9646 6238
rect 9680 6204 9696 6238
rect 9834 6204 9850 6238
rect 9884 6204 9900 6238
rect 10038 6204 10054 6238
rect 10088 6204 10104 6238
rect 10242 6204 10258 6238
rect 10292 6204 10308 6238
rect 10446 6204 10462 6238
rect 10496 6204 10512 6238
rect 10650 6204 10666 6238
rect 10700 6204 10716 6238
rect 10854 6204 10870 6238
rect 10904 6204 10920 6238
rect 11058 6204 11074 6238
rect 11108 6204 11124 6238
rect 11262 6204 11278 6238
rect 11312 6204 11328 6238
rect 11466 6204 11482 6238
rect 11516 6204 11532 6238
rect 11670 6204 11686 6238
rect 11720 6204 11736 6238
rect 11874 6204 11890 6238
rect 11924 6204 11940 6238
rect 12078 6204 12094 6238
rect 12128 6204 12144 6238
rect 12282 6204 12298 6238
rect 12332 6204 12348 6238
rect 12486 6204 12502 6238
rect 12536 6204 12552 6238
rect 12690 6204 12706 6238
rect 12740 6204 12756 6238
rect 12894 6204 12910 6238
rect 12944 6204 12960 6238
rect 13098 6204 13114 6238
rect 13148 6204 13164 6238
rect 13302 6204 13318 6238
rect 13352 6204 13368 6238
rect 13506 6204 13522 6238
rect 13556 6204 13572 6238
rect 13710 6204 13726 6238
rect 13760 6204 13776 6238
rect 13914 6204 13930 6238
rect 13964 6204 13980 6238
rect 14118 6204 14134 6238
rect 14168 6204 14184 6238
rect 14322 6204 14338 6238
rect 14372 6204 14388 6238
rect 14526 6204 14542 6238
rect 14576 6204 14592 6238
rect 14730 6204 14746 6238
rect 14780 6204 14796 6238
rect 14934 6204 14950 6238
rect 14984 6204 15000 6238
rect 15138 6204 15154 6238
rect 15188 6204 15204 6238
rect 15342 6204 15358 6238
rect 15392 6204 15408 6238
rect 15546 6204 15562 6238
rect 15596 6204 15612 6238
rect 15750 6204 15766 6238
rect 15800 6204 15816 6238
rect 15954 6204 15970 6238
rect 16004 6204 16020 6238
rect 16158 6204 16174 6238
rect 16208 6204 16224 6238
rect 16362 6204 16378 6238
rect 16412 6204 16428 6238
rect 16566 6204 16582 6238
rect 16616 6204 16632 6238
rect 16770 6204 16786 6238
rect 16820 6204 16836 6238
rect 16974 6204 16990 6238
rect 17024 6204 17040 6238
rect 17178 6204 17194 6238
rect 17228 6204 17244 6238
rect 17382 6204 17398 6238
rect 17432 6204 17448 6238
rect 17586 6204 17602 6238
rect 17636 6204 17652 6238
rect 17790 6204 17806 6238
rect 17840 6204 17856 6238
rect 17994 6204 18010 6238
rect 18044 6204 18060 6238
rect 18198 6204 18214 6238
rect 18248 6204 18264 6238
rect 18402 6204 18418 6238
rect 18452 6204 18468 6238
rect 18606 6204 18622 6238
rect 18656 6204 18672 6238
rect 18810 6204 18826 6238
rect 18860 6204 18876 6238
rect 19014 6204 19030 6238
rect 19064 6204 19080 6238
rect 19218 6204 19234 6238
rect 19268 6204 19284 6238
rect 19422 6204 19438 6238
rect 19472 6204 19488 6238
rect 19626 6204 19642 6238
rect 19676 6204 19692 6238
rect 19830 6204 19846 6238
rect 19880 6204 19896 6238
rect 337 5563 371 5579
rect 337 5513 371 5529
rect 745 5563 779 5579
rect 745 5513 779 5529
rect 1153 5563 1187 5579
rect 1153 5513 1187 5529
rect 1561 5563 1595 5579
rect 1561 5513 1595 5529
rect 1969 5563 2003 5579
rect 1969 5513 2003 5529
rect 6723 4883 6757 4899
rect 6723 4833 6757 4849
rect 6723 4679 6757 4695
rect 6723 4629 6757 4645
rect 6723 4475 6757 4491
rect 6723 4425 6757 4441
rect 6723 4271 6757 4287
rect 6723 4221 6757 4237
rect 2513 4092 2547 4108
rect 2513 4042 2547 4058
rect 6723 4067 6757 4083
rect 6723 4017 6757 4033
rect 6723 3863 6757 3879
rect 6723 3813 6757 3829
rect 6723 3659 6757 3675
rect 6723 3609 6757 3625
rect 6723 3455 6757 3471
rect 6723 3405 6757 3421
rect 8560 2129 8594 2145
rect 8560 2079 8594 2095
rect 8868 2129 8902 2145
rect 8868 2079 8902 2095
rect 9176 2129 9210 2145
rect 9176 2079 9210 2095
rect 9484 2129 9518 2145
rect 9484 2079 9518 2095
rect 9792 2129 9826 2145
rect 9792 2079 9826 2095
rect 10100 2129 10134 2145
rect 10100 2079 10134 2095
rect 10408 2129 10442 2145
rect 10408 2079 10442 2095
rect 10716 2129 10750 2145
rect 10716 2079 10750 2095
rect 490 1427 524 1443
rect 490 1377 524 1393
rect 2037 1365 2071 1381
rect 2037 1315 2071 1331
rect 2550 420 2584 436
rect 8544 390 8560 424
rect 8594 390 8610 424
rect 8852 390 8868 424
rect 8902 390 8918 424
rect 9160 390 9176 424
rect 9210 390 9226 424
rect 9468 390 9484 424
rect 9518 390 9534 424
rect 9776 390 9792 424
rect 9826 390 9842 424
rect 10084 390 10100 424
rect 10134 390 10150 424
rect 10392 390 10408 424
rect 10442 390 10458 424
rect 10700 390 10716 424
rect 10750 390 10766 424
rect 2550 370 2584 386
rect 3599 94 3633 110
rect 3599 44 3633 60
rect 4007 94 4041 110
rect 4007 44 4041 60
rect 4415 94 4449 110
rect 4415 44 4449 60
<< viali >>
rect 6723 15526 6757 15560
rect 6723 15322 6757 15356
rect 6723 15118 6757 15152
rect 6723 14914 6757 14948
rect 6723 14710 6757 14744
rect 6723 14506 6757 14540
rect 6723 14302 6757 14336
rect 6723 14098 6757 14132
rect 6723 13790 6757 13824
rect 6723 13586 6757 13620
rect 6723 13382 6757 13416
rect 6723 13178 6757 13212
rect 6723 12974 6757 13008
rect 6723 12770 6757 12804
rect 6723 12566 6757 12600
rect 6723 12362 6757 12396
rect 6723 12054 6757 12088
rect 6723 11850 6757 11884
rect 6723 11646 6757 11680
rect 6723 11442 6757 11476
rect 6723 11238 6757 11272
rect 6723 11034 6757 11068
rect 6723 10830 6757 10864
rect 6723 10626 6757 10660
rect 6723 10318 6757 10352
rect 6723 10114 6757 10148
rect 6723 9910 6757 9944
rect 6723 9706 6757 9740
rect 6723 9502 6757 9536
rect 6723 9298 6757 9332
rect 6723 9094 6757 9128
rect 6723 8890 6757 8924
rect 6994 7799 7028 7833
rect 7198 7799 7232 7833
rect 7402 7799 7436 7833
rect 7606 7799 7640 7833
rect 7810 7799 7844 7833
rect 8014 7799 8048 7833
rect 8218 7799 8252 7833
rect 8422 7799 8456 7833
rect 8626 7799 8660 7833
rect 8830 7799 8864 7833
rect 9034 7799 9068 7833
rect 9238 7799 9272 7833
rect 9442 7799 9476 7833
rect 9646 7799 9680 7833
rect 9850 7799 9884 7833
rect 10054 7799 10088 7833
rect 10258 7799 10292 7833
rect 10462 7799 10496 7833
rect 10666 7799 10700 7833
rect 10870 7799 10904 7833
rect 11074 7799 11108 7833
rect 11278 7799 11312 7833
rect 11482 7799 11516 7833
rect 11686 7799 11720 7833
rect 11890 7799 11924 7833
rect 12094 7799 12128 7833
rect 12298 7799 12332 7833
rect 12502 7799 12536 7833
rect 12706 7799 12740 7833
rect 12910 7799 12944 7833
rect 13114 7799 13148 7833
rect 13318 7799 13352 7833
rect 13522 7799 13556 7833
rect 13726 7799 13760 7833
rect 13930 7799 13964 7833
rect 14134 7799 14168 7833
rect 14338 7799 14372 7833
rect 14542 7799 14576 7833
rect 14746 7799 14780 7833
rect 14950 7799 14984 7833
rect 15154 7799 15188 7833
rect 15358 7799 15392 7833
rect 15562 7799 15596 7833
rect 15766 7799 15800 7833
rect 15970 7799 16004 7833
rect 16174 7799 16208 7833
rect 16378 7799 16412 7833
rect 16582 7799 16616 7833
rect 16786 7799 16820 7833
rect 16990 7799 17024 7833
rect 17194 7799 17228 7833
rect 17398 7799 17432 7833
rect 17602 7799 17636 7833
rect 17806 7799 17840 7833
rect 18010 7799 18044 7833
rect 18214 7799 18248 7833
rect 18418 7799 18452 7833
rect 18622 7799 18656 7833
rect 18826 7799 18860 7833
rect 19030 7799 19064 7833
rect 19234 7799 19268 7833
rect 19438 7799 19472 7833
rect 19642 7799 19676 7833
rect 19846 7799 19880 7833
rect 6994 6204 7028 6238
rect 7198 6204 7232 6238
rect 7402 6204 7436 6238
rect 7606 6204 7640 6238
rect 7810 6204 7844 6238
rect 8014 6204 8048 6238
rect 8218 6204 8252 6238
rect 8422 6204 8456 6238
rect 8626 6204 8660 6238
rect 8830 6204 8864 6238
rect 9034 6204 9068 6238
rect 9238 6204 9272 6238
rect 9442 6204 9476 6238
rect 9646 6204 9680 6238
rect 9850 6204 9884 6238
rect 10054 6204 10088 6238
rect 10258 6204 10292 6238
rect 10462 6204 10496 6238
rect 10666 6204 10700 6238
rect 10870 6204 10904 6238
rect 11074 6204 11108 6238
rect 11278 6204 11312 6238
rect 11482 6204 11516 6238
rect 11686 6204 11720 6238
rect 11890 6204 11924 6238
rect 12094 6204 12128 6238
rect 12298 6204 12332 6238
rect 12502 6204 12536 6238
rect 12706 6204 12740 6238
rect 12910 6204 12944 6238
rect 13114 6204 13148 6238
rect 13318 6204 13352 6238
rect 13522 6204 13556 6238
rect 13726 6204 13760 6238
rect 13930 6204 13964 6238
rect 14134 6204 14168 6238
rect 14338 6204 14372 6238
rect 14542 6204 14576 6238
rect 14746 6204 14780 6238
rect 14950 6204 14984 6238
rect 15154 6204 15188 6238
rect 15358 6204 15392 6238
rect 15562 6204 15596 6238
rect 15766 6204 15800 6238
rect 15970 6204 16004 6238
rect 16174 6204 16208 6238
rect 16378 6204 16412 6238
rect 16582 6204 16616 6238
rect 16786 6204 16820 6238
rect 16990 6204 17024 6238
rect 17194 6204 17228 6238
rect 17398 6204 17432 6238
rect 17602 6204 17636 6238
rect 17806 6204 17840 6238
rect 18010 6204 18044 6238
rect 18214 6204 18248 6238
rect 18418 6204 18452 6238
rect 18622 6204 18656 6238
rect 18826 6204 18860 6238
rect 19030 6204 19064 6238
rect 19234 6204 19268 6238
rect 19438 6204 19472 6238
rect 19642 6204 19676 6238
rect 19846 6204 19880 6238
rect 337 5529 371 5563
rect 745 5529 779 5563
rect 1153 5529 1187 5563
rect 1561 5529 1595 5563
rect 1969 5529 2003 5563
rect 6723 4849 6757 4883
rect 6723 4645 6757 4679
rect 6723 4441 6757 4475
rect 6723 4237 6757 4271
rect 2513 4058 2547 4092
rect 6723 4033 6757 4067
rect 6723 3829 6757 3863
rect 6723 3625 6757 3659
rect 6723 3421 6757 3455
rect 8560 2095 8594 2129
rect 8868 2095 8902 2129
rect 9176 2095 9210 2129
rect 9484 2095 9518 2129
rect 9792 2095 9826 2129
rect 10100 2095 10134 2129
rect 10408 2095 10442 2129
rect 10716 2095 10750 2129
rect 490 1393 524 1427
rect 2037 1331 2071 1365
rect 2550 386 2584 420
rect 8560 390 8594 424
rect 8868 390 8902 424
rect 9176 390 9210 424
rect 9484 390 9518 424
rect 9792 390 9826 424
rect 10100 390 10134 424
rect 10408 390 10442 424
rect 10716 390 10750 424
rect 3599 60 3633 94
rect 4007 60 4041 94
rect 4415 60 4449 94
<< metal1 >>
rect 6965 15848 6971 15900
rect 7023 15848 7029 15900
rect 19845 15848 19851 15900
rect 19903 15848 19909 15900
rect 3321 15637 3327 15689
rect 3379 15637 3385 15689
rect 3943 15637 3949 15689
rect 4001 15637 4007 15689
rect 4741 15637 4747 15689
rect 4799 15637 4805 15689
rect 5989 15637 5995 15689
rect 6047 15637 6053 15689
rect 6711 15560 6769 15566
rect 6711 15526 6723 15560
rect 6757 15557 6769 15560
rect 6870 15557 6876 15569
rect 6757 15529 6876 15557
rect 6757 15526 6769 15529
rect 6711 15520 6769 15526
rect 6870 15517 6876 15529
rect 6928 15517 6934 15569
rect 6711 15356 6769 15362
rect 6711 15322 6723 15356
rect 6757 15353 6769 15356
rect 6870 15353 6876 15365
rect 6757 15325 6876 15353
rect 6757 15322 6769 15325
rect 6711 15316 6769 15322
rect 6870 15313 6876 15325
rect 6928 15313 6934 15365
rect 6711 15152 6769 15158
rect 6711 15118 6723 15152
rect 6757 15149 6769 15152
rect 6870 15149 6876 15161
rect 6757 15121 6876 15149
rect 6757 15118 6769 15121
rect 6711 15112 6769 15118
rect 6870 15109 6876 15121
rect 6928 15109 6934 15161
rect 6711 14948 6769 14954
rect 6711 14914 6723 14948
rect 6757 14945 6769 14948
rect 6870 14945 6876 14957
rect 6757 14917 6876 14945
rect 6757 14914 6769 14917
rect 6711 14908 6769 14914
rect 6870 14905 6876 14917
rect 6928 14905 6934 14957
rect 6711 14744 6769 14750
rect 6711 14710 6723 14744
rect 6757 14741 6769 14744
rect 6870 14741 6876 14753
rect 6757 14713 6876 14741
rect 6757 14710 6769 14713
rect 6711 14704 6769 14710
rect 6870 14701 6876 14713
rect 6928 14701 6934 14753
rect 6711 14540 6769 14546
rect 6711 14506 6723 14540
rect 6757 14537 6769 14540
rect 6870 14537 6876 14549
rect 6757 14509 6876 14537
rect 6757 14506 6769 14509
rect 6711 14500 6769 14506
rect 6870 14497 6876 14509
rect 6928 14497 6934 14549
rect 6711 14336 6769 14342
rect 6711 14302 6723 14336
rect 6757 14333 6769 14336
rect 6870 14333 6876 14345
rect 6757 14305 6876 14333
rect 6757 14302 6769 14305
rect 6711 14296 6769 14302
rect 6870 14293 6876 14305
rect 6928 14293 6934 14345
rect 6711 14132 6769 14138
rect 6711 14098 6723 14132
rect 6757 14129 6769 14132
rect 6870 14129 6876 14141
rect 6757 14101 6876 14129
rect 6757 14098 6769 14101
rect 6711 14092 6769 14098
rect 6870 14089 6876 14101
rect 6928 14089 6934 14141
rect 6711 13824 6769 13830
rect 6711 13790 6723 13824
rect 6757 13821 6769 13824
rect 6870 13821 6876 13833
rect 6757 13793 6876 13821
rect 6757 13790 6769 13793
rect 6711 13784 6769 13790
rect 6870 13781 6876 13793
rect 6928 13781 6934 13833
rect 6711 13620 6769 13626
rect 6711 13586 6723 13620
rect 6757 13617 6769 13620
rect 6870 13617 6876 13629
rect 6757 13589 6876 13617
rect 6757 13586 6769 13589
rect 6711 13580 6769 13586
rect 6870 13577 6876 13589
rect 6928 13577 6934 13629
rect 6711 13416 6769 13422
rect 6711 13382 6723 13416
rect 6757 13413 6769 13416
rect 6870 13413 6876 13425
rect 6757 13385 6876 13413
rect 6757 13382 6769 13385
rect 6711 13376 6769 13382
rect 6870 13373 6876 13385
rect 6928 13373 6934 13425
rect 6711 13212 6769 13218
rect 6711 13178 6723 13212
rect 6757 13209 6769 13212
rect 6870 13209 6876 13221
rect 6757 13181 6876 13209
rect 6757 13178 6769 13181
rect 6711 13172 6769 13178
rect 6870 13169 6876 13181
rect 6928 13169 6934 13221
rect 6711 13008 6769 13014
rect 6711 12974 6723 13008
rect 6757 13005 6769 13008
rect 6870 13005 6876 13017
rect 6757 12977 6876 13005
rect 6757 12974 6769 12977
rect 6711 12968 6769 12974
rect 6870 12965 6876 12977
rect 6928 12965 6934 13017
rect 6711 12804 6769 12810
rect 6711 12770 6723 12804
rect 6757 12801 6769 12804
rect 6870 12801 6876 12813
rect 6757 12773 6876 12801
rect 6757 12770 6769 12773
rect 6711 12764 6769 12770
rect 6870 12761 6876 12773
rect 6928 12761 6934 12813
rect 6711 12600 6769 12606
rect 6711 12566 6723 12600
rect 6757 12597 6769 12600
rect 6870 12597 6876 12609
rect 6757 12569 6876 12597
rect 6757 12566 6769 12569
rect 6711 12560 6769 12566
rect 6870 12557 6876 12569
rect 6928 12557 6934 12609
rect 6711 12396 6769 12402
rect 6711 12362 6723 12396
rect 6757 12393 6769 12396
rect 6870 12393 6876 12405
rect 6757 12365 6876 12393
rect 6757 12362 6769 12365
rect 6711 12356 6769 12362
rect 6870 12353 6876 12365
rect 6928 12353 6934 12405
rect 6711 12088 6769 12094
rect 6711 12054 6723 12088
rect 6757 12085 6769 12088
rect 6870 12085 6876 12097
rect 6757 12057 6876 12085
rect 6757 12054 6769 12057
rect 6711 12048 6769 12054
rect 6870 12045 6876 12057
rect 6928 12045 6934 12097
rect 6711 11884 6769 11890
rect 6711 11850 6723 11884
rect 6757 11881 6769 11884
rect 6870 11881 6876 11893
rect 6757 11853 6876 11881
rect 6757 11850 6769 11853
rect 6711 11844 6769 11850
rect 6870 11841 6876 11853
rect 6928 11841 6934 11893
rect 6711 11680 6769 11686
rect 6711 11646 6723 11680
rect 6757 11677 6769 11680
rect 6870 11677 6876 11689
rect 6757 11649 6876 11677
rect 6757 11646 6769 11649
rect 6711 11640 6769 11646
rect 6870 11637 6876 11649
rect 6928 11637 6934 11689
rect 6711 11476 6769 11482
rect 6711 11442 6723 11476
rect 6757 11473 6769 11476
rect 6870 11473 6876 11485
rect 6757 11445 6876 11473
rect 6757 11442 6769 11445
rect 6711 11436 6769 11442
rect 6870 11433 6876 11445
rect 6928 11433 6934 11485
rect 6711 11272 6769 11278
rect 6711 11238 6723 11272
rect 6757 11269 6769 11272
rect 6870 11269 6876 11281
rect 6757 11241 6876 11269
rect 6757 11238 6769 11241
rect 6711 11232 6769 11238
rect 6870 11229 6876 11241
rect 6928 11229 6934 11281
rect 6711 11068 6769 11074
rect 6711 11034 6723 11068
rect 6757 11065 6769 11068
rect 6870 11065 6876 11077
rect 6757 11037 6876 11065
rect 6757 11034 6769 11037
rect 6711 11028 6769 11034
rect 6870 11025 6876 11037
rect 6928 11025 6934 11077
rect 6711 10864 6769 10870
rect 6711 10830 6723 10864
rect 6757 10861 6769 10864
rect 6870 10861 6876 10873
rect 6757 10833 6876 10861
rect 6757 10830 6769 10833
rect 6711 10824 6769 10830
rect 6870 10821 6876 10833
rect 6928 10821 6934 10873
rect 6711 10660 6769 10666
rect 6711 10626 6723 10660
rect 6757 10657 6769 10660
rect 6870 10657 6876 10669
rect 6757 10629 6876 10657
rect 6757 10626 6769 10629
rect 6711 10620 6769 10626
rect 6870 10617 6876 10629
rect 6928 10617 6934 10669
rect 6711 10352 6769 10358
rect 6711 10318 6723 10352
rect 6757 10349 6769 10352
rect 6870 10349 6876 10361
rect 6757 10321 6876 10349
rect 6757 10318 6769 10321
rect 6711 10312 6769 10318
rect 6870 10309 6876 10321
rect 6928 10309 6934 10361
rect 6711 10148 6769 10154
rect 6711 10114 6723 10148
rect 6757 10145 6769 10148
rect 6870 10145 6876 10157
rect 6757 10117 6876 10145
rect 6757 10114 6769 10117
rect 6711 10108 6769 10114
rect 6870 10105 6876 10117
rect 6928 10105 6934 10157
rect 6711 9944 6769 9950
rect 6711 9910 6723 9944
rect 6757 9941 6769 9944
rect 6870 9941 6876 9953
rect 6757 9913 6876 9941
rect 6757 9910 6769 9913
rect 6711 9904 6769 9910
rect 6870 9901 6876 9913
rect 6928 9901 6934 9953
rect 6711 9740 6769 9746
rect 6711 9706 6723 9740
rect 6757 9737 6769 9740
rect 6870 9737 6876 9749
rect 6757 9709 6876 9737
rect 6757 9706 6769 9709
rect 6711 9700 6769 9706
rect 6870 9697 6876 9709
rect 6928 9697 6934 9749
rect 6711 9536 6769 9542
rect 6711 9502 6723 9536
rect 6757 9533 6769 9536
rect 6870 9533 6876 9545
rect 6757 9505 6876 9533
rect 6757 9502 6769 9505
rect 6711 9496 6769 9502
rect 6870 9493 6876 9505
rect 6928 9493 6934 9545
rect 6711 9332 6769 9338
rect 6711 9298 6723 9332
rect 6757 9329 6769 9332
rect 6870 9329 6876 9341
rect 6757 9301 6876 9329
rect 6757 9298 6769 9301
rect 6711 9292 6769 9298
rect 6870 9289 6876 9301
rect 6928 9289 6934 9341
rect 6711 9128 6769 9134
rect 6711 9094 6723 9128
rect 6757 9125 6769 9128
rect 6870 9125 6876 9137
rect 6757 9097 6876 9125
rect 6757 9094 6769 9097
rect 6711 9088 6769 9094
rect 6870 9085 6876 9097
rect 6928 9085 6934 9137
rect 6711 8924 6769 8930
rect 6711 8890 6723 8924
rect 6757 8921 6769 8924
rect 6870 8921 6876 8933
rect 6757 8893 6876 8921
rect 6757 8890 6769 8893
rect 6711 8884 6769 8890
rect 6870 8881 6876 8893
rect 6928 8881 6934 8933
rect 3321 8713 3327 8765
rect 3379 8713 3385 8765
rect 3943 8713 3949 8765
rect 4001 8713 4007 8765
rect 4741 8713 4747 8765
rect 4799 8713 4805 8765
rect 5989 8713 5995 8765
rect 6047 8713 6053 8765
rect 109 8290 115 8342
rect 167 8290 173 8342
rect 6912 8276 6918 8288
rect 5139 8248 6918 8276
rect 2149 7865 2155 7917
rect 2207 7865 2213 7917
rect 2219 7657 2225 7669
rect 2167 7629 2225 7657
rect 2219 7617 2225 7629
rect 2277 7617 2283 7669
rect 109 7338 115 7390
rect 167 7338 173 7390
rect 2149 6913 2155 6965
rect 2207 6913 2213 6965
rect 109 6301 115 6353
rect 167 6301 173 6353
rect 2149 5679 2155 5731
rect 2207 5679 2213 5731
rect 322 5520 328 5572
rect 380 5520 386 5572
rect 730 5520 736 5572
rect 788 5520 794 5572
rect 1138 5520 1144 5572
rect 1196 5520 1202 5572
rect 1546 5520 1552 5572
rect 1604 5520 1610 5572
rect 1954 5520 1960 5572
rect 2012 5520 2018 5572
rect 5139 5257 5167 8248
rect 6912 8236 6918 8248
rect 6970 8236 6976 8288
rect 6997 7845 7025 7894
rect 7201 7845 7229 7894
rect 7405 7845 7433 7894
rect 7609 7845 7637 7894
rect 7813 7845 7841 7894
rect 8017 7845 8045 7894
rect 8221 7845 8249 7894
rect 8425 7845 8453 7894
rect 8629 7845 8657 7894
rect 8833 7845 8861 7894
rect 9037 7845 9065 7894
rect 9241 7845 9269 7894
rect 9445 7845 9473 7894
rect 9649 7845 9677 7894
rect 9853 7845 9881 7894
rect 10057 7845 10085 7894
rect 10261 7845 10289 7894
rect 10465 7845 10493 7894
rect 10669 7845 10697 7894
rect 10873 7845 10901 7894
rect 11077 7845 11105 7894
rect 11281 7845 11309 7894
rect 11485 7845 11513 7894
rect 11689 7845 11717 7894
rect 11893 7845 11921 7894
rect 12097 7845 12125 7894
rect 12301 7845 12329 7894
rect 12505 7845 12533 7894
rect 12709 7845 12737 7894
rect 12913 7845 12941 7894
rect 13117 7845 13145 7894
rect 13321 7845 13349 7894
rect 13525 7845 13553 7894
rect 13729 7845 13757 7894
rect 13933 7845 13961 7894
rect 14137 7845 14165 7894
rect 14341 7845 14369 7894
rect 14545 7845 14573 7894
rect 14749 7845 14777 7894
rect 14953 7845 14981 7894
rect 15157 7845 15185 7894
rect 15361 7845 15389 7894
rect 15565 7845 15593 7894
rect 15769 7845 15797 7894
rect 15973 7845 16001 7894
rect 16177 7845 16205 7894
rect 16381 7845 16409 7894
rect 16585 7845 16613 7894
rect 16789 7845 16817 7894
rect 16993 7845 17021 7894
rect 17197 7845 17225 7894
rect 17401 7845 17429 7894
rect 17605 7845 17633 7894
rect 17809 7845 17837 7894
rect 18013 7845 18041 7894
rect 18217 7845 18245 7894
rect 18421 7845 18449 7894
rect 18625 7845 18653 7894
rect 18829 7845 18857 7894
rect 19033 7845 19061 7894
rect 19237 7845 19265 7894
rect 19441 7845 19469 7894
rect 19645 7845 19673 7894
rect 19849 7845 19877 7894
rect 6988 7833 7034 7845
rect 6988 7799 6994 7833
rect 7028 7799 7034 7833
rect 6988 7787 7034 7799
rect 7192 7833 7238 7845
rect 7192 7799 7198 7833
rect 7232 7799 7238 7833
rect 7192 7787 7238 7799
rect 7396 7833 7442 7845
rect 7396 7799 7402 7833
rect 7436 7799 7442 7833
rect 7396 7787 7442 7799
rect 7600 7833 7646 7845
rect 7600 7799 7606 7833
rect 7640 7799 7646 7833
rect 7600 7787 7646 7799
rect 7804 7833 7850 7845
rect 7804 7799 7810 7833
rect 7844 7799 7850 7833
rect 7804 7787 7850 7799
rect 8008 7833 8054 7845
rect 8008 7799 8014 7833
rect 8048 7799 8054 7833
rect 8008 7787 8054 7799
rect 8212 7833 8258 7845
rect 8212 7799 8218 7833
rect 8252 7799 8258 7833
rect 8212 7787 8258 7799
rect 8416 7833 8462 7845
rect 8416 7799 8422 7833
rect 8456 7799 8462 7833
rect 8416 7787 8462 7799
rect 8620 7833 8666 7845
rect 8620 7799 8626 7833
rect 8660 7799 8666 7833
rect 8620 7787 8666 7799
rect 8824 7833 8870 7845
rect 8824 7799 8830 7833
rect 8864 7799 8870 7833
rect 8824 7787 8870 7799
rect 9028 7833 9074 7845
rect 9028 7799 9034 7833
rect 9068 7799 9074 7833
rect 9028 7787 9074 7799
rect 9232 7833 9278 7845
rect 9232 7799 9238 7833
rect 9272 7799 9278 7833
rect 9232 7787 9278 7799
rect 9436 7833 9482 7845
rect 9436 7799 9442 7833
rect 9476 7799 9482 7833
rect 9436 7787 9482 7799
rect 9640 7833 9686 7845
rect 9640 7799 9646 7833
rect 9680 7799 9686 7833
rect 9640 7787 9686 7799
rect 9844 7833 9890 7845
rect 9844 7799 9850 7833
rect 9884 7799 9890 7833
rect 9844 7787 9890 7799
rect 10048 7833 10094 7845
rect 10048 7799 10054 7833
rect 10088 7799 10094 7833
rect 10048 7787 10094 7799
rect 10252 7833 10298 7845
rect 10252 7799 10258 7833
rect 10292 7799 10298 7833
rect 10252 7787 10298 7799
rect 10456 7833 10502 7845
rect 10456 7799 10462 7833
rect 10496 7799 10502 7833
rect 10456 7787 10502 7799
rect 10660 7833 10706 7845
rect 10660 7799 10666 7833
rect 10700 7799 10706 7833
rect 10660 7787 10706 7799
rect 10864 7833 10910 7845
rect 10864 7799 10870 7833
rect 10904 7799 10910 7833
rect 10864 7787 10910 7799
rect 11068 7833 11114 7845
rect 11068 7799 11074 7833
rect 11108 7799 11114 7833
rect 11068 7787 11114 7799
rect 11272 7833 11318 7845
rect 11272 7799 11278 7833
rect 11312 7799 11318 7833
rect 11272 7787 11318 7799
rect 11476 7833 11522 7845
rect 11476 7799 11482 7833
rect 11516 7799 11522 7833
rect 11476 7787 11522 7799
rect 11680 7833 11726 7845
rect 11680 7799 11686 7833
rect 11720 7799 11726 7833
rect 11680 7787 11726 7799
rect 11884 7833 11930 7845
rect 11884 7799 11890 7833
rect 11924 7799 11930 7833
rect 11884 7787 11930 7799
rect 12088 7833 12134 7845
rect 12088 7799 12094 7833
rect 12128 7799 12134 7833
rect 12088 7787 12134 7799
rect 12292 7833 12338 7845
rect 12292 7799 12298 7833
rect 12332 7799 12338 7833
rect 12292 7787 12338 7799
rect 12496 7833 12542 7845
rect 12496 7799 12502 7833
rect 12536 7799 12542 7833
rect 12496 7787 12542 7799
rect 12700 7833 12746 7845
rect 12700 7799 12706 7833
rect 12740 7799 12746 7833
rect 12700 7787 12746 7799
rect 12904 7833 12950 7845
rect 12904 7799 12910 7833
rect 12944 7799 12950 7833
rect 12904 7787 12950 7799
rect 13108 7833 13154 7845
rect 13108 7799 13114 7833
rect 13148 7799 13154 7833
rect 13108 7787 13154 7799
rect 13312 7833 13358 7845
rect 13312 7799 13318 7833
rect 13352 7799 13358 7833
rect 13312 7787 13358 7799
rect 13516 7833 13562 7845
rect 13516 7799 13522 7833
rect 13556 7799 13562 7833
rect 13516 7787 13562 7799
rect 13720 7833 13766 7845
rect 13720 7799 13726 7833
rect 13760 7799 13766 7833
rect 13720 7787 13766 7799
rect 13924 7833 13970 7845
rect 13924 7799 13930 7833
rect 13964 7799 13970 7833
rect 13924 7787 13970 7799
rect 14128 7833 14174 7845
rect 14128 7799 14134 7833
rect 14168 7799 14174 7833
rect 14128 7787 14174 7799
rect 14332 7833 14378 7845
rect 14332 7799 14338 7833
rect 14372 7799 14378 7833
rect 14332 7787 14378 7799
rect 14536 7833 14582 7845
rect 14536 7799 14542 7833
rect 14576 7799 14582 7833
rect 14536 7787 14582 7799
rect 14740 7833 14786 7845
rect 14740 7799 14746 7833
rect 14780 7799 14786 7833
rect 14740 7787 14786 7799
rect 14944 7833 14990 7845
rect 14944 7799 14950 7833
rect 14984 7799 14990 7833
rect 14944 7787 14990 7799
rect 15148 7833 15194 7845
rect 15148 7799 15154 7833
rect 15188 7799 15194 7833
rect 15148 7787 15194 7799
rect 15352 7833 15398 7845
rect 15352 7799 15358 7833
rect 15392 7799 15398 7833
rect 15352 7787 15398 7799
rect 15556 7833 15602 7845
rect 15556 7799 15562 7833
rect 15596 7799 15602 7833
rect 15556 7787 15602 7799
rect 15760 7833 15806 7845
rect 15760 7799 15766 7833
rect 15800 7799 15806 7833
rect 15760 7787 15806 7799
rect 15964 7833 16010 7845
rect 15964 7799 15970 7833
rect 16004 7799 16010 7833
rect 15964 7787 16010 7799
rect 16168 7833 16214 7845
rect 16168 7799 16174 7833
rect 16208 7799 16214 7833
rect 16168 7787 16214 7799
rect 16372 7833 16418 7845
rect 16372 7799 16378 7833
rect 16412 7799 16418 7833
rect 16372 7787 16418 7799
rect 16576 7833 16622 7845
rect 16576 7799 16582 7833
rect 16616 7799 16622 7833
rect 16576 7787 16622 7799
rect 16780 7833 16826 7845
rect 16780 7799 16786 7833
rect 16820 7799 16826 7833
rect 16780 7787 16826 7799
rect 16984 7833 17030 7845
rect 16984 7799 16990 7833
rect 17024 7799 17030 7833
rect 16984 7787 17030 7799
rect 17188 7833 17234 7845
rect 17188 7799 17194 7833
rect 17228 7799 17234 7833
rect 17188 7787 17234 7799
rect 17392 7833 17438 7845
rect 17392 7799 17398 7833
rect 17432 7799 17438 7833
rect 17392 7787 17438 7799
rect 17596 7833 17642 7845
rect 17596 7799 17602 7833
rect 17636 7799 17642 7833
rect 17596 7787 17642 7799
rect 17800 7833 17846 7845
rect 17800 7799 17806 7833
rect 17840 7799 17846 7833
rect 17800 7787 17846 7799
rect 18004 7833 18050 7845
rect 18004 7799 18010 7833
rect 18044 7799 18050 7833
rect 18004 7787 18050 7799
rect 18208 7833 18254 7845
rect 18208 7799 18214 7833
rect 18248 7799 18254 7833
rect 18208 7787 18254 7799
rect 18412 7833 18458 7845
rect 18412 7799 18418 7833
rect 18452 7799 18458 7833
rect 18412 7787 18458 7799
rect 18616 7833 18662 7845
rect 18616 7799 18622 7833
rect 18656 7799 18662 7833
rect 18616 7787 18662 7799
rect 18820 7833 18866 7845
rect 18820 7799 18826 7833
rect 18860 7799 18866 7833
rect 18820 7787 18866 7799
rect 19024 7833 19070 7845
rect 19024 7799 19030 7833
rect 19064 7799 19070 7833
rect 19024 7787 19070 7799
rect 19228 7833 19274 7845
rect 19228 7799 19234 7833
rect 19268 7799 19274 7833
rect 19228 7787 19274 7799
rect 19432 7833 19478 7845
rect 19432 7799 19438 7833
rect 19472 7799 19478 7833
rect 19432 7787 19478 7799
rect 19636 7833 19682 7845
rect 19636 7799 19642 7833
rect 19676 7799 19682 7833
rect 19636 7787 19682 7799
rect 19840 7833 19886 7845
rect 19840 7799 19846 7833
rect 19880 7799 19886 7833
rect 19840 7787 19886 7799
rect 6859 7198 6865 7250
rect 6917 7198 6923 7250
rect 19915 7198 19921 7250
rect 19973 7198 19979 7250
rect 6859 6282 6865 6334
rect 6917 6282 6923 6334
rect 19915 6282 19921 6334
rect 19973 6282 19979 6334
rect 6988 6238 7034 6250
rect 6988 6204 6994 6238
rect 7028 6204 7034 6238
rect 6988 6192 7034 6204
rect 7192 6238 7238 6250
rect 7192 6204 7198 6238
rect 7232 6204 7238 6238
rect 7192 6192 7238 6204
rect 7396 6238 7442 6250
rect 7396 6204 7402 6238
rect 7436 6204 7442 6238
rect 7396 6192 7442 6204
rect 7600 6238 7646 6250
rect 7600 6204 7606 6238
rect 7640 6204 7646 6238
rect 7600 6192 7646 6204
rect 7804 6238 7850 6250
rect 7804 6204 7810 6238
rect 7844 6204 7850 6238
rect 7804 6192 7850 6204
rect 8008 6238 8054 6250
rect 8008 6204 8014 6238
rect 8048 6204 8054 6238
rect 8008 6192 8054 6204
rect 8212 6238 8258 6250
rect 8212 6204 8218 6238
rect 8252 6204 8258 6238
rect 8212 6192 8258 6204
rect 8416 6238 8462 6250
rect 8416 6204 8422 6238
rect 8456 6204 8462 6238
rect 8416 6192 8462 6204
rect 8620 6238 8666 6250
rect 8620 6204 8626 6238
rect 8660 6204 8666 6238
rect 8620 6192 8666 6204
rect 8824 6238 8870 6250
rect 8824 6204 8830 6238
rect 8864 6204 8870 6238
rect 8824 6192 8870 6204
rect 9028 6238 9074 6250
rect 9028 6204 9034 6238
rect 9068 6204 9074 6238
rect 9028 6192 9074 6204
rect 9232 6238 9278 6250
rect 9232 6204 9238 6238
rect 9272 6204 9278 6238
rect 9232 6192 9278 6204
rect 9436 6238 9482 6250
rect 9436 6204 9442 6238
rect 9476 6204 9482 6238
rect 9436 6192 9482 6204
rect 9640 6238 9686 6250
rect 9640 6204 9646 6238
rect 9680 6204 9686 6238
rect 9640 6192 9686 6204
rect 9844 6238 9890 6250
rect 9844 6204 9850 6238
rect 9884 6204 9890 6238
rect 9844 6192 9890 6204
rect 10048 6238 10094 6250
rect 10048 6204 10054 6238
rect 10088 6204 10094 6238
rect 10048 6192 10094 6204
rect 10252 6238 10298 6250
rect 10252 6204 10258 6238
rect 10292 6204 10298 6238
rect 10252 6192 10298 6204
rect 10456 6238 10502 6250
rect 10456 6204 10462 6238
rect 10496 6204 10502 6238
rect 10456 6192 10502 6204
rect 10660 6238 10706 6250
rect 10660 6204 10666 6238
rect 10700 6204 10706 6238
rect 10660 6192 10706 6204
rect 10864 6238 10910 6250
rect 10864 6204 10870 6238
rect 10904 6204 10910 6238
rect 10864 6192 10910 6204
rect 11068 6238 11114 6250
rect 11068 6204 11074 6238
rect 11108 6204 11114 6238
rect 11068 6192 11114 6204
rect 11272 6238 11318 6250
rect 11272 6204 11278 6238
rect 11312 6204 11318 6238
rect 11272 6192 11318 6204
rect 11476 6238 11522 6250
rect 11476 6204 11482 6238
rect 11516 6204 11522 6238
rect 11476 6192 11522 6204
rect 11680 6238 11726 6250
rect 11680 6204 11686 6238
rect 11720 6204 11726 6238
rect 11680 6192 11726 6204
rect 11884 6238 11930 6250
rect 11884 6204 11890 6238
rect 11924 6204 11930 6238
rect 11884 6192 11930 6204
rect 12088 6238 12134 6250
rect 12088 6204 12094 6238
rect 12128 6204 12134 6238
rect 12088 6192 12134 6204
rect 12292 6238 12338 6250
rect 12292 6204 12298 6238
rect 12332 6204 12338 6238
rect 12292 6192 12338 6204
rect 12496 6238 12542 6250
rect 12496 6204 12502 6238
rect 12536 6204 12542 6238
rect 12496 6192 12542 6204
rect 12700 6238 12746 6250
rect 12700 6204 12706 6238
rect 12740 6204 12746 6238
rect 12700 6192 12746 6204
rect 12904 6238 12950 6250
rect 12904 6204 12910 6238
rect 12944 6204 12950 6238
rect 12904 6192 12950 6204
rect 13108 6238 13154 6250
rect 13108 6204 13114 6238
rect 13148 6204 13154 6238
rect 13108 6192 13154 6204
rect 13312 6238 13358 6250
rect 13312 6204 13318 6238
rect 13352 6204 13358 6238
rect 13312 6192 13358 6204
rect 13516 6238 13562 6250
rect 13516 6204 13522 6238
rect 13556 6204 13562 6238
rect 13516 6192 13562 6204
rect 13720 6238 13766 6250
rect 13720 6204 13726 6238
rect 13760 6204 13766 6238
rect 13720 6192 13766 6204
rect 13924 6238 13970 6250
rect 13924 6204 13930 6238
rect 13964 6204 13970 6238
rect 13924 6192 13970 6204
rect 14128 6238 14174 6250
rect 14128 6204 14134 6238
rect 14168 6204 14174 6238
rect 14128 6192 14174 6204
rect 14332 6238 14378 6250
rect 14332 6204 14338 6238
rect 14372 6204 14378 6238
rect 14332 6192 14378 6204
rect 14536 6238 14582 6250
rect 14536 6204 14542 6238
rect 14576 6204 14582 6238
rect 14536 6192 14582 6204
rect 14740 6238 14786 6250
rect 14740 6204 14746 6238
rect 14780 6204 14786 6238
rect 14740 6192 14786 6204
rect 14944 6238 14990 6250
rect 14944 6204 14950 6238
rect 14984 6204 14990 6238
rect 14944 6192 14990 6204
rect 15148 6238 15194 6250
rect 15148 6204 15154 6238
rect 15188 6204 15194 6238
rect 15148 6192 15194 6204
rect 15352 6238 15398 6250
rect 15352 6204 15358 6238
rect 15392 6204 15398 6238
rect 15352 6192 15398 6204
rect 15556 6238 15602 6250
rect 15556 6204 15562 6238
rect 15596 6204 15602 6238
rect 15556 6192 15602 6204
rect 15760 6238 15806 6250
rect 15760 6204 15766 6238
rect 15800 6204 15806 6238
rect 15760 6192 15806 6204
rect 15964 6238 16010 6250
rect 15964 6204 15970 6238
rect 16004 6204 16010 6238
rect 15964 6192 16010 6204
rect 16168 6238 16214 6250
rect 16168 6204 16174 6238
rect 16208 6204 16214 6238
rect 16168 6192 16214 6204
rect 16372 6238 16418 6250
rect 16372 6204 16378 6238
rect 16412 6204 16418 6238
rect 16372 6192 16418 6204
rect 16576 6238 16622 6250
rect 16576 6204 16582 6238
rect 16616 6204 16622 6238
rect 16576 6192 16622 6204
rect 16780 6238 16826 6250
rect 16780 6204 16786 6238
rect 16820 6204 16826 6238
rect 16780 6192 16826 6204
rect 16984 6238 17030 6250
rect 16984 6204 16990 6238
rect 17024 6204 17030 6238
rect 16984 6192 17030 6204
rect 17188 6238 17234 6250
rect 17188 6204 17194 6238
rect 17228 6204 17234 6238
rect 17188 6192 17234 6204
rect 17392 6238 17438 6250
rect 17392 6204 17398 6238
rect 17432 6204 17438 6238
rect 17392 6192 17438 6204
rect 17596 6238 17642 6250
rect 17596 6204 17602 6238
rect 17636 6204 17642 6238
rect 17596 6192 17642 6204
rect 17800 6238 17846 6250
rect 17800 6204 17806 6238
rect 17840 6204 17846 6238
rect 17800 6192 17846 6204
rect 18004 6238 18050 6250
rect 18004 6204 18010 6238
rect 18044 6204 18050 6238
rect 18004 6192 18050 6204
rect 18208 6238 18254 6250
rect 18208 6204 18214 6238
rect 18248 6204 18254 6238
rect 18208 6192 18254 6204
rect 18412 6238 18458 6250
rect 18412 6204 18418 6238
rect 18452 6204 18458 6238
rect 18412 6192 18458 6204
rect 18616 6238 18662 6250
rect 18616 6204 18622 6238
rect 18656 6204 18662 6238
rect 18616 6192 18662 6204
rect 18820 6238 18866 6250
rect 18820 6204 18826 6238
rect 18860 6204 18866 6238
rect 18820 6192 18866 6204
rect 19024 6238 19070 6250
rect 19024 6204 19030 6238
rect 19064 6204 19070 6238
rect 19024 6192 19070 6204
rect 19228 6238 19274 6250
rect 19228 6204 19234 6238
rect 19268 6204 19274 6238
rect 19228 6192 19274 6204
rect 19432 6238 19478 6250
rect 19432 6204 19438 6238
rect 19472 6204 19478 6238
rect 19432 6192 19478 6204
rect 19636 6238 19682 6250
rect 19636 6204 19642 6238
rect 19676 6204 19682 6238
rect 19636 6192 19682 6204
rect 19840 6238 19886 6250
rect 19840 6204 19846 6238
rect 19880 6204 19886 6238
rect 19840 6192 19886 6204
rect 6997 5686 7025 6192
rect 7201 5686 7229 6192
rect 7405 5686 7433 6192
rect 7609 5686 7637 6192
rect 7813 5686 7841 6192
rect 8017 5686 8045 6192
rect 8221 5686 8249 6192
rect 8425 5686 8453 6192
rect 8629 5686 8657 6192
rect 8833 5686 8861 6192
rect 9037 5686 9065 6192
rect 9241 5686 9269 6192
rect 9445 5686 9473 6192
rect 9649 5686 9677 6192
rect 9853 5686 9881 6192
rect 10057 5686 10085 6192
rect 10261 5686 10289 6192
rect 10465 5686 10493 6192
rect 10669 5686 10697 6192
rect 10873 5686 10901 6192
rect 11077 5686 11105 6192
rect 11281 5686 11309 6192
rect 11485 5686 11513 6192
rect 11689 5686 11717 6192
rect 11893 5686 11921 6192
rect 12097 5686 12125 6192
rect 12301 5686 12329 6192
rect 12505 5686 12533 6192
rect 12709 5686 12737 6192
rect 12913 5686 12941 6192
rect 13117 5686 13145 6192
rect 13321 5686 13349 6192
rect 13525 5686 13553 6192
rect 13729 5686 13757 6192
rect 13933 5686 13961 6192
rect 14137 5686 14165 6192
rect 14341 5686 14369 6192
rect 14545 5686 14573 6192
rect 14749 5686 14777 6192
rect 14953 5686 14981 6192
rect 15157 5686 15185 6192
rect 15361 5686 15389 6192
rect 15565 5686 15593 6192
rect 15769 5686 15797 6192
rect 15973 5686 16001 6192
rect 16177 5686 16205 6192
rect 16381 5686 16409 6192
rect 16585 5686 16613 6192
rect 16789 5686 16817 6192
rect 16993 5686 17021 6192
rect 17197 5686 17225 6192
rect 17401 5686 17429 6192
rect 17605 5686 17633 6192
rect 17809 5686 17837 6192
rect 18013 5686 18041 6192
rect 18217 5686 18245 6192
rect 18421 5686 18449 6192
rect 18625 5686 18653 6192
rect 18829 5686 18857 6192
rect 19033 5686 19061 6192
rect 19237 5686 19265 6192
rect 19441 5686 19469 6192
rect 19645 5686 19673 6192
rect 19849 5686 19877 6192
rect 3042 5229 5167 5257
rect 2501 4092 2559 4098
rect 2501 4058 2513 4092
rect 2547 4089 2559 4092
rect 3042 4089 3070 5229
rect 5767 4960 5773 5012
rect 5825 4960 5831 5012
rect 6389 4960 6395 5012
rect 6447 4960 6453 5012
rect 6708 4840 6714 4892
rect 6766 4840 6772 4892
rect 6708 4636 6714 4688
rect 6766 4636 6772 4688
rect 6708 4432 6714 4484
rect 6766 4432 6772 4484
rect 6708 4228 6714 4280
rect 6766 4228 6772 4280
rect 2547 4061 3070 4089
rect 2547 4058 2559 4061
rect 2501 4052 2559 4058
rect 3042 2188 3070 4061
rect 6708 4024 6714 4076
rect 6766 4024 6772 4076
rect 6708 3820 6714 3872
rect 6766 3820 6772 3872
rect 6708 3616 6714 3668
rect 6766 3616 6772 3668
rect 6708 3412 6714 3464
rect 6766 3412 6772 3464
rect 5767 3244 5773 3296
rect 5825 3244 5831 3296
rect 6389 3244 6395 3296
rect 6447 3244 6453 3296
rect 6979 3194 6985 3246
rect 7037 3194 7043 3246
rect 8611 3194 8617 3246
rect 8669 3194 8675 3246
rect 10243 3194 10249 3246
rect 10301 3194 10307 3246
rect 11875 3194 11881 3246
rect 11933 3194 11939 3246
rect 13507 3194 13513 3246
rect 13565 3194 13571 3246
rect 15139 3194 15145 3246
rect 15197 3194 15203 3246
rect 16771 3194 16777 3246
rect 16829 3194 16835 3246
rect 18403 3194 18409 3246
rect 18461 3194 18467 3246
rect 3371 2821 3377 2873
rect 3429 2821 3435 2873
rect 10701 2717 10707 2769
rect 10759 2757 10765 2769
rect 18403 2757 18409 2769
rect 10759 2729 18409 2757
rect 10759 2717 10765 2729
rect 18403 2717 18409 2729
rect 18461 2717 18467 2769
rect 10085 2615 10091 2667
rect 10143 2655 10149 2667
rect 15139 2655 15145 2667
rect 10143 2627 15145 2655
rect 10143 2615 10149 2627
rect 15139 2615 15145 2627
rect 15197 2615 15203 2667
rect 9777 2513 9783 2565
rect 9835 2553 9841 2565
rect 13507 2553 13513 2565
rect 9835 2525 13513 2553
rect 9835 2513 9841 2525
rect 13507 2513 13513 2525
rect 13565 2513 13571 2565
rect 4595 2396 4601 2448
rect 4653 2396 4659 2448
rect 8611 2411 8617 2463
rect 8669 2451 8675 2463
rect 8853 2451 8859 2463
rect 8669 2423 8859 2451
rect 8669 2411 8675 2423
rect 8853 2411 8859 2423
rect 8911 2411 8917 2463
rect 9469 2411 9475 2463
rect 9527 2451 9533 2463
rect 11875 2451 11881 2463
rect 9527 2423 11881 2451
rect 9527 2411 9533 2423
rect 11875 2411 11881 2423
rect 11933 2411 11939 2463
rect 6979 2309 6985 2361
rect 7037 2349 7043 2361
rect 8545 2349 8551 2361
rect 7037 2321 8551 2349
rect 7037 2309 7043 2321
rect 8545 2309 8551 2321
rect 8603 2309 8609 2361
rect 9161 2309 9167 2361
rect 9219 2349 9225 2361
rect 10243 2349 10249 2361
rect 9219 2321 10249 2349
rect 9219 2309 9225 2321
rect 10243 2309 10249 2321
rect 10301 2309 10307 2361
rect 10393 2309 10399 2361
rect 10451 2349 10457 2361
rect 16771 2349 16777 2361
rect 10451 2321 16777 2349
rect 10451 2309 10457 2321
rect 16771 2309 16777 2321
rect 16829 2309 16835 2361
rect 3042 2160 4001 2188
rect 8545 2086 8551 2138
rect 8603 2086 8609 2138
rect 8853 2086 8859 2138
rect 8911 2086 8917 2138
rect 9161 2086 9167 2138
rect 9219 2086 9225 2138
rect 9469 2086 9475 2138
rect 9527 2086 9533 2138
rect 9777 2086 9783 2138
rect 9835 2086 9841 2138
rect 10085 2086 10091 2138
rect 10143 2086 10149 2138
rect 10393 2086 10399 2138
rect 10451 2086 10457 2138
rect 10701 2086 10707 2138
rect 10759 2086 10765 2138
rect 3371 1869 3377 1921
rect 3429 1869 3435 1921
rect 8377 1816 8383 1868
rect 8435 1816 8441 1868
rect 10821 1816 10827 1868
rect 10879 1816 10885 1868
rect 4595 1444 4601 1496
rect 4653 1444 4659 1496
rect 475 1384 481 1436
rect 533 1384 539 1436
rect 2022 1322 2028 1374
rect 2080 1322 2086 1374
rect 8377 900 8383 952
rect 8435 900 8441 952
rect 10821 900 10827 952
rect 10879 900 10885 952
rect 3371 832 3377 884
rect 3429 832 3435 884
rect 8551 433 8603 439
rect 2535 377 2541 429
rect 2593 377 2599 429
rect 8551 375 8603 381
rect 8859 433 8911 439
rect 8859 375 8911 381
rect 9167 433 9219 439
rect 9167 375 9219 381
rect 9475 433 9527 439
rect 9475 375 9527 381
rect 9783 433 9835 439
rect 9783 375 9835 381
rect 10091 433 10143 439
rect 10091 375 10143 381
rect 10399 433 10451 439
rect 10399 375 10451 381
rect 10707 433 10759 439
rect 10707 375 10759 381
rect 4595 210 4601 262
rect 4653 210 4659 262
rect 3584 51 3590 103
rect 3642 51 3648 103
rect 3992 51 3998 103
rect 4050 51 4056 103
rect 4400 51 4406 103
rect 4458 51 4464 103
<< via1 >>
rect 6971 15848 7023 15900
rect 19851 15848 19903 15900
rect 3327 15637 3379 15689
rect 3949 15637 4001 15689
rect 4747 15637 4799 15689
rect 5995 15637 6047 15689
rect 6876 15517 6928 15569
rect 6876 15313 6928 15365
rect 6876 15109 6928 15161
rect 6876 14905 6928 14957
rect 6876 14701 6928 14753
rect 6876 14497 6928 14549
rect 6876 14293 6928 14345
rect 6876 14089 6928 14141
rect 6876 13781 6928 13833
rect 6876 13577 6928 13629
rect 6876 13373 6928 13425
rect 6876 13169 6928 13221
rect 6876 12965 6928 13017
rect 6876 12761 6928 12813
rect 6876 12557 6928 12609
rect 6876 12353 6928 12405
rect 6876 12045 6928 12097
rect 6876 11841 6928 11893
rect 6876 11637 6928 11689
rect 6876 11433 6928 11485
rect 6876 11229 6928 11281
rect 6876 11025 6928 11077
rect 6876 10821 6928 10873
rect 6876 10617 6928 10669
rect 6876 10309 6928 10361
rect 6876 10105 6928 10157
rect 6876 9901 6928 9953
rect 6876 9697 6928 9749
rect 6876 9493 6928 9545
rect 6876 9289 6928 9341
rect 6876 9085 6928 9137
rect 6876 8881 6928 8933
rect 3327 8713 3379 8765
rect 3949 8713 4001 8765
rect 4747 8713 4799 8765
rect 5995 8713 6047 8765
rect 115 8290 167 8342
rect 2155 7865 2207 7917
rect 2225 7617 2277 7669
rect 115 7338 167 7390
rect 2155 6913 2207 6965
rect 115 6301 167 6353
rect 2155 5679 2207 5731
rect 328 5563 380 5572
rect 328 5529 337 5563
rect 337 5529 371 5563
rect 371 5529 380 5563
rect 328 5520 380 5529
rect 736 5563 788 5572
rect 736 5529 745 5563
rect 745 5529 779 5563
rect 779 5529 788 5563
rect 736 5520 788 5529
rect 1144 5563 1196 5572
rect 1144 5529 1153 5563
rect 1153 5529 1187 5563
rect 1187 5529 1196 5563
rect 1144 5520 1196 5529
rect 1552 5563 1604 5572
rect 1552 5529 1561 5563
rect 1561 5529 1595 5563
rect 1595 5529 1604 5563
rect 1552 5520 1604 5529
rect 1960 5563 2012 5572
rect 1960 5529 1969 5563
rect 1969 5529 2003 5563
rect 2003 5529 2012 5563
rect 1960 5520 2012 5529
rect 6918 8236 6970 8288
rect 6865 7198 6917 7250
rect 19921 7198 19973 7250
rect 6865 6282 6917 6334
rect 19921 6282 19973 6334
rect 5773 4960 5825 5012
rect 6395 4960 6447 5012
rect 6714 4883 6766 4892
rect 6714 4849 6723 4883
rect 6723 4849 6757 4883
rect 6757 4849 6766 4883
rect 6714 4840 6766 4849
rect 6714 4679 6766 4688
rect 6714 4645 6723 4679
rect 6723 4645 6757 4679
rect 6757 4645 6766 4679
rect 6714 4636 6766 4645
rect 6714 4475 6766 4484
rect 6714 4441 6723 4475
rect 6723 4441 6757 4475
rect 6757 4441 6766 4475
rect 6714 4432 6766 4441
rect 6714 4271 6766 4280
rect 6714 4237 6723 4271
rect 6723 4237 6757 4271
rect 6757 4237 6766 4271
rect 6714 4228 6766 4237
rect 6714 4067 6766 4076
rect 6714 4033 6723 4067
rect 6723 4033 6757 4067
rect 6757 4033 6766 4067
rect 6714 4024 6766 4033
rect 6714 3863 6766 3872
rect 6714 3829 6723 3863
rect 6723 3829 6757 3863
rect 6757 3829 6766 3863
rect 6714 3820 6766 3829
rect 6714 3659 6766 3668
rect 6714 3625 6723 3659
rect 6723 3625 6757 3659
rect 6757 3625 6766 3659
rect 6714 3616 6766 3625
rect 6714 3455 6766 3464
rect 6714 3421 6723 3455
rect 6723 3421 6757 3455
rect 6757 3421 6766 3455
rect 6714 3412 6766 3421
rect 5773 3244 5825 3296
rect 6395 3244 6447 3296
rect 6985 3194 7037 3246
rect 8617 3194 8669 3246
rect 10249 3194 10301 3246
rect 11881 3194 11933 3246
rect 13513 3194 13565 3246
rect 15145 3194 15197 3246
rect 16777 3194 16829 3246
rect 18409 3194 18461 3246
rect 3377 2821 3429 2873
rect 10707 2717 10759 2769
rect 18409 2717 18461 2769
rect 10091 2615 10143 2667
rect 15145 2615 15197 2667
rect 9783 2513 9835 2565
rect 13513 2513 13565 2565
rect 4601 2396 4653 2448
rect 8617 2411 8669 2463
rect 8859 2411 8911 2463
rect 9475 2411 9527 2463
rect 11881 2411 11933 2463
rect 6985 2309 7037 2361
rect 8551 2309 8603 2361
rect 9167 2309 9219 2361
rect 10249 2309 10301 2361
rect 10399 2309 10451 2361
rect 16777 2309 16829 2361
rect 8551 2129 8603 2138
rect 8551 2095 8560 2129
rect 8560 2095 8594 2129
rect 8594 2095 8603 2129
rect 8551 2086 8603 2095
rect 8859 2129 8911 2138
rect 8859 2095 8868 2129
rect 8868 2095 8902 2129
rect 8902 2095 8911 2129
rect 8859 2086 8911 2095
rect 9167 2129 9219 2138
rect 9167 2095 9176 2129
rect 9176 2095 9210 2129
rect 9210 2095 9219 2129
rect 9167 2086 9219 2095
rect 9475 2129 9527 2138
rect 9475 2095 9484 2129
rect 9484 2095 9518 2129
rect 9518 2095 9527 2129
rect 9475 2086 9527 2095
rect 9783 2129 9835 2138
rect 9783 2095 9792 2129
rect 9792 2095 9826 2129
rect 9826 2095 9835 2129
rect 9783 2086 9835 2095
rect 10091 2129 10143 2138
rect 10091 2095 10100 2129
rect 10100 2095 10134 2129
rect 10134 2095 10143 2129
rect 10091 2086 10143 2095
rect 10399 2129 10451 2138
rect 10399 2095 10408 2129
rect 10408 2095 10442 2129
rect 10442 2095 10451 2129
rect 10399 2086 10451 2095
rect 10707 2129 10759 2138
rect 10707 2095 10716 2129
rect 10716 2095 10750 2129
rect 10750 2095 10759 2129
rect 10707 2086 10759 2095
rect 3377 1869 3429 1921
rect 8383 1816 8435 1868
rect 10827 1816 10879 1868
rect 4601 1444 4653 1496
rect 481 1427 533 1436
rect 481 1393 490 1427
rect 490 1393 524 1427
rect 524 1393 533 1427
rect 481 1384 533 1393
rect 2028 1365 2080 1374
rect 2028 1331 2037 1365
rect 2037 1331 2071 1365
rect 2071 1331 2080 1365
rect 2028 1322 2080 1331
rect 8383 900 8435 952
rect 10827 900 10879 952
rect 3377 832 3429 884
rect 2541 420 2593 429
rect 2541 386 2550 420
rect 2550 386 2584 420
rect 2584 386 2593 420
rect 2541 377 2593 386
rect 8551 424 8603 433
rect 8551 390 8560 424
rect 8560 390 8594 424
rect 8594 390 8603 424
rect 8551 381 8603 390
rect 8859 424 8911 433
rect 8859 390 8868 424
rect 8868 390 8902 424
rect 8902 390 8911 424
rect 8859 381 8911 390
rect 9167 424 9219 433
rect 9167 390 9176 424
rect 9176 390 9210 424
rect 9210 390 9219 424
rect 9167 381 9219 390
rect 9475 424 9527 433
rect 9475 390 9484 424
rect 9484 390 9518 424
rect 9518 390 9527 424
rect 9475 381 9527 390
rect 9783 424 9835 433
rect 9783 390 9792 424
rect 9792 390 9826 424
rect 9826 390 9835 424
rect 9783 381 9835 390
rect 10091 424 10143 433
rect 10091 390 10100 424
rect 10100 390 10134 424
rect 10134 390 10143 424
rect 10091 381 10143 390
rect 10399 424 10451 433
rect 10399 390 10408 424
rect 10408 390 10442 424
rect 10442 390 10451 424
rect 10399 381 10451 390
rect 10707 424 10759 433
rect 10707 390 10716 424
rect 10716 390 10750 424
rect 10750 390 10759 424
rect 10707 381 10759 390
rect 4601 210 4653 262
rect 3590 94 3642 103
rect 3590 60 3599 94
rect 3599 60 3633 94
rect 3633 60 3642 94
rect 3590 51 3642 60
rect 3998 94 4050 103
rect 3998 60 4007 94
rect 4007 60 4041 94
rect 4041 60 4050 94
rect 3998 51 4050 60
rect 4406 94 4458 103
rect 4406 60 4415 94
rect 4415 60 4449 94
rect 4449 60 4458 94
rect 4406 51 4458 60
<< metal2 >>
rect 6969 15902 7025 15911
rect 6969 15837 7025 15846
rect 19849 15902 19905 15911
rect 19849 15837 19905 15846
rect 3325 15691 3381 15700
rect 3325 15626 3381 15635
rect 3947 15691 4003 15700
rect 3947 15626 4003 15635
rect 4745 15691 4801 15700
rect 4745 15626 4801 15635
rect 5993 15691 6049 15700
rect 5993 15626 6049 15635
rect 6876 15569 6928 15575
rect 6870 15522 6876 15565
rect 6928 15522 6934 15565
rect 6876 15511 6928 15517
rect 6876 15365 6928 15371
rect 6870 15318 6876 15361
rect 6928 15318 6934 15361
rect 6876 15307 6928 15313
rect 6876 15161 6928 15167
rect 6870 15114 6876 15157
rect 6928 15114 6934 15157
rect 6876 15103 6928 15109
rect 6876 14957 6928 14963
rect 6870 14910 6876 14953
rect 6928 14910 6934 14953
rect 6876 14899 6928 14905
rect 6876 14753 6928 14759
rect 6870 14706 6876 14749
rect 6928 14706 6934 14749
rect 6876 14695 6928 14701
rect 6876 14549 6928 14555
rect 6870 14502 6876 14545
rect 6928 14502 6934 14545
rect 6876 14491 6928 14497
rect 6876 14345 6928 14351
rect 6870 14298 6876 14341
rect 6928 14298 6934 14341
rect 6876 14287 6928 14293
rect 6876 14141 6928 14147
rect 6870 14094 6876 14137
rect 6928 14094 6934 14137
rect 6876 14083 6928 14089
rect 13518 13989 13574 13998
rect 13518 13924 13574 13933
rect 6876 13833 6928 13839
rect 6870 13786 6876 13829
rect 6928 13786 6934 13829
rect 6876 13775 6928 13781
rect 6876 13629 6928 13635
rect 6870 13582 6876 13625
rect 6928 13582 6934 13625
rect 6876 13571 6928 13577
rect 6876 13425 6928 13431
rect 6870 13378 6876 13421
rect 6928 13378 6934 13421
rect 6876 13367 6928 13373
rect 6876 13221 6928 13227
rect 6870 13174 6876 13217
rect 6928 13174 6934 13217
rect 6876 13163 6928 13169
rect 6876 13017 6928 13023
rect 6870 12970 6876 13013
rect 6928 12970 6934 13013
rect 6876 12959 6928 12965
rect 6876 12813 6928 12819
rect 6870 12766 6876 12809
rect 6928 12766 6934 12809
rect 6876 12755 6928 12761
rect 6876 12609 6928 12615
rect 6870 12562 6876 12605
rect 6928 12562 6934 12605
rect 6876 12551 6928 12557
rect 6876 12405 6928 12411
rect 6870 12358 6876 12401
rect 6928 12358 6934 12401
rect 6876 12347 6928 12353
rect 13518 12253 13574 12262
rect 13518 12188 13574 12197
rect 6876 12097 6928 12103
rect 6870 12050 6876 12093
rect 6928 12050 6934 12093
rect 6876 12039 6928 12045
rect 6876 11893 6928 11899
rect 6870 11846 6876 11889
rect 6928 11846 6934 11889
rect 6876 11835 6928 11841
rect 6876 11689 6928 11695
rect 6870 11642 6876 11685
rect 6928 11642 6934 11685
rect 6876 11631 6928 11637
rect 6876 11485 6928 11491
rect 6870 11438 6876 11481
rect 6928 11438 6934 11481
rect 6876 11427 6928 11433
rect 6876 11281 6928 11287
rect 6870 11234 6876 11277
rect 6928 11234 6934 11277
rect 6876 11223 6928 11229
rect 6876 11077 6928 11083
rect 6870 11030 6876 11073
rect 6928 11030 6934 11073
rect 6876 11019 6928 11025
rect 6876 10873 6928 10879
rect 6870 10826 6876 10869
rect 6928 10826 6934 10869
rect 6876 10815 6928 10821
rect 6876 10669 6928 10675
rect 6870 10622 6876 10665
rect 6928 10622 6934 10665
rect 6876 10611 6928 10617
rect 13518 10517 13574 10526
rect 13518 10452 13574 10461
rect 6876 10361 6928 10367
rect 6870 10314 6876 10357
rect 6928 10314 6934 10357
rect 6876 10303 6928 10309
rect 6876 10157 6928 10163
rect 6870 10110 6876 10153
rect 6928 10110 6934 10153
rect 6876 10099 6928 10105
rect 6876 9953 6928 9959
rect 6870 9906 6876 9949
rect 6928 9906 6934 9949
rect 6876 9895 6928 9901
rect 6876 9749 6928 9755
rect 6870 9702 6876 9745
rect 6928 9702 6934 9745
rect 6876 9691 6928 9697
rect 6876 9545 6928 9551
rect 6870 9498 6876 9541
rect 6928 9498 6934 9541
rect 6876 9487 6928 9493
rect 6876 9341 6928 9347
rect 6870 9294 6876 9337
rect 6928 9294 6934 9337
rect 6876 9283 6928 9289
rect 6876 9137 6928 9143
rect 6870 9090 6876 9133
rect 6928 9090 6934 9133
rect 6876 9079 6928 9085
rect 6876 8933 6928 8939
rect 6870 8886 6876 8929
rect 6928 8886 6934 8929
rect 6876 8875 6928 8881
rect 13518 8781 13574 8790
rect 3325 8767 3381 8776
rect 2237 8722 2721 8750
rect 113 8344 169 8353
rect 113 8279 169 8288
rect 2153 7919 2209 7928
rect 2153 7854 2209 7863
rect 2237 7675 2265 8722
rect 3061 8715 3117 8724
rect 3325 8702 3381 8711
rect 3947 8767 4003 8776
rect 3947 8702 4003 8711
rect 4745 8767 4801 8776
rect 4745 8702 4801 8711
rect 5993 8767 6049 8776
rect 13518 8716 13574 8725
rect 5993 8702 6049 8711
rect 3061 8650 3117 8659
rect 6918 8288 6970 8294
rect 6918 8230 6970 8236
rect 6867 7908 6923 7917
rect 6867 7843 6923 7852
rect 2225 7669 2277 7675
rect 2277 7629 3116 7657
rect 2225 7611 2277 7617
rect 113 7392 169 7401
rect 113 7327 169 7336
rect 2153 6967 2209 6976
rect 2153 6902 2209 6911
rect 113 6355 169 6364
rect 113 6290 169 6299
rect 2153 5733 2209 5742
rect 2153 5668 2209 5677
rect 326 5574 382 5583
rect 326 5509 382 5518
rect 734 5574 790 5583
rect 734 5509 790 5518
rect 1142 5574 1198 5583
rect 1142 5509 1198 5518
rect 1550 5574 1606 5583
rect 1550 5509 1606 5518
rect 1958 5574 2014 5583
rect 1958 5509 2014 5518
rect 479 1438 535 1447
rect 479 1373 535 1382
rect 2028 1374 2080 1380
rect 3088 1362 3116 7629
rect 6863 7252 6919 7261
rect 6863 7187 6919 7196
rect 19919 7252 19975 7261
rect 19919 7187 19975 7196
rect 6863 6336 6919 6345
rect 6863 6271 6919 6280
rect 19919 6336 19975 6345
rect 19919 6271 19975 6280
rect 13450 5834 13506 5843
rect 13450 5769 13506 5778
rect 5771 5014 5827 5023
rect 5771 4949 5827 4958
rect 6393 5014 6449 5023
rect 6393 4949 6449 4958
rect 6714 4892 6766 4898
rect 6766 4852 19973 4880
rect 6714 4834 6766 4840
rect 6714 4688 6766 4694
rect 6766 4648 19973 4676
rect 6714 4630 6766 4636
rect 6714 4484 6766 4490
rect 6766 4444 19973 4472
rect 6714 4426 6766 4432
rect 6714 4280 6766 4286
rect 6766 4240 19973 4268
rect 6714 4222 6766 4228
rect 6714 4076 6766 4082
rect 6766 4036 19973 4064
rect 6714 4018 6766 4024
rect 6714 3872 6766 3878
rect 6766 3832 19973 3860
rect 6714 3814 6766 3820
rect 6714 3668 6766 3674
rect 6766 3628 19973 3656
rect 6714 3610 6766 3616
rect 6714 3464 6766 3470
rect 6766 3424 19973 3452
rect 6714 3406 6766 3412
rect 5771 3298 5827 3307
rect 5507 3246 5563 3255
rect 5771 3233 5827 3242
rect 6393 3298 6449 3307
rect 6393 3233 6449 3242
rect 6985 3246 7037 3252
rect 5507 3181 5563 3190
rect 6985 3188 7037 3194
rect 8617 3246 8669 3252
rect 8617 3188 8669 3194
rect 10249 3246 10301 3252
rect 10249 3188 10301 3194
rect 11881 3246 11933 3252
rect 11881 3188 11933 3194
rect 13513 3246 13565 3252
rect 13513 3188 13565 3194
rect 15145 3246 15197 3252
rect 15145 3188 15197 3194
rect 16777 3246 16829 3252
rect 16777 3188 16829 3194
rect 18409 3246 18461 3252
rect 18409 3188 18461 3194
rect 3375 2875 3431 2884
rect 3375 2810 3431 2819
rect 4599 2450 4655 2459
rect 4599 2385 4655 2394
rect 6997 2367 7025 3188
rect 8629 2469 8657 3188
rect 10091 2667 10143 2673
rect 10091 2609 10143 2615
rect 9783 2565 9835 2571
rect 9783 2507 9835 2513
rect 8617 2463 8669 2469
rect 8617 2405 8669 2411
rect 8859 2463 8911 2469
rect 8859 2405 8911 2411
rect 9475 2463 9527 2469
rect 9475 2405 9527 2411
rect 6985 2361 7037 2367
rect 6985 2303 7037 2309
rect 8551 2361 8603 2367
rect 8551 2303 8603 2309
rect 8563 2144 8591 2303
rect 8871 2144 8899 2405
rect 9167 2361 9219 2367
rect 9167 2303 9219 2309
rect 9179 2144 9207 2303
rect 9487 2144 9515 2405
rect 9795 2144 9823 2507
rect 10103 2144 10131 2609
rect 10261 2367 10289 3188
rect 10707 2769 10759 2775
rect 10707 2711 10759 2717
rect 10249 2361 10301 2367
rect 10249 2303 10301 2309
rect 10399 2361 10451 2367
rect 10399 2303 10451 2309
rect 10411 2144 10439 2303
rect 10719 2144 10747 2711
rect 11893 2469 11921 3188
rect 13525 2571 13553 3188
rect 15157 2673 15185 3188
rect 15145 2667 15197 2673
rect 15145 2609 15197 2615
rect 13513 2565 13565 2571
rect 13513 2507 13565 2513
rect 11881 2463 11933 2469
rect 11881 2405 11933 2411
rect 16789 2367 16817 3188
rect 18421 2775 18449 3188
rect 18409 2769 18461 2775
rect 18409 2711 18461 2717
rect 16777 2361 16829 2367
rect 16777 2303 16829 2309
rect 8551 2138 8603 2144
rect 8551 2080 8603 2086
rect 8859 2138 8911 2144
rect 8859 2080 8911 2086
rect 9167 2138 9219 2144
rect 9167 2080 9219 2086
rect 9475 2138 9527 2144
rect 9475 2080 9527 2086
rect 9783 2138 9835 2144
rect 9783 2080 9835 2086
rect 10091 2138 10143 2144
rect 10091 2080 10143 2086
rect 10399 2138 10451 2144
rect 10399 2080 10451 2086
rect 10707 2138 10759 2144
rect 10707 2080 10759 2086
rect 3375 1923 3431 1932
rect 3375 1858 3431 1867
rect 8381 1870 8437 1879
rect 8381 1805 8437 1814
rect 10825 1870 10881 1879
rect 10825 1805 10881 1814
rect 4599 1498 4655 1507
rect 4599 1433 4655 1442
rect 2080 1334 3116 1362
rect 2028 1316 2080 1322
rect 8381 954 8437 963
rect 3375 886 3431 895
rect 8381 889 8437 898
rect 10825 954 10881 963
rect 10825 889 10881 898
rect 3375 821 3431 830
rect 2539 431 2595 440
rect 8540 379 8549 435
rect 8605 379 8614 435
rect 8848 379 8857 435
rect 8913 379 8922 435
rect 9156 379 9165 435
rect 9221 379 9230 435
rect 9464 379 9473 435
rect 9529 379 9538 435
rect 9772 379 9781 435
rect 9837 379 9846 435
rect 10080 379 10089 435
rect 10145 379 10154 435
rect 10388 379 10397 435
rect 10453 379 10462 435
rect 10696 379 10705 435
rect 10761 379 10770 435
rect 2539 366 2595 375
rect 4599 264 4655 273
rect 4599 199 4655 208
rect 3588 105 3644 114
rect 3588 40 3644 49
rect 3996 105 4052 114
rect 3996 40 4052 49
rect 4404 105 4460 114
rect 4404 40 4460 49
<< via2 >>
rect 6969 15900 7025 15902
rect 6969 15848 6971 15900
rect 6971 15848 7023 15900
rect 7023 15848 7025 15900
rect 6969 15846 7025 15848
rect 19849 15900 19905 15902
rect 19849 15848 19851 15900
rect 19851 15848 19903 15900
rect 19903 15848 19905 15900
rect 19849 15846 19905 15848
rect 3325 15689 3381 15691
rect 3325 15637 3327 15689
rect 3327 15637 3379 15689
rect 3379 15637 3381 15689
rect 3325 15635 3381 15637
rect 3947 15689 4003 15691
rect 3947 15637 3949 15689
rect 3949 15637 4001 15689
rect 4001 15637 4003 15689
rect 3947 15635 4003 15637
rect 4745 15689 4801 15691
rect 4745 15637 4747 15689
rect 4747 15637 4799 15689
rect 4799 15637 4801 15689
rect 4745 15635 4801 15637
rect 5993 15689 6049 15691
rect 5993 15637 5995 15689
rect 5995 15637 6047 15689
rect 6047 15637 6049 15689
rect 5993 15635 6049 15637
rect 13518 13933 13574 13989
rect 13518 12197 13574 12253
rect 13518 10461 13574 10517
rect 3325 8765 3381 8767
rect 113 8342 169 8344
rect 113 8290 115 8342
rect 115 8290 167 8342
rect 167 8290 169 8342
rect 113 8288 169 8290
rect 2153 7917 2209 7919
rect 2153 7865 2155 7917
rect 2155 7865 2207 7917
rect 2207 7865 2209 7917
rect 2153 7863 2209 7865
rect 3061 8659 3117 8715
rect 3325 8713 3327 8765
rect 3327 8713 3379 8765
rect 3379 8713 3381 8765
rect 3325 8711 3381 8713
rect 3947 8765 4003 8767
rect 3947 8713 3949 8765
rect 3949 8713 4001 8765
rect 4001 8713 4003 8765
rect 3947 8711 4003 8713
rect 4745 8765 4801 8767
rect 4745 8713 4747 8765
rect 4747 8713 4799 8765
rect 4799 8713 4801 8765
rect 4745 8711 4801 8713
rect 5993 8765 6049 8767
rect 5993 8713 5995 8765
rect 5995 8713 6047 8765
rect 6047 8713 6049 8765
rect 13518 8725 13574 8781
rect 5993 8711 6049 8713
rect 6867 7852 6923 7908
rect 113 7390 169 7392
rect 113 7338 115 7390
rect 115 7338 167 7390
rect 167 7338 169 7390
rect 113 7336 169 7338
rect 2153 6965 2209 6967
rect 2153 6913 2155 6965
rect 2155 6913 2207 6965
rect 2207 6913 2209 6965
rect 2153 6911 2209 6913
rect 113 6353 169 6355
rect 113 6301 115 6353
rect 115 6301 167 6353
rect 167 6301 169 6353
rect 113 6299 169 6301
rect 2153 5731 2209 5733
rect 2153 5679 2155 5731
rect 2155 5679 2207 5731
rect 2207 5679 2209 5731
rect 2153 5677 2209 5679
rect 326 5572 382 5574
rect 326 5520 328 5572
rect 328 5520 380 5572
rect 380 5520 382 5572
rect 326 5518 382 5520
rect 734 5572 790 5574
rect 734 5520 736 5572
rect 736 5520 788 5572
rect 788 5520 790 5572
rect 734 5518 790 5520
rect 1142 5572 1198 5574
rect 1142 5520 1144 5572
rect 1144 5520 1196 5572
rect 1196 5520 1198 5572
rect 1142 5518 1198 5520
rect 1550 5572 1606 5574
rect 1550 5520 1552 5572
rect 1552 5520 1604 5572
rect 1604 5520 1606 5572
rect 1550 5518 1606 5520
rect 1958 5572 2014 5574
rect 1958 5520 1960 5572
rect 1960 5520 2012 5572
rect 2012 5520 2014 5572
rect 1958 5518 2014 5520
rect 479 1436 535 1438
rect 479 1384 481 1436
rect 481 1384 533 1436
rect 533 1384 535 1436
rect 479 1382 535 1384
rect 6863 7250 6919 7252
rect 6863 7198 6865 7250
rect 6865 7198 6917 7250
rect 6917 7198 6919 7250
rect 6863 7196 6919 7198
rect 19919 7250 19975 7252
rect 19919 7198 19921 7250
rect 19921 7198 19973 7250
rect 19973 7198 19975 7250
rect 19919 7196 19975 7198
rect 6863 6334 6919 6336
rect 6863 6282 6865 6334
rect 6865 6282 6917 6334
rect 6917 6282 6919 6334
rect 6863 6280 6919 6282
rect 19919 6334 19975 6336
rect 19919 6282 19921 6334
rect 19921 6282 19973 6334
rect 19973 6282 19975 6334
rect 19919 6280 19975 6282
rect 13450 5778 13506 5834
rect 5771 5012 5827 5014
rect 5771 4960 5773 5012
rect 5773 4960 5825 5012
rect 5825 4960 5827 5012
rect 5771 4958 5827 4960
rect 6393 5012 6449 5014
rect 6393 4960 6395 5012
rect 6395 4960 6447 5012
rect 6447 4960 6449 5012
rect 6393 4958 6449 4960
rect 5771 3296 5827 3298
rect 5507 3190 5563 3246
rect 5771 3244 5773 3296
rect 5773 3244 5825 3296
rect 5825 3244 5827 3296
rect 5771 3242 5827 3244
rect 6393 3296 6449 3298
rect 6393 3244 6395 3296
rect 6395 3244 6447 3296
rect 6447 3244 6449 3296
rect 6393 3242 6449 3244
rect 3375 2873 3431 2875
rect 3375 2821 3377 2873
rect 3377 2821 3429 2873
rect 3429 2821 3431 2873
rect 3375 2819 3431 2821
rect 4599 2448 4655 2450
rect 4599 2396 4601 2448
rect 4601 2396 4653 2448
rect 4653 2396 4655 2448
rect 4599 2394 4655 2396
rect 3375 1921 3431 1923
rect 3375 1869 3377 1921
rect 3377 1869 3429 1921
rect 3429 1869 3431 1921
rect 3375 1867 3431 1869
rect 8381 1868 8437 1870
rect 8381 1816 8383 1868
rect 8383 1816 8435 1868
rect 8435 1816 8437 1868
rect 8381 1814 8437 1816
rect 10825 1868 10881 1870
rect 10825 1816 10827 1868
rect 10827 1816 10879 1868
rect 10879 1816 10881 1868
rect 10825 1814 10881 1816
rect 4599 1496 4655 1498
rect 4599 1444 4601 1496
rect 4601 1444 4653 1496
rect 4653 1444 4655 1496
rect 4599 1442 4655 1444
rect 8381 952 8437 954
rect 8381 900 8383 952
rect 8383 900 8435 952
rect 8435 900 8437 952
rect 8381 898 8437 900
rect 10825 952 10881 954
rect 10825 900 10827 952
rect 10827 900 10879 952
rect 10879 900 10881 952
rect 10825 898 10881 900
rect 3375 884 3431 886
rect 3375 832 3377 884
rect 3377 832 3429 884
rect 3429 832 3431 884
rect 3375 830 3431 832
rect 2539 429 2595 431
rect 2539 377 2541 429
rect 2541 377 2593 429
rect 2593 377 2595 429
rect 8549 433 8605 435
rect 8549 381 8551 433
rect 8551 381 8603 433
rect 8603 381 8605 433
rect 8549 379 8605 381
rect 8857 433 8913 435
rect 8857 381 8859 433
rect 8859 381 8911 433
rect 8911 381 8913 433
rect 8857 379 8913 381
rect 9165 433 9221 435
rect 9165 381 9167 433
rect 9167 381 9219 433
rect 9219 381 9221 433
rect 9165 379 9221 381
rect 9473 433 9529 435
rect 9473 381 9475 433
rect 9475 381 9527 433
rect 9527 381 9529 433
rect 9473 379 9529 381
rect 9781 433 9837 435
rect 9781 381 9783 433
rect 9783 381 9835 433
rect 9835 381 9837 433
rect 9781 379 9837 381
rect 10089 433 10145 435
rect 10089 381 10091 433
rect 10091 381 10143 433
rect 10143 381 10145 433
rect 10089 379 10145 381
rect 10397 433 10453 435
rect 10397 381 10399 433
rect 10399 381 10451 433
rect 10451 381 10453 433
rect 10397 379 10453 381
rect 10705 433 10761 435
rect 10705 381 10707 433
rect 10707 381 10759 433
rect 10759 381 10761 433
rect 10705 379 10761 381
rect 2539 375 2595 377
rect 4599 262 4655 264
rect 4599 210 4601 262
rect 4601 210 4653 262
rect 4653 210 4655 262
rect 4599 208 4655 210
rect 3588 103 3644 105
rect 3588 51 3590 103
rect 3590 51 3642 103
rect 3642 51 3644 103
rect 3588 49 3644 51
rect 3996 103 4052 105
rect 3996 51 3998 103
rect 3998 51 4050 103
rect 4050 51 4052 103
rect 3996 49 4052 51
rect 4404 103 4460 105
rect 4404 51 4406 103
rect 4406 51 4458 103
rect 4458 51 4460 103
rect 4404 49 4460 51
<< metal3 >>
rect -1496 17424 21670 17430
rect -1496 17360 -1490 17424
rect -1426 17360 -1354 17424
rect -1290 17360 -1218 17424
rect -1154 17360 21328 17424
rect 21392 17360 21464 17424
rect 21528 17360 21600 17424
rect 21664 17360 21670 17424
rect -1496 17288 21670 17360
rect -1496 17224 -1490 17288
rect -1426 17224 -1354 17288
rect -1290 17224 -1218 17288
rect -1154 17224 21328 17288
rect 21392 17224 21464 17288
rect 21528 17224 21600 17288
rect 21664 17224 21670 17288
rect -1496 17152 21670 17224
rect -1496 17088 -1490 17152
rect -1426 17088 -1354 17152
rect -1290 17088 -1218 17152
rect -1154 17088 3943 17152
rect 4007 17088 5989 17152
rect 6053 17088 16819 17152
rect 16883 17088 21328 17152
rect 21392 17088 21464 17152
rect 21528 17088 21600 17152
rect 21664 17088 21670 17152
rect -1496 17082 21670 17088
rect -800 16728 20974 16734
rect -800 16664 -794 16728
rect -730 16664 -658 16728
rect -594 16664 -522 16728
rect -458 16664 20632 16728
rect 20696 16664 20768 16728
rect 20832 16664 20904 16728
rect 20968 16664 20974 16728
rect -800 16592 20974 16664
rect -800 16528 -794 16592
rect -730 16528 -658 16592
rect -594 16528 -522 16592
rect -458 16528 20632 16592
rect 20696 16528 20768 16592
rect 20832 16528 20904 16592
rect 20968 16528 20974 16592
rect -800 16456 20974 16528
rect -800 16392 -794 16456
rect -730 16392 -658 16456
rect -594 16392 -522 16456
rect -458 16392 3321 16456
rect 3385 16392 4741 16456
rect 4805 16392 7940 16456
rect 8004 16392 12170 16456
rect 12234 16392 16401 16456
rect 16465 16392 19845 16456
rect 19909 16392 20632 16456
rect 20696 16392 20768 16456
rect 20832 16392 20904 16456
rect 20968 16392 20974 16456
rect -800 16386 20974 16392
rect 6948 15912 7046 15923
rect 19828 15912 19926 15923
rect 4735 15906 8010 15912
rect 4735 15902 7940 15906
rect 2026 15774 3391 15850
rect 2026 15704 2102 15774
rect 3315 15712 3391 15774
rect 4735 15846 6969 15902
rect 7025 15846 7940 15902
rect 4735 15842 7940 15846
rect 8004 15842 8010 15906
rect 4735 15836 8010 15842
rect 19828 15906 20702 15912
rect 19828 15842 19845 15906
rect 19909 15842 20632 15906
rect 20696 15842 20702 15906
rect 19828 15836 20702 15842
rect 4735 15712 4811 15836
rect 6948 15825 7046 15836
rect 19828 15825 19926 15836
rect 2026 15701 3242 15704
rect 3304 15701 3402 15712
rect 3926 15701 4024 15712
rect 2026 15698 3402 15701
rect -40 15634 -34 15698
rect 30 15634 36 15698
rect 2026 15634 2032 15698
rect 2096 15695 3402 15698
rect 2096 15634 3321 15695
rect 2026 15631 3321 15634
rect 3385 15631 3402 15695
rect 2026 15628 3402 15631
rect 3166 15625 3402 15628
rect 3304 15614 3402 15625
rect 3464 15695 4024 15701
rect 3464 15631 3943 15695
rect 4007 15631 4024 15695
rect 3464 15625 4024 15631
rect 3464 15552 3540 15625
rect 3926 15614 4024 15625
rect 4724 15695 4822 15712
rect 5972 15701 6070 15712
rect 4724 15631 4741 15695
rect 4805 15631 4822 15695
rect 4724 15614 4822 15631
rect 4884 15695 6070 15701
rect 4884 15631 5989 15695
rect 6053 15631 6070 15695
rect 4884 15625 6070 15631
rect -1224 15546 3540 15552
rect -1224 15482 -1218 15546
rect -1154 15482 3540 15546
rect -1224 15476 3540 15482
rect 3937 15552 4013 15614
rect 4884 15552 4960 15625
rect 5972 15614 6070 15625
rect 3937 15476 4960 15552
rect 13497 13999 13595 14010
rect 12164 13993 16471 13999
rect -528 13962 45 13968
rect -528 13898 -522 13962
rect -458 13898 -34 13962
rect 30 13898 45 13962
rect 2026 13898 2032 13962
rect 2096 13960 2102 13962
rect 2096 13900 2111 13960
rect 12164 13929 12170 13993
rect 12234 13929 13514 13993
rect 13578 13929 16401 13993
rect 16465 13929 16471 13993
rect 12164 13923 16471 13929
rect 13497 13912 13595 13923
rect 2096 13898 2102 13900
rect -528 13892 45 13898
rect 13497 12257 13595 12274
rect -528 12226 45 12232
rect -528 12162 -522 12226
rect -458 12162 -34 12226
rect 30 12162 45 12226
rect 2026 12162 2032 12226
rect 2096 12224 2102 12226
rect 2096 12164 2111 12224
rect 13497 12193 13514 12257
rect 13578 12193 13595 12257
rect 13497 12176 13595 12193
rect 2096 12162 2102 12164
rect -528 12156 45 12162
rect 13497 10527 13595 10538
rect 13497 10521 13733 10527
rect -528 10490 45 10496
rect -528 10426 -522 10490
rect -458 10426 -34 10490
rect 30 10426 45 10490
rect 2026 10426 2032 10490
rect 2096 10488 2102 10490
rect 2096 10428 2111 10488
rect 13497 10457 13514 10521
rect 13578 10457 13663 10521
rect 13727 10457 13733 10521
rect 13497 10451 13733 10457
rect 13497 10440 13595 10451
rect 2096 10426 2102 10428
rect -528 10420 45 10426
rect 3051 8850 4013 8926
rect -528 8754 45 8760
rect 2035 8754 2978 8760
rect -528 8690 -522 8754
rect -458 8690 45 8754
rect 1822 8690 1828 8754
rect 1892 8690 1898 8754
rect 2026 8690 2032 8754
rect 2096 8690 2978 8754
rect 3051 8736 3127 8850
rect 3937 8788 4013 8850
rect 13497 8791 13595 8802
rect 3304 8777 3402 8788
rect 3926 8777 4024 8788
rect 3304 8771 3864 8777
rect 3304 8767 3794 8771
rect -528 8684 45 8690
rect 2035 8684 2978 8690
rect 2902 8576 2978 8684
rect 3040 8719 3138 8736
rect 3040 8655 3057 8719
rect 3121 8655 3138 8719
rect 3304 8711 3325 8767
rect 3381 8711 3794 8767
rect 3304 8707 3794 8711
rect 3858 8707 3864 8771
rect 3304 8701 3864 8707
rect 3926 8767 4662 8777
rect 3926 8711 3947 8767
rect 4003 8711 4662 8767
rect 3926 8701 4662 8711
rect 3304 8690 3402 8701
rect 3926 8690 4024 8701
rect 3040 8638 3138 8655
rect 3315 8576 3391 8690
rect 2902 8500 3391 8576
rect 4586 8628 4662 8701
rect 4724 8771 4822 8788
rect 4724 8707 4741 8771
rect 4805 8707 4822 8771
rect 4724 8690 4822 8707
rect 5972 8777 6070 8788
rect 13497 8785 13733 8791
rect 5972 8771 6933 8777
rect 5972 8767 6863 8771
rect 5972 8711 5993 8767
rect 6049 8711 6863 8767
rect 5972 8707 6863 8711
rect 6927 8707 6933 8771
rect 5972 8701 6933 8707
rect 13497 8721 13514 8785
rect 13578 8721 13663 8785
rect 13727 8721 13733 8785
rect 13497 8715 13733 8721
rect 13497 8704 13595 8715
rect 5972 8690 6070 8701
rect 5983 8628 6059 8690
rect 4586 8552 6059 8628
rect 3788 8484 4811 8490
rect 3788 8420 3794 8484
rect 3858 8420 4741 8484
rect 4805 8420 4811 8484
rect 3788 8414 4811 8420
rect 92 8354 190 8365
rect -1224 8348 3127 8354
rect -1224 8284 -1218 8348
rect -1154 8284 109 8348
rect 173 8284 3057 8348
rect 3121 8284 3127 8348
rect -1224 8278 3127 8284
rect 92 8267 190 8278
rect 2132 7929 2230 7940
rect 1822 7923 2368 7929
rect 1822 7859 1828 7923
rect 1892 7859 2000 7923
rect 2064 7919 2298 7923
rect 2064 7863 2153 7919
rect 2209 7863 2298 7919
rect 2064 7859 2298 7863
rect 2362 7859 2368 7923
rect 1822 7853 2368 7859
rect 6846 7912 6944 7929
rect 2132 7842 2230 7853
rect 6846 7848 6863 7912
rect 6927 7848 6944 7912
rect 6846 7831 6944 7848
rect 92 7396 190 7413
rect 92 7332 109 7396
rect 173 7332 190 7396
rect 92 7315 190 7332
rect 6842 7262 6940 7273
rect 19898 7262 19996 7273
rect 6383 7256 6940 7262
rect 6383 7192 6389 7256
rect 6453 7192 6859 7256
rect 6923 7192 6940 7256
rect 6383 7186 6940 7192
rect 16813 7256 21398 7262
rect 16813 7192 16819 7256
rect 16883 7192 19915 7256
rect 19979 7192 21328 7256
rect 21392 7192 21398 7256
rect 16813 7186 21398 7192
rect 6842 7175 6940 7186
rect 19898 7175 19996 7186
rect 2132 6977 2230 6988
rect 2132 6971 2368 6977
rect 2132 6907 2149 6971
rect 2213 6907 2298 6971
rect 2362 6907 2368 6971
rect 2132 6901 2368 6907
rect 2132 6890 2230 6901
rect 92 6365 190 6376
rect -1224 6359 190 6365
rect -1224 6295 -1218 6359
rect -1154 6295 109 6359
rect 173 6295 190 6359
rect 6842 6346 6940 6357
rect -1224 6289 190 6295
rect 92 6278 190 6289
rect 5761 6340 6940 6346
rect 5761 6276 5767 6340
rect 5831 6336 6940 6340
rect 5831 6280 6863 6336
rect 6919 6280 6940 6336
rect 5831 6276 6940 6280
rect 5761 6270 6940 6276
rect 6842 6259 6940 6270
rect 19898 6346 19996 6357
rect 20898 6347 20974 6353
rect 20898 6346 20904 6347
rect 19898 6340 20904 6346
rect 19898 6336 20632 6340
rect 19898 6280 19919 6336
rect 19975 6280 20632 6336
rect 19898 6276 20632 6280
rect 20696 6283 20904 6340
rect 20968 6283 20974 6347
rect 20696 6276 20974 6283
rect 19898 6270 20974 6276
rect 19898 6259 19996 6270
rect -1496 6003 2024 6009
rect -1496 5939 1954 6003
rect 2018 5939 2024 6003
rect -1496 5933 2024 5939
rect -1496 5865 949 5871
rect -1496 5801 879 5865
rect 943 5801 949 5865
rect -1496 5795 949 5801
rect 13429 5838 13527 5855
rect 13429 5774 13446 5838
rect 13510 5774 13527 5838
rect 13429 5757 13527 5774
rect 2132 5743 2230 5754
rect 1686 5737 3298 5743
rect -1496 5657 541 5733
rect 1686 5673 1692 5737
rect 1756 5673 2149 5737
rect 2213 5673 2298 5737
rect 2362 5673 3228 5737
rect 3292 5673 3298 5737
rect 1686 5667 3298 5673
rect 305 5584 403 5595
rect -1496 5574 403 5584
rect -1496 5518 326 5574
rect 382 5518 403 5574
rect -1496 5508 403 5518
rect 465 5584 541 5657
rect 2132 5656 2230 5667
rect 713 5584 811 5595
rect 1121 5584 1219 5595
rect 1529 5584 1627 5595
rect 465 5574 811 5584
rect 465 5518 734 5574
rect 790 5518 811 5574
rect 465 5508 811 5518
rect 873 5578 1219 5584
rect 873 5514 879 5578
rect 943 5574 1219 5578
rect 943 5518 1142 5574
rect 1198 5518 1219 5574
rect 943 5514 1219 5518
rect 873 5508 1219 5514
rect 1281 5578 1627 5584
rect 1281 5514 1287 5578
rect 1351 5574 1627 5578
rect 1351 5518 1550 5574
rect 1606 5518 1627 5574
rect 1351 5514 1627 5518
rect 1281 5508 1627 5514
rect 305 5497 403 5508
rect 713 5497 811 5508
rect 1121 5497 1219 5508
rect 1529 5497 1627 5508
rect 1937 5578 2035 5595
rect 1937 5514 1954 5578
rect 2018 5514 2035 5578
rect 1937 5497 2035 5514
rect 1675 5428 1773 5439
rect -528 5422 1773 5428
rect -528 5358 -522 5422
rect -458 5358 1692 5422
rect 1756 5358 1773 5422
rect -528 5352 1773 5358
rect 1675 5341 1773 5352
rect -1496 5284 1357 5290
rect -1496 5220 1287 5284
rect 1351 5220 1357 5284
rect -1496 5214 1357 5220
rect 2292 5024 5688 5027
rect 5750 5024 5848 5035
rect 2292 5021 5848 5024
rect 2292 4957 2298 5021
rect 2362 4957 3228 5021
rect 3292 5018 5848 5021
rect 3292 4957 5767 5018
rect 2292 4954 5767 4957
rect 5831 4954 5848 5018
rect 2292 4951 5848 4954
rect 5612 4948 5848 4951
rect 5750 4937 5848 4948
rect 6372 5018 6470 5035
rect 6372 4954 6389 5018
rect 6453 4954 6470 5018
rect 6372 4937 6470 4954
rect 5497 3381 5986 3457
rect 3222 3285 4557 3291
rect 3222 3221 4274 3285
rect 4338 3221 4487 3285
rect 4551 3221 4557 3285
rect 5497 3267 5573 3381
rect 5750 3302 5848 3319
rect 5486 3256 5584 3267
rect 3222 3215 4557 3221
rect 4481 3107 4557 3215
rect 4627 3250 5584 3256
rect 4627 3186 4633 3250
rect 4697 3246 5584 3250
rect 4697 3190 5507 3246
rect 5563 3190 5584 3246
rect 5750 3238 5767 3302
rect 5831 3238 5848 3302
rect 5750 3221 5848 3238
rect 5910 3308 5986 3381
rect 6372 3308 6470 3319
rect 5910 3302 8447 3308
rect 5910 3238 6389 3302
rect 6453 3238 8377 3302
rect 8441 3238 8447 3302
rect 5910 3232 8447 3238
rect 6372 3221 6470 3232
rect 4697 3186 5584 3190
rect 4627 3180 5584 3186
rect 5486 3169 5584 3180
rect 5761 3107 5837 3221
rect 4481 3031 5837 3107
rect 3354 2885 3452 2896
rect 1543 2879 4703 2885
rect 1543 2815 3371 2879
rect 3435 2815 4633 2879
rect 4697 2815 4703 2879
rect 1383 2799 1481 2810
rect 1543 2809 4703 2815
rect 1543 2799 1619 2809
rect -1224 2793 1619 2799
rect 3354 2798 3452 2809
rect -1224 2729 -1218 2793
rect -1154 2729 1619 2793
rect -1224 2723 1619 2729
rect 1383 2712 1481 2723
rect 4578 2460 4676 2471
rect 4268 2454 4814 2460
rect 4268 2390 4274 2454
rect 4338 2390 4446 2454
rect 4510 2450 4744 2454
rect 4510 2394 4599 2450
rect 4655 2394 4744 2450
rect 4510 2390 4744 2394
rect 4808 2390 4814 2454
rect 4268 2384 4814 2390
rect 4578 2373 4676 2384
rect 3354 1927 3452 1944
rect 3354 1863 3371 1927
rect 3435 1863 3452 1927
rect 8360 1880 8458 1891
rect 10804 1880 10902 1891
rect 3354 1846 3452 1863
rect 5761 1874 16471 1880
rect 5761 1810 5767 1874
rect 5831 1810 7940 1874
rect 8004 1870 12170 1874
rect 8004 1814 8381 1870
rect 8437 1814 10825 1870
rect 10881 1814 12170 1870
rect 8004 1810 12170 1814
rect 12234 1810 13446 1874
rect 13510 1810 16401 1874
rect 16465 1810 16471 1874
rect 5761 1804 16471 1810
rect 8360 1793 8458 1804
rect 10804 1793 10902 1804
rect 4578 1508 4676 1519
rect 4578 1502 4814 1508
rect 458 1448 556 1459
rect -1496 1438 556 1448
rect -1496 1382 479 1438
rect 535 1382 556 1438
rect 4578 1438 4595 1502
rect 4659 1438 4744 1502
rect 4808 1438 4814 1502
rect 4578 1432 4814 1438
rect 4578 1421 4676 1432
rect -1496 1372 556 1382
rect 458 1361 556 1372
rect 8360 964 8458 975
rect 10804 964 10902 975
rect 7794 958 16889 964
rect 3354 890 3452 907
rect 3354 826 3371 890
rect 3435 826 3452 890
rect 7794 894 7800 958
rect 7864 894 8377 958
rect 8441 954 12310 958
rect 8441 898 10825 954
rect 10881 898 12310 954
rect 8441 894 12310 898
rect 12374 894 16819 958
rect 16883 894 16889 958
rect 7794 888 16889 894
rect 8360 877 8458 888
rect 10804 877 10902 888
rect 3354 809 3452 826
rect 2518 435 2616 452
rect 2518 371 2535 435
rect 2599 371 2616 435
rect 2518 354 2616 371
rect 8528 439 8626 456
rect 8528 375 8545 439
rect 8609 375 8626 439
rect 8528 358 8626 375
rect 8836 439 8934 456
rect 8836 375 8853 439
rect 8917 375 8934 439
rect 8836 358 8934 375
rect 9144 439 9242 456
rect 9144 375 9161 439
rect 9225 375 9242 439
rect 9144 358 9242 375
rect 9452 439 9550 456
rect 9452 375 9469 439
rect 9533 375 9550 439
rect 9452 358 9550 375
rect 9760 439 9858 456
rect 9760 375 9777 439
rect 9841 375 9858 439
rect 9760 358 9858 375
rect 10068 439 10166 456
rect 10068 375 10085 439
rect 10149 375 10166 439
rect 10068 358 10166 375
rect 10376 439 10474 456
rect 10376 375 10393 439
rect 10457 375 10474 439
rect 10376 358 10474 375
rect 10684 439 10782 456
rect 10684 375 10701 439
rect 10765 375 10782 439
rect 10684 358 10782 375
rect 4578 274 4676 285
rect 3703 268 4676 274
rect 3703 204 3709 268
rect 3773 204 4595 268
rect 4659 204 4676 268
rect 3703 198 4676 204
rect 4578 187 4676 198
rect 1383 165 1481 182
rect 1383 101 1400 165
rect 1464 101 1481 165
rect 1383 84 1481 101
rect 3567 105 3665 126
rect 3567 49 3588 105
rect 3644 49 3665 105
rect 3567 28 3665 49
rect 3975 109 4073 126
rect 3975 45 3992 109
rect 4056 45 4073 109
rect 3975 28 4073 45
rect 4383 109 4481 126
rect 4383 45 4400 109
rect 4464 45 4481 109
rect 4383 28 4481 45
rect 3578 -34 3654 28
rect 3565 -40 3654 -34
rect 3565 -104 3571 -40
rect 3635 -104 3654 -40
rect 3565 -110 3654 -104
rect -800 -458 20974 -452
rect -800 -522 -794 -458
rect -730 -522 -658 -458
rect -594 -522 -522 -458
rect -458 -522 1400 -458
rect 1464 -522 3709 -458
rect 3773 -522 7940 -458
rect 8004 -522 12170 -458
rect 12234 -522 16401 -458
rect 16465 -522 20632 -458
rect 20696 -522 20768 -458
rect 20832 -522 20904 -458
rect 20968 -522 20974 -458
rect -800 -594 20974 -522
rect -800 -658 -794 -594
rect -730 -658 -658 -594
rect -594 -658 -522 -594
rect -458 -658 20632 -594
rect 20696 -658 20768 -594
rect 20832 -658 20904 -594
rect 20968 -658 20974 -594
rect -800 -730 20974 -658
rect -800 -794 -794 -730
rect -730 -794 -658 -730
rect -594 -794 -522 -730
rect -458 -794 20632 -730
rect 20696 -794 20768 -730
rect 20832 -794 20904 -730
rect 20968 -794 20974 -730
rect -800 -800 20974 -794
rect -1496 -1154 21670 -1148
rect -1496 -1218 -1490 -1154
rect -1426 -1218 -1354 -1154
rect -1290 -1218 -1218 -1154
rect -1154 -1218 3371 -1154
rect 3435 -1218 7800 -1154
rect 7864 -1218 12310 -1154
rect 12374 -1218 16819 -1154
rect 16883 -1218 19915 -1154
rect 19979 -1218 21328 -1154
rect 21392 -1218 21464 -1154
rect 21528 -1218 21600 -1154
rect 21664 -1218 21670 -1154
rect -1496 -1290 21670 -1218
rect -1496 -1354 -1490 -1290
rect -1426 -1354 -1354 -1290
rect -1290 -1354 -1218 -1290
rect -1154 -1354 21328 -1290
rect 21392 -1354 21464 -1290
rect 21528 -1354 21600 -1290
rect 21664 -1354 21670 -1290
rect -1496 -1426 21670 -1354
rect -1496 -1490 -1490 -1426
rect -1426 -1490 -1354 -1426
rect -1290 -1490 -1218 -1426
rect -1154 -1490 21328 -1426
rect 21392 -1490 21464 -1426
rect 21528 -1490 21600 -1426
rect 21664 -1490 21670 -1426
rect -1496 -1496 21670 -1490
<< via3 >>
rect -1490 17360 -1426 17424
rect -1354 17360 -1290 17424
rect -1218 17360 -1154 17424
rect 21328 17360 21392 17424
rect 21464 17360 21528 17424
rect 21600 17360 21664 17424
rect -1490 17224 -1426 17288
rect -1354 17224 -1290 17288
rect -1218 17224 -1154 17288
rect 21328 17224 21392 17288
rect 21464 17224 21528 17288
rect 21600 17224 21664 17288
rect -1490 17088 -1426 17152
rect -1354 17088 -1290 17152
rect -1218 17088 -1154 17152
rect 3943 17088 4007 17152
rect 5989 17088 6053 17152
rect 16819 17088 16883 17152
rect 21328 17088 21392 17152
rect 21464 17088 21528 17152
rect 21600 17088 21664 17152
rect -794 16664 -730 16728
rect -658 16664 -594 16728
rect -522 16664 -458 16728
rect 20632 16664 20696 16728
rect 20768 16664 20832 16728
rect 20904 16664 20968 16728
rect -794 16528 -730 16592
rect -658 16528 -594 16592
rect -522 16528 -458 16592
rect 20632 16528 20696 16592
rect 20768 16528 20832 16592
rect 20904 16528 20968 16592
rect -794 16392 -730 16456
rect -658 16392 -594 16456
rect -522 16392 -458 16456
rect 3321 16392 3385 16456
rect 4741 16392 4805 16456
rect 7940 16392 8004 16456
rect 12170 16392 12234 16456
rect 16401 16392 16465 16456
rect 19845 16392 19909 16456
rect 20632 16392 20696 16456
rect 20768 16392 20832 16456
rect 20904 16392 20968 16456
rect 7940 15842 8004 15906
rect 19845 15902 19909 15906
rect 19845 15846 19849 15902
rect 19849 15846 19905 15902
rect 19905 15846 19909 15902
rect 19845 15842 19909 15846
rect 20632 15842 20696 15906
rect -34 15634 30 15698
rect 2032 15634 2096 15698
rect 3321 15691 3385 15695
rect 3321 15635 3325 15691
rect 3325 15635 3381 15691
rect 3381 15635 3385 15691
rect 3321 15631 3385 15635
rect 3943 15691 4007 15695
rect 3943 15635 3947 15691
rect 3947 15635 4003 15691
rect 4003 15635 4007 15691
rect 3943 15631 4007 15635
rect 4741 15691 4805 15695
rect 4741 15635 4745 15691
rect 4745 15635 4801 15691
rect 4801 15635 4805 15691
rect 4741 15631 4805 15635
rect 5989 15691 6053 15695
rect 5989 15635 5993 15691
rect 5993 15635 6049 15691
rect 6049 15635 6053 15691
rect 5989 15631 6053 15635
rect -1218 15482 -1154 15546
rect -522 13898 -458 13962
rect -34 13898 30 13962
rect 2032 13898 2096 13962
rect 12170 13929 12234 13993
rect 13514 13989 13578 13993
rect 13514 13933 13518 13989
rect 13518 13933 13574 13989
rect 13574 13933 13578 13989
rect 13514 13929 13578 13933
rect 16401 13929 16465 13993
rect -522 12162 -458 12226
rect -34 12162 30 12226
rect 2032 12162 2096 12226
rect 13514 12253 13578 12257
rect 13514 12197 13518 12253
rect 13518 12197 13574 12253
rect 13574 12197 13578 12253
rect 13514 12193 13578 12197
rect -522 10426 -458 10490
rect -34 10426 30 10490
rect 2032 10426 2096 10490
rect 13514 10517 13578 10521
rect 13514 10461 13518 10517
rect 13518 10461 13574 10517
rect 13574 10461 13578 10517
rect 13514 10457 13578 10461
rect 13663 10457 13727 10521
rect -522 8690 -458 8754
rect 1828 8690 1892 8754
rect 2032 8690 2096 8754
rect 3057 8715 3121 8719
rect 3057 8659 3061 8715
rect 3061 8659 3117 8715
rect 3117 8659 3121 8715
rect 3057 8655 3121 8659
rect 3794 8707 3858 8771
rect 4741 8767 4805 8771
rect 4741 8711 4745 8767
rect 4745 8711 4801 8767
rect 4801 8711 4805 8767
rect 4741 8707 4805 8711
rect 6863 8707 6927 8771
rect 13514 8781 13578 8785
rect 13514 8725 13518 8781
rect 13518 8725 13574 8781
rect 13574 8725 13578 8781
rect 13514 8721 13578 8725
rect 13663 8721 13727 8785
rect 3794 8420 3858 8484
rect 4741 8420 4805 8484
rect -1218 8284 -1154 8348
rect 109 8344 173 8348
rect 109 8288 113 8344
rect 113 8288 169 8344
rect 169 8288 173 8344
rect 109 8284 173 8288
rect 3057 8284 3121 8348
rect 1828 7859 1892 7923
rect 2000 7859 2064 7923
rect 2298 7859 2362 7923
rect 6863 7908 6927 7912
rect 6863 7852 6867 7908
rect 6867 7852 6923 7908
rect 6923 7852 6927 7908
rect 6863 7848 6927 7852
rect 109 7392 173 7396
rect 109 7336 113 7392
rect 113 7336 169 7392
rect 169 7336 173 7392
rect 109 7332 173 7336
rect 6389 7192 6453 7256
rect 6859 7252 6923 7256
rect 6859 7196 6863 7252
rect 6863 7196 6919 7252
rect 6919 7196 6923 7252
rect 6859 7192 6923 7196
rect 16819 7192 16883 7256
rect 19915 7252 19979 7256
rect 19915 7196 19919 7252
rect 19919 7196 19975 7252
rect 19975 7196 19979 7252
rect 19915 7192 19979 7196
rect 21328 7192 21392 7256
rect 2149 6967 2213 6971
rect 2149 6911 2153 6967
rect 2153 6911 2209 6967
rect 2209 6911 2213 6967
rect 2149 6907 2213 6911
rect 2298 6907 2362 6971
rect -1218 6295 -1154 6359
rect 109 6355 173 6359
rect 109 6299 113 6355
rect 113 6299 169 6355
rect 169 6299 173 6355
rect 109 6295 173 6299
rect 5767 6276 5831 6340
rect 20632 6276 20696 6340
rect 20904 6283 20968 6347
rect 1954 5939 2018 6003
rect 879 5801 943 5865
rect 13446 5834 13510 5838
rect 13446 5778 13450 5834
rect 13450 5778 13506 5834
rect 13506 5778 13510 5834
rect 13446 5774 13510 5778
rect 1692 5673 1756 5737
rect 2149 5733 2213 5737
rect 2149 5677 2153 5733
rect 2153 5677 2209 5733
rect 2209 5677 2213 5733
rect 2149 5673 2213 5677
rect 2298 5673 2362 5737
rect 3228 5673 3292 5737
rect 879 5514 943 5578
rect 1287 5514 1351 5578
rect 1954 5574 2018 5578
rect 1954 5518 1958 5574
rect 1958 5518 2014 5574
rect 2014 5518 2018 5574
rect 1954 5514 2018 5518
rect -522 5358 -458 5422
rect 1692 5358 1756 5422
rect 1287 5220 1351 5284
rect 2298 4957 2362 5021
rect 3228 4957 3292 5021
rect 5767 5014 5831 5018
rect 5767 4958 5771 5014
rect 5771 4958 5827 5014
rect 5827 4958 5831 5014
rect 5767 4954 5831 4958
rect 6389 5014 6453 5018
rect 6389 4958 6393 5014
rect 6393 4958 6449 5014
rect 6449 4958 6453 5014
rect 6389 4954 6453 4958
rect 4274 3221 4338 3285
rect 4487 3221 4551 3285
rect 4633 3186 4697 3250
rect 5767 3298 5831 3302
rect 5767 3242 5771 3298
rect 5771 3242 5827 3298
rect 5827 3242 5831 3298
rect 5767 3238 5831 3242
rect 6389 3298 6453 3302
rect 6389 3242 6393 3298
rect 6393 3242 6449 3298
rect 6449 3242 6453 3298
rect 6389 3238 6453 3242
rect 8377 3238 8441 3302
rect 3371 2875 3435 2879
rect 3371 2819 3375 2875
rect 3375 2819 3431 2875
rect 3431 2819 3435 2875
rect 3371 2815 3435 2819
rect 4633 2815 4697 2879
rect -1218 2729 -1154 2793
rect 4274 2390 4338 2454
rect 4446 2390 4510 2454
rect 4744 2390 4808 2454
rect 3371 1923 3435 1927
rect 3371 1867 3375 1923
rect 3375 1867 3431 1923
rect 3431 1867 3435 1923
rect 3371 1863 3435 1867
rect 5767 1810 5831 1874
rect 7940 1810 8004 1874
rect 12170 1810 12234 1874
rect 13446 1810 13510 1874
rect 16401 1810 16465 1874
rect 4595 1498 4659 1502
rect 4595 1442 4599 1498
rect 4599 1442 4655 1498
rect 4655 1442 4659 1498
rect 4595 1438 4659 1442
rect 4744 1438 4808 1502
rect 3371 886 3435 890
rect 3371 830 3375 886
rect 3375 830 3431 886
rect 3431 830 3435 886
rect 3371 826 3435 830
rect 7800 894 7864 958
rect 8377 954 8441 958
rect 8377 898 8381 954
rect 8381 898 8437 954
rect 8437 898 8441 954
rect 8377 894 8441 898
rect 12310 894 12374 958
rect 16819 894 16883 958
rect 2535 431 2599 435
rect 2535 375 2539 431
rect 2539 375 2595 431
rect 2595 375 2599 431
rect 2535 371 2599 375
rect 8545 435 8609 439
rect 8545 379 8549 435
rect 8549 379 8605 435
rect 8605 379 8609 435
rect 8545 375 8609 379
rect 8853 435 8917 439
rect 8853 379 8857 435
rect 8857 379 8913 435
rect 8913 379 8917 435
rect 8853 375 8917 379
rect 9161 435 9225 439
rect 9161 379 9165 435
rect 9165 379 9221 435
rect 9221 379 9225 435
rect 9161 375 9225 379
rect 9469 435 9533 439
rect 9469 379 9473 435
rect 9473 379 9529 435
rect 9529 379 9533 435
rect 9469 375 9533 379
rect 9777 435 9841 439
rect 9777 379 9781 435
rect 9781 379 9837 435
rect 9837 379 9841 435
rect 9777 375 9841 379
rect 10085 435 10149 439
rect 10085 379 10089 435
rect 10089 379 10145 435
rect 10145 379 10149 435
rect 10085 375 10149 379
rect 10393 435 10457 439
rect 10393 379 10397 435
rect 10397 379 10453 435
rect 10453 379 10457 435
rect 10393 375 10457 379
rect 10701 435 10765 439
rect 10701 379 10705 435
rect 10705 379 10761 435
rect 10761 379 10765 435
rect 10701 375 10765 379
rect 3709 204 3773 268
rect 4595 264 4659 268
rect 4595 208 4599 264
rect 4599 208 4655 264
rect 4655 208 4659 264
rect 4595 204 4659 208
rect 1400 101 1464 165
rect 3992 105 4056 109
rect 3992 49 3996 105
rect 3996 49 4052 105
rect 4052 49 4056 105
rect 3992 45 4056 49
rect 4400 105 4464 109
rect 4400 49 4404 105
rect 4404 49 4460 105
rect 4460 49 4464 105
rect 4400 45 4464 49
rect 3571 -104 3635 -40
rect -794 -522 -730 -458
rect -658 -522 -594 -458
rect -522 -522 -458 -458
rect 1400 -522 1464 -458
rect 3709 -522 3773 -458
rect 7940 -522 8004 -458
rect 12170 -522 12234 -458
rect 16401 -522 16465 -458
rect 20632 -522 20696 -458
rect 20768 -522 20832 -458
rect 20904 -522 20968 -458
rect -794 -658 -730 -594
rect -658 -658 -594 -594
rect -522 -658 -458 -594
rect 20632 -658 20696 -594
rect 20768 -658 20832 -594
rect 20904 -658 20968 -594
rect -794 -794 -730 -730
rect -658 -794 -594 -730
rect -522 -794 -458 -730
rect 20632 -794 20696 -730
rect 20768 -794 20832 -730
rect 20904 -794 20968 -730
rect -1490 -1218 -1426 -1154
rect -1354 -1218 -1290 -1154
rect -1218 -1218 -1154 -1154
rect 3371 -1218 3435 -1154
rect 7800 -1218 7864 -1154
rect 12310 -1218 12374 -1154
rect 16819 -1218 16883 -1154
rect 19915 -1218 19979 -1154
rect 21328 -1218 21392 -1154
rect 21464 -1218 21528 -1154
rect 21600 -1218 21664 -1154
rect -1490 -1354 -1426 -1290
rect -1354 -1354 -1290 -1290
rect -1218 -1354 -1154 -1290
rect 21328 -1354 21392 -1290
rect 21464 -1354 21528 -1290
rect 21600 -1354 21664 -1290
rect -1490 -1490 -1426 -1426
rect -1354 -1490 -1290 -1426
rect -1218 -1490 -1154 -1426
rect 21328 -1490 21392 -1426
rect 21464 -1490 21528 -1426
rect 21600 -1490 21664 -1426
<< metal4 >>
rect -1496 17424 -1148 17430
rect -1496 17360 -1490 17424
rect -1426 17360 -1354 17424
rect -1290 17360 -1218 17424
rect -1154 17360 -1148 17424
rect -1496 17288 -1148 17360
rect -1496 17224 -1490 17288
rect -1426 17224 -1354 17288
rect -1290 17224 -1218 17288
rect -1154 17224 -1148 17288
rect -1496 17152 -1148 17224
rect 21322 17424 21670 17430
rect 21322 17360 21328 17424
rect 21392 17360 21464 17424
rect 21528 17360 21600 17424
rect 21664 17360 21670 17424
rect 21322 17288 21670 17360
rect 21322 17224 21328 17288
rect 21392 17224 21464 17288
rect 21528 17224 21600 17288
rect 21664 17224 21670 17288
rect -1496 17088 -1490 17152
rect -1426 17088 -1354 17152
rect -1290 17088 -1218 17152
rect -1154 17088 -1148 17152
rect -1496 15546 -1148 17088
rect 3937 17152 4013 17158
rect 3937 17088 3943 17152
rect 4007 17088 4013 17152
rect -1496 15482 -1218 15546
rect -1154 15482 -1148 15546
rect -1496 8348 -1148 15482
rect -1496 8284 -1218 8348
rect -1154 8284 -1148 8348
rect -1496 6359 -1148 8284
rect -1496 6295 -1218 6359
rect -1154 6295 -1148 6359
rect -1496 2793 -1148 6295
rect -1496 2729 -1218 2793
rect -1154 2729 -1148 2793
rect -1496 -1154 -1148 2729
rect -800 16728 -452 16734
rect -800 16664 -794 16728
rect -730 16664 -658 16728
rect -594 16664 -522 16728
rect -458 16664 -452 16728
rect -800 16592 -452 16664
rect -800 16528 -794 16592
rect -730 16528 -658 16592
rect -594 16528 -522 16592
rect -458 16528 -452 16592
rect -800 16456 -452 16528
rect -800 16392 -794 16456
rect -730 16392 -658 16456
rect -594 16392 -522 16456
rect -458 16392 -452 16456
rect -800 13962 -452 16392
rect 3315 16456 3391 16462
rect 3315 16392 3321 16456
rect 3385 16392 3391 16456
rect -800 13898 -522 13962
rect -458 13898 -452 13962
rect -800 12226 -452 13898
rect -40 15698 36 15704
rect -40 15634 -34 15698
rect 30 15634 36 15698
rect -40 13962 36 15634
rect -40 13898 -34 13962
rect 30 13898 36 13962
rect -40 13892 36 13898
rect 2026 15698 2102 15704
rect 2026 15634 2032 15698
rect 2096 15634 2102 15698
rect 2026 13962 2102 15634
rect 3315 15695 3391 16392
rect 3315 15631 3321 15695
rect 3385 15631 3391 15695
rect 3315 15625 3391 15631
rect 3937 15695 4013 17088
rect 5983 17152 6059 17158
rect 5983 17088 5989 17152
rect 6053 17088 6059 17152
rect 3937 15631 3943 15695
rect 4007 15631 4013 15695
rect 3937 15625 4013 15631
rect 4735 16456 4811 16462
rect 4735 16392 4741 16456
rect 4805 16392 4811 16456
rect 4735 15695 4811 16392
rect 4735 15631 4741 15695
rect 4805 15631 4811 15695
rect 4735 15625 4811 15631
rect 5983 15695 6059 17088
rect 16813 17152 16889 17158
rect 16813 17088 16819 17152
rect 16883 17088 16889 17152
rect 7934 16456 8010 16462
rect 7934 16392 7940 16456
rect 8004 16392 8010 16456
rect 7934 15906 8010 16392
rect 7934 15842 7940 15906
rect 8004 15842 8010 15906
rect 7934 15836 8010 15842
rect 12164 16456 12240 16462
rect 12164 16392 12170 16456
rect 12234 16392 12240 16456
rect 5983 15631 5989 15695
rect 6053 15631 6059 15695
rect 5983 15625 6059 15631
rect 2026 13898 2032 13962
rect 2096 13898 2102 13962
rect 12164 13993 12240 16392
rect 16395 16456 16471 16462
rect 16395 16392 16401 16456
rect 16465 16392 16471 16456
rect 12164 13929 12170 13993
rect 12234 13929 12240 13993
rect 12164 13923 12240 13929
rect 13508 13993 13584 13999
rect 13508 13929 13514 13993
rect 13578 13929 13584 13993
rect -800 12162 -522 12226
rect -458 12162 -452 12226
rect -800 10490 -452 12162
rect -800 10426 -522 10490
rect -458 10426 -452 10490
rect -800 8754 -452 10426
rect -40 12226 36 12232
rect -40 12162 -34 12226
rect 30 12162 36 12226
rect -40 10490 36 12162
rect -40 10426 -34 10490
rect 30 10426 36 10490
rect -40 10420 36 10426
rect 2026 12226 2102 13898
rect 2026 12162 2032 12226
rect 2096 12162 2102 12226
rect 2026 10490 2102 12162
rect 2026 10426 2032 10490
rect 2096 10426 2102 10490
rect 13508 12257 13584 13929
rect 16395 13993 16471 16392
rect 16395 13929 16401 13993
rect 16465 13929 16471 13993
rect 16395 13923 16471 13929
rect 13508 12193 13514 12257
rect 13578 12193 13584 12257
rect 13508 10521 13584 12193
rect 13508 10457 13514 10521
rect 13578 10457 13584 10521
rect 13508 10451 13584 10457
rect 13657 10521 13733 10527
rect 13657 10457 13663 10521
rect 13727 10457 13733 10521
rect -800 8690 -522 8754
rect -458 8690 -452 8754
rect -800 5422 -452 8690
rect 1822 8754 1898 8760
rect 1822 8690 1828 8754
rect 1892 8690 1898 8754
rect 103 8348 179 8354
rect 103 8284 109 8348
rect 173 8284 179 8348
rect 103 7396 179 8284
rect 1822 7923 1898 8690
rect 2026 8754 2102 10426
rect 13440 8785 13584 8791
rect 2026 8690 2032 8754
rect 2096 8690 2102 8754
rect 3788 8771 3864 8777
rect 2026 7929 2102 8690
rect 3051 8719 3127 8725
rect 3051 8655 3057 8719
rect 3121 8655 3127 8719
rect 3051 8348 3127 8655
rect 3788 8707 3794 8771
rect 3858 8707 3864 8771
rect 3788 8484 3864 8707
rect 3788 8420 3794 8484
rect 3858 8420 3864 8484
rect 3788 8414 3864 8420
rect 4735 8771 4811 8777
rect 4735 8707 4741 8771
rect 4805 8707 4811 8771
rect 4735 8484 4811 8707
rect 4735 8420 4741 8484
rect 4805 8420 4811 8484
rect 4735 8414 4811 8420
rect 6857 8771 6933 8777
rect 6857 8707 6863 8771
rect 6927 8707 6933 8771
rect 3051 8284 3057 8348
rect 3121 8284 3127 8348
rect 3051 8278 3127 8284
rect 1822 7859 1828 7923
rect 1892 7859 1898 7923
rect 1822 7853 1898 7859
rect 1994 7923 2102 7929
rect 1994 7859 2000 7923
rect 2064 7859 2102 7923
rect 1994 7853 2102 7859
rect 2292 7923 2368 7929
rect 2292 7859 2298 7923
rect 2362 7859 2368 7923
rect 103 7332 109 7396
rect 173 7332 179 7396
rect 103 6359 179 7332
rect 103 6295 109 6359
rect 173 6295 179 6359
rect 103 6289 179 6295
rect 2143 6971 2219 6977
rect 2143 6907 2149 6971
rect 2213 6907 2219 6971
rect 1948 6003 2024 6009
rect 1948 5939 1954 6003
rect 2018 5939 2024 6003
rect 873 5865 949 5871
rect 873 5801 879 5865
rect 943 5801 949 5865
rect 873 5578 949 5801
rect 1686 5737 1762 5743
rect 1686 5673 1692 5737
rect 1756 5673 1762 5737
rect 873 5514 879 5578
rect 943 5514 949 5578
rect 873 5508 949 5514
rect 1281 5578 1357 5584
rect 1281 5514 1287 5578
rect 1351 5514 1357 5578
rect -800 5358 -522 5422
rect -458 5358 -452 5422
rect -800 -458 -452 5358
rect 1281 5284 1357 5514
rect 1686 5422 1762 5673
rect 1948 5578 2024 5939
rect 2143 5737 2219 6907
rect 2292 6971 2368 7859
rect 6857 7912 6933 8707
rect 6857 7848 6863 7912
rect 6927 7848 6933 7912
rect 6857 7262 6933 7848
rect 2292 6907 2298 6971
rect 2362 6907 2368 6971
rect 2292 6901 2368 6907
rect 6383 7256 6459 7262
rect 6383 7192 6389 7256
rect 6453 7192 6459 7256
rect 5761 6340 5837 6346
rect 5761 6276 5767 6340
rect 5831 6276 5837 6340
rect 2143 5673 2149 5737
rect 2213 5673 2219 5737
rect 2143 5667 2219 5673
rect 2292 5737 2368 5743
rect 2292 5673 2298 5737
rect 2362 5673 2368 5737
rect 1948 5514 1954 5578
rect 2018 5514 2024 5578
rect 1948 5508 2024 5514
rect 1686 5358 1692 5422
rect 1756 5358 1762 5422
rect 1686 5352 1762 5358
rect 1281 5220 1287 5284
rect 1351 5220 1357 5284
rect 1281 5214 1357 5220
rect 2292 5021 2368 5673
rect 2292 4957 2298 5021
rect 2362 4957 2368 5021
rect 2292 4951 2368 4957
rect 3222 5737 3298 5743
rect 3222 5673 3228 5737
rect 3292 5673 3298 5737
rect 3222 5021 3298 5673
rect 3222 4957 3228 5021
rect 3292 4957 3298 5021
rect 3222 4951 3298 4957
rect 5761 5018 5837 6276
rect 5761 4954 5767 5018
rect 5831 4954 5837 5018
rect 5761 3302 5837 4954
rect 4268 3285 4344 3291
rect 4268 3221 4274 3285
rect 4338 3221 4344 3285
rect 3365 2879 3441 2885
rect 3365 2815 3371 2879
rect 3435 2815 3441 2879
rect 3365 1927 3441 2815
rect 4268 2454 4344 3221
rect 4481 3285 4557 3291
rect 4481 3221 4487 3285
rect 4551 3221 4557 3285
rect 4481 2460 4557 3221
rect 4627 3250 4703 3256
rect 4627 3186 4633 3250
rect 4697 3186 4703 3250
rect 4627 2879 4703 3186
rect 4627 2815 4633 2879
rect 4697 2815 4703 2879
rect 4627 2809 4703 2815
rect 5761 3238 5767 3302
rect 5831 3238 5837 3302
rect 4268 2390 4274 2454
rect 4338 2390 4344 2454
rect 4268 2384 4344 2390
rect 4440 2454 4557 2460
rect 4440 2390 4446 2454
rect 4510 2390 4557 2454
rect 4440 2384 4557 2390
rect 4738 2454 4814 2460
rect 4738 2390 4744 2454
rect 4808 2390 4814 2454
rect 3365 1863 3371 1927
rect 3435 1863 3441 1927
rect 3365 890 3441 1863
rect 3365 826 3371 890
rect 3435 826 3441 890
rect 2529 435 2605 441
rect 2529 371 2535 435
rect 2599 371 2605 435
rect -800 -522 -794 -458
rect -730 -522 -658 -458
rect -594 -522 -522 -458
rect -458 -522 -452 -458
rect -800 -594 -452 -522
rect 1394 165 1470 171
rect 1394 101 1400 165
rect 1464 101 1470 165
rect 1394 -458 1470 101
rect 1394 -522 1400 -458
rect 1464 -522 1470 -458
rect 1394 -528 1470 -522
rect -800 -658 -794 -594
rect -730 -658 -658 -594
rect -594 -658 -522 -594
rect -458 -658 -452 -594
rect -800 -730 -452 -658
rect -800 -794 -794 -730
rect -730 -794 -658 -730
rect -594 -794 -522 -730
rect -458 -794 -452 -730
rect -800 -800 -452 -794
rect -1496 -1218 -1490 -1154
rect -1426 -1218 -1354 -1154
rect -1290 -1218 -1218 -1154
rect -1154 -1218 -1148 -1154
rect -1496 -1290 -1148 -1218
rect -1496 -1354 -1490 -1290
rect -1426 -1354 -1354 -1290
rect -1290 -1354 -1218 -1290
rect -1154 -1354 -1148 -1290
rect -1496 -1426 -1148 -1354
rect -1496 -1490 -1490 -1426
rect -1426 -1490 -1354 -1426
rect -1290 -1490 -1218 -1426
rect -1154 -1490 -1148 -1426
rect -1496 -1496 -1148 -1490
rect 2529 -1496 2605 371
rect 3365 -1154 3441 826
rect 4589 1502 4665 1508
rect 4589 1438 4595 1502
rect 4659 1438 4665 1502
rect 3703 268 3779 274
rect 3703 204 3709 268
rect 3773 204 3779 268
rect 3365 -1218 3371 -1154
rect 3435 -1218 3441 -1154
rect 3365 -1224 3441 -1218
rect 3565 -40 3641 -34
rect 3565 -104 3571 -40
rect 3635 -104 3641 -40
rect 3565 -1496 3641 -104
rect 3703 -458 3779 204
rect 4589 268 4665 1438
rect 4738 1502 4814 2390
rect 5761 1874 5837 3238
rect 6383 5018 6459 7192
rect 6853 7256 6933 7262
rect 6853 7192 6859 7256
rect 6923 7192 6933 7256
rect 6853 7186 6933 7192
rect 13440 8721 13514 8785
rect 13578 8721 13584 8785
rect 13440 8715 13584 8721
rect 13657 8785 13733 10457
rect 13657 8721 13663 8785
rect 13727 8721 13733 8785
rect 13657 8715 13733 8721
rect 6383 4954 6389 5018
rect 6453 4954 6459 5018
rect 6383 3302 6459 4954
rect 13440 5838 13516 8715
rect 16813 7256 16889 17088
rect 21322 17152 21670 17224
rect 21322 17088 21328 17152
rect 21392 17088 21464 17152
rect 21528 17088 21600 17152
rect 21664 17088 21670 17152
rect 20626 16728 20974 16734
rect 20626 16664 20632 16728
rect 20696 16664 20768 16728
rect 20832 16664 20904 16728
rect 20968 16664 20974 16728
rect 20626 16592 20974 16664
rect 20626 16528 20632 16592
rect 20696 16528 20768 16592
rect 20832 16528 20904 16592
rect 20968 16528 20974 16592
rect 19839 16456 19915 16462
rect 19839 16392 19845 16456
rect 19909 16392 19915 16456
rect 19839 15906 19915 16392
rect 19839 15842 19845 15906
rect 19909 15842 19915 15906
rect 19839 15836 19915 15842
rect 20626 16456 20974 16528
rect 20626 16392 20632 16456
rect 20696 16392 20768 16456
rect 20832 16392 20904 16456
rect 20968 16392 20974 16456
rect 20626 15906 20974 16392
rect 20626 15842 20632 15906
rect 20696 15842 20974 15906
rect 16813 7192 16819 7256
rect 16883 7192 16889 7256
rect 16813 7186 16889 7192
rect 19909 7256 19985 7262
rect 19909 7192 19915 7256
rect 19979 7192 19985 7256
rect 13440 5774 13446 5838
rect 13510 5774 13516 5838
rect 6383 3238 6389 3302
rect 6453 3238 6459 3302
rect 6383 3232 6459 3238
rect 8371 3302 8447 3308
rect 8371 3238 8377 3302
rect 8441 3238 8447 3302
rect 5761 1810 5767 1874
rect 5831 1810 5837 1874
rect 5761 1804 5837 1810
rect 7934 1874 8010 1880
rect 7934 1810 7940 1874
rect 8004 1810 8010 1874
rect 4738 1438 4744 1502
rect 4808 1438 4814 1502
rect 4738 1432 4814 1438
rect 4589 204 4595 268
rect 4659 204 4665 268
rect 4589 198 4665 204
rect 7794 958 7870 964
rect 7794 894 7800 958
rect 7864 894 7870 958
rect 3703 -522 3709 -458
rect 3773 -522 3779 -458
rect 3703 -528 3779 -522
rect 3986 109 4062 115
rect 3986 45 3992 109
rect 4056 45 4062 109
rect 3986 -1496 4062 45
rect 4394 109 4470 115
rect 4394 45 4400 109
rect 4464 45 4470 109
rect 4394 -1496 4470 45
rect 7794 -1154 7870 894
rect 7934 -458 8010 1810
rect 8371 958 8447 3238
rect 8371 894 8377 958
rect 8441 894 8447 958
rect 8371 888 8447 894
rect 12164 1874 12240 1880
rect 12164 1810 12170 1874
rect 12234 1810 12240 1874
rect 7934 -522 7940 -458
rect 8004 -522 8010 -458
rect 7934 -528 8010 -522
rect 8539 439 8615 445
rect 8539 375 8545 439
rect 8609 375 8615 439
rect 7794 -1218 7800 -1154
rect 7864 -1218 7870 -1154
rect 7794 -1224 7870 -1218
rect 8539 -1496 8615 375
rect 8847 439 8923 445
rect 8847 375 8853 439
rect 8917 375 8923 439
rect 8847 -1496 8923 375
rect 9155 439 9231 445
rect 9155 375 9161 439
rect 9225 375 9231 439
rect 9155 -1496 9231 375
rect 9463 439 9539 445
rect 9463 375 9469 439
rect 9533 375 9539 439
rect 9463 -1496 9539 375
rect 9771 439 9847 445
rect 9771 375 9777 439
rect 9841 375 9847 439
rect 9771 -1496 9847 375
rect 10079 439 10155 445
rect 10079 375 10085 439
rect 10149 375 10155 439
rect 10079 -1496 10155 375
rect 10387 439 10463 445
rect 10387 375 10393 439
rect 10457 375 10463 439
rect 10387 -1496 10463 375
rect 10695 439 10771 445
rect 10695 375 10701 439
rect 10765 375 10771 439
rect 10695 -1496 10771 375
rect 12164 -458 12240 1810
rect 13440 1874 13516 5774
rect 13440 1810 13446 1874
rect 13510 1810 13516 1874
rect 13440 1804 13516 1810
rect 16395 1874 16471 1880
rect 16395 1810 16401 1874
rect 16465 1810 16471 1874
rect 12164 -522 12170 -458
rect 12234 -522 12240 -458
rect 12164 -528 12240 -522
rect 12304 958 12380 964
rect 12304 894 12310 958
rect 12374 894 12380 958
rect 12304 -1154 12380 894
rect 16395 -458 16471 1810
rect 16395 -522 16401 -458
rect 16465 -522 16471 -458
rect 16395 -528 16471 -522
rect 16813 958 16889 964
rect 16813 894 16819 958
rect 16883 894 16889 958
rect 12304 -1218 12310 -1154
rect 12374 -1218 12380 -1154
rect 12304 -1224 12380 -1218
rect 16813 -1154 16889 894
rect 16813 -1218 16819 -1154
rect 16883 -1218 16889 -1154
rect 16813 -1224 16889 -1218
rect 19909 -1154 19985 7192
rect 20626 6347 20974 15842
rect 20626 6340 20904 6347
rect 20626 6276 20632 6340
rect 20696 6283 20904 6340
rect 20968 6283 20974 6347
rect 20696 6276 20974 6283
rect 20626 -458 20974 6276
rect 20626 -522 20632 -458
rect 20696 -522 20768 -458
rect 20832 -522 20904 -458
rect 20968 -522 20974 -458
rect 20626 -594 20974 -522
rect 20626 -658 20632 -594
rect 20696 -658 20768 -594
rect 20832 -658 20904 -594
rect 20968 -658 20974 -594
rect 20626 -730 20974 -658
rect 20626 -794 20632 -730
rect 20696 -794 20768 -730
rect 20832 -794 20904 -730
rect 20968 -794 20974 -730
rect 20626 -800 20974 -794
rect 21322 7256 21670 17088
rect 21322 7192 21328 7256
rect 21392 7192 21670 7256
rect 19909 -1218 19915 -1154
rect 19979 -1218 19985 -1154
rect 19909 -1224 19985 -1218
rect 21322 -1154 21670 7192
rect 21322 -1218 21328 -1154
rect 21392 -1218 21464 -1154
rect 21528 -1218 21600 -1154
rect 21664 -1218 21670 -1154
rect 21322 -1290 21670 -1218
rect 21322 -1354 21328 -1290
rect 21392 -1354 21464 -1290
rect 21528 -1354 21600 -1290
rect 21664 -1354 21670 -1290
rect 21322 -1426 21670 -1354
rect 21322 -1490 21328 -1426
rect 21392 -1490 21464 -1426
rect 21528 -1490 21600 -1426
rect 21664 -1490 21670 -1426
rect 21322 -1496 21670 -1490
use sky130_rom_krom_rom_base_array  sky130_rom_krom_rom_base_array_0
timestamp 1581320205
transform 1 0 6869 0 1 7880
box 0 -84 13305 8021
use sky130_rom_krom_rom_bitline_inverter  sky130_rom_krom_rom_bitline_inverter_0
timestamp 1581320207
transform 0 -1 19947 1 0 5978
box 136 -79 1879 13151
use sky130_rom_krom_rom_column_decode  sky130_rom_krom_rom_column_decode_0
timestamp 1581320207
transform 1 0 3262 0 1 0
box -39 44 3513 5257
use sky130_rom_krom_rom_column_mux_array  sky130_rom_krom_rom_column_mux_array_0
timestamp 1581320207
transform 1 0 6917 0 1 2812
box 0 382 13107 3061
use sky130_rom_krom_rom_control_logic  sky130_rom_krom_rom_control_logic_0
timestamp 1581320207
transform 1 0 426 0 1 133
box -36 -49 2632 5306
use sky130_rom_krom_rom_output_buffer  sky130_rom_krom_rom_output_buffer_0
timestamp 1581320207
transform 0 1 8389 -1 0 2172
box 44 -50 1800 2559
use sky130_rom_krom_rom_row_decode  sky130_rom_krom_rom_row_decode_0
timestamp 1581320207
transform 1 0 0 0 1 5469
box -39 44 6775 10465
<< labels >>
rlabel metal4 s 2529 -1496 2605 -1420 4 cs0
port 3 nsew
rlabel metal3 s -1496 1372 -1420 1448 4 clk0
port 5 nsew
rlabel metal4 s 8539 -1496 8615 -1420 4 dout0[0]
port 7 nsew
rlabel metal4 s 8847 -1496 8923 -1420 4 dout0[1]
port 9 nsew
rlabel metal4 s 9155 -1496 9231 -1420 4 dout0[2]
port 11 nsew
rlabel metal4 s 9463 -1496 9539 -1420 4 dout0[3]
port 13 nsew
rlabel metal4 s 9771 -1496 9847 -1420 4 dout0[4]
port 15 nsew
rlabel metal4 s 10079 -1496 10155 -1420 4 dout0[5]
port 17 nsew
rlabel metal4 s 10387 -1496 10463 -1420 4 dout0[6]
port 19 nsew
rlabel metal4 s 10695 -1496 10771 -1420 4 dout0[7]
port 21 nsew
rlabel metal4 s 3565 -1496 3641 -1420 4 addr0[0]
port 23 nsew
rlabel metal4 s 3986 -1496 4062 -1420 4 addr0[1]
port 25 nsew
rlabel metal4 s 4394 -1496 4470 -1420 4 addr0[2]
port 27 nsew
rlabel metal3 s -1496 5508 -1420 5584 4 addr0[3]
port 29 nsew
rlabel metal3 s -1496 5657 -1420 5733 4 addr0[4]
port 31 nsew
rlabel metal3 s -1496 5795 -1420 5871 4 addr0[5]
port 33 nsew
rlabel metal3 s -1496 5214 -1420 5290 4 addr0[6]
port 35 nsew
rlabel metal3 s -1496 5933 -1420 6009 4 addr0[7]
port 37 nsew
rlabel metal3 s -1496 -1496 21670 -1148 4 vccd1
port 39 nsew
rlabel metal3 s -1496 17082 21670 17430 4 vccd1
port 39 nsew
rlabel metal4 s 21322 -1496 21670 17430 4 vccd1
port 39 nsew
rlabel metal4 s -1496 -1496 -1148 17430 4 vccd1
port 39 nsew
rlabel metal4 s -800 -800 -452 16734 4 vssd1
port 41 nsew
rlabel metal3 s -800 16386 20974 16734 4 vssd1
port 41 nsew
rlabel metal3 s -800 -800 20974 -452 4 vssd1
port 41 nsew
rlabel metal4 s 20626 -800 20974 16734 4 vssd1
port 41 nsew
<< properties >>
string FIXED_BBOX 21594 -1491 21670 -1425
<< end >>
