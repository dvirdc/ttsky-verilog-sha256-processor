magic
tech sky130A
magscale 1 2
timestamp 1581321262
<< checkpaint >>
rect -1260 -1344 11301 11529
<< pwell >>
rect 177 9502 9913 9604
rect 177 7766 9913 7868
rect 177 6030 9913 6132
rect 177 4294 9913 4396
rect 177 2558 9913 2660
rect 177 822 9913 924
<< psubdiff >>
rect 203 9570 285 9578
rect 203 9536 227 9570
rect 261 9536 285 9570
rect 203 9528 285 9536
rect 407 9570 489 9578
rect 407 9536 431 9570
rect 465 9536 489 9570
rect 407 9528 489 9536
rect 611 9570 693 9578
rect 611 9536 635 9570
rect 669 9536 693 9570
rect 611 9528 693 9536
rect 815 9570 897 9578
rect 815 9536 839 9570
rect 873 9536 897 9570
rect 815 9528 897 9536
rect 1019 9570 1101 9578
rect 1019 9536 1043 9570
rect 1077 9536 1101 9570
rect 1019 9528 1101 9536
rect 1223 9570 1305 9578
rect 1223 9536 1247 9570
rect 1281 9536 1305 9570
rect 1223 9528 1305 9536
rect 1427 9570 1509 9578
rect 1427 9536 1451 9570
rect 1485 9536 1509 9570
rect 1427 9528 1509 9536
rect 1631 9570 1713 9578
rect 1631 9536 1655 9570
rect 1689 9536 1713 9570
rect 1631 9528 1713 9536
rect 1835 9570 1917 9578
rect 1835 9536 1859 9570
rect 1893 9536 1917 9570
rect 1835 9528 1917 9536
rect 2039 9570 2121 9578
rect 2039 9536 2063 9570
rect 2097 9536 2121 9570
rect 2039 9528 2121 9536
rect 2243 9570 2325 9578
rect 2243 9536 2267 9570
rect 2301 9536 2325 9570
rect 2243 9528 2325 9536
rect 2447 9570 2529 9578
rect 2447 9536 2471 9570
rect 2505 9536 2529 9570
rect 2447 9528 2529 9536
rect 2651 9570 2733 9578
rect 2651 9536 2675 9570
rect 2709 9536 2733 9570
rect 2651 9528 2733 9536
rect 2855 9570 2937 9578
rect 2855 9536 2879 9570
rect 2913 9536 2937 9570
rect 2855 9528 2937 9536
rect 3059 9570 3141 9578
rect 3059 9536 3083 9570
rect 3117 9536 3141 9570
rect 3059 9528 3141 9536
rect 3263 9570 3345 9578
rect 3263 9536 3287 9570
rect 3321 9536 3345 9570
rect 3263 9528 3345 9536
rect 3467 9570 3549 9578
rect 3467 9536 3491 9570
rect 3525 9536 3549 9570
rect 3467 9528 3549 9536
rect 3671 9570 3753 9578
rect 3671 9536 3695 9570
rect 3729 9536 3753 9570
rect 3671 9528 3753 9536
rect 3875 9570 3957 9578
rect 3875 9536 3899 9570
rect 3933 9536 3957 9570
rect 3875 9528 3957 9536
rect 4079 9570 4161 9578
rect 4079 9536 4103 9570
rect 4137 9536 4161 9570
rect 4079 9528 4161 9536
rect 4283 9570 4365 9578
rect 4283 9536 4307 9570
rect 4341 9536 4365 9570
rect 4283 9528 4365 9536
rect 4487 9570 4569 9578
rect 4487 9536 4511 9570
rect 4545 9536 4569 9570
rect 4487 9528 4569 9536
rect 4691 9570 4773 9578
rect 4691 9536 4715 9570
rect 4749 9536 4773 9570
rect 4691 9528 4773 9536
rect 4895 9570 4977 9578
rect 4895 9536 4919 9570
rect 4953 9536 4977 9570
rect 4895 9528 4977 9536
rect 5099 9570 5181 9578
rect 5099 9536 5123 9570
rect 5157 9536 5181 9570
rect 5099 9528 5181 9536
rect 5303 9570 5385 9578
rect 5303 9536 5327 9570
rect 5361 9536 5385 9570
rect 5303 9528 5385 9536
rect 5507 9570 5589 9578
rect 5507 9536 5531 9570
rect 5565 9536 5589 9570
rect 5507 9528 5589 9536
rect 5711 9570 5793 9578
rect 5711 9536 5735 9570
rect 5769 9536 5793 9570
rect 5711 9528 5793 9536
rect 5915 9570 5997 9578
rect 5915 9536 5939 9570
rect 5973 9536 5997 9570
rect 5915 9528 5997 9536
rect 6119 9570 6201 9578
rect 6119 9536 6143 9570
rect 6177 9536 6201 9570
rect 6119 9528 6201 9536
rect 6323 9570 6405 9578
rect 6323 9536 6347 9570
rect 6381 9536 6405 9570
rect 6323 9528 6405 9536
rect 6527 9570 6609 9578
rect 6527 9536 6551 9570
rect 6585 9536 6609 9570
rect 6527 9528 6609 9536
rect 6731 9570 6813 9578
rect 6731 9536 6755 9570
rect 6789 9536 6813 9570
rect 6731 9528 6813 9536
rect 6935 9570 7017 9578
rect 6935 9536 6959 9570
rect 6993 9536 7017 9570
rect 6935 9528 7017 9536
rect 7139 9570 7221 9578
rect 7139 9536 7163 9570
rect 7197 9536 7221 9570
rect 7139 9528 7221 9536
rect 7343 9570 7425 9578
rect 7343 9536 7367 9570
rect 7401 9536 7425 9570
rect 7343 9528 7425 9536
rect 7547 9570 7629 9578
rect 7547 9536 7571 9570
rect 7605 9536 7629 9570
rect 7547 9528 7629 9536
rect 7751 9570 7833 9578
rect 7751 9536 7775 9570
rect 7809 9536 7833 9570
rect 7751 9528 7833 9536
rect 7955 9570 8037 9578
rect 7955 9536 7979 9570
rect 8013 9536 8037 9570
rect 7955 9528 8037 9536
rect 8159 9570 8241 9578
rect 8159 9536 8183 9570
rect 8217 9536 8241 9570
rect 8159 9528 8241 9536
rect 8363 9570 8445 9578
rect 8363 9536 8387 9570
rect 8421 9536 8445 9570
rect 8363 9528 8445 9536
rect 8567 9570 8649 9578
rect 8567 9536 8591 9570
rect 8625 9536 8649 9570
rect 8567 9528 8649 9536
rect 8771 9570 8853 9578
rect 8771 9536 8795 9570
rect 8829 9536 8853 9570
rect 8771 9528 8853 9536
rect 8975 9570 9057 9578
rect 8975 9536 8999 9570
rect 9033 9536 9057 9570
rect 8975 9528 9057 9536
rect 9179 9570 9261 9578
rect 9179 9536 9203 9570
rect 9237 9536 9261 9570
rect 9179 9528 9261 9536
rect 9383 9570 9465 9578
rect 9383 9536 9407 9570
rect 9441 9536 9465 9570
rect 9383 9528 9465 9536
rect 9587 9570 9669 9578
rect 9587 9536 9611 9570
rect 9645 9536 9669 9570
rect 9587 9528 9669 9536
rect 9805 9570 9887 9578
rect 9805 9536 9829 9570
rect 9863 9536 9887 9570
rect 9805 9528 9887 9536
rect 203 7834 285 7842
rect 203 7800 227 7834
rect 261 7800 285 7834
rect 203 7792 285 7800
rect 407 7834 489 7842
rect 407 7800 431 7834
rect 465 7800 489 7834
rect 407 7792 489 7800
rect 611 7834 693 7842
rect 611 7800 635 7834
rect 669 7800 693 7834
rect 611 7792 693 7800
rect 815 7834 897 7842
rect 815 7800 839 7834
rect 873 7800 897 7834
rect 815 7792 897 7800
rect 1019 7834 1101 7842
rect 1019 7800 1043 7834
rect 1077 7800 1101 7834
rect 1019 7792 1101 7800
rect 1223 7834 1305 7842
rect 1223 7800 1247 7834
rect 1281 7800 1305 7834
rect 1223 7792 1305 7800
rect 1427 7834 1509 7842
rect 1427 7800 1451 7834
rect 1485 7800 1509 7834
rect 1427 7792 1509 7800
rect 1631 7834 1713 7842
rect 1631 7800 1655 7834
rect 1689 7800 1713 7834
rect 1631 7792 1713 7800
rect 1835 7834 1917 7842
rect 1835 7800 1859 7834
rect 1893 7800 1917 7834
rect 1835 7792 1917 7800
rect 2039 7834 2121 7842
rect 2039 7800 2063 7834
rect 2097 7800 2121 7834
rect 2039 7792 2121 7800
rect 2243 7834 2325 7842
rect 2243 7800 2267 7834
rect 2301 7800 2325 7834
rect 2243 7792 2325 7800
rect 2447 7834 2529 7842
rect 2447 7800 2471 7834
rect 2505 7800 2529 7834
rect 2447 7792 2529 7800
rect 2651 7834 2733 7842
rect 2651 7800 2675 7834
rect 2709 7800 2733 7834
rect 2651 7792 2733 7800
rect 2855 7834 2937 7842
rect 2855 7800 2879 7834
rect 2913 7800 2937 7834
rect 2855 7792 2937 7800
rect 3059 7834 3141 7842
rect 3059 7800 3083 7834
rect 3117 7800 3141 7834
rect 3059 7792 3141 7800
rect 3263 7834 3345 7842
rect 3263 7800 3287 7834
rect 3321 7800 3345 7834
rect 3263 7792 3345 7800
rect 3467 7834 3549 7842
rect 3467 7800 3491 7834
rect 3525 7800 3549 7834
rect 3467 7792 3549 7800
rect 3671 7834 3753 7842
rect 3671 7800 3695 7834
rect 3729 7800 3753 7834
rect 3671 7792 3753 7800
rect 3875 7834 3957 7842
rect 3875 7800 3899 7834
rect 3933 7800 3957 7834
rect 3875 7792 3957 7800
rect 4079 7834 4161 7842
rect 4079 7800 4103 7834
rect 4137 7800 4161 7834
rect 4079 7792 4161 7800
rect 4283 7834 4365 7842
rect 4283 7800 4307 7834
rect 4341 7800 4365 7834
rect 4283 7792 4365 7800
rect 4487 7834 4569 7842
rect 4487 7800 4511 7834
rect 4545 7800 4569 7834
rect 4487 7792 4569 7800
rect 4691 7834 4773 7842
rect 4691 7800 4715 7834
rect 4749 7800 4773 7834
rect 4691 7792 4773 7800
rect 4895 7834 4977 7842
rect 4895 7800 4919 7834
rect 4953 7800 4977 7834
rect 4895 7792 4977 7800
rect 5099 7834 5181 7842
rect 5099 7800 5123 7834
rect 5157 7800 5181 7834
rect 5099 7792 5181 7800
rect 5303 7834 5385 7842
rect 5303 7800 5327 7834
rect 5361 7800 5385 7834
rect 5303 7792 5385 7800
rect 5507 7834 5589 7842
rect 5507 7800 5531 7834
rect 5565 7800 5589 7834
rect 5507 7792 5589 7800
rect 5711 7834 5793 7842
rect 5711 7800 5735 7834
rect 5769 7800 5793 7834
rect 5711 7792 5793 7800
rect 5915 7834 5997 7842
rect 5915 7800 5939 7834
rect 5973 7800 5997 7834
rect 5915 7792 5997 7800
rect 6119 7834 6201 7842
rect 6119 7800 6143 7834
rect 6177 7800 6201 7834
rect 6119 7792 6201 7800
rect 6323 7834 6405 7842
rect 6323 7800 6347 7834
rect 6381 7800 6405 7834
rect 6323 7792 6405 7800
rect 6527 7834 6609 7842
rect 6527 7800 6551 7834
rect 6585 7800 6609 7834
rect 6527 7792 6609 7800
rect 6731 7834 6813 7842
rect 6731 7800 6755 7834
rect 6789 7800 6813 7834
rect 6731 7792 6813 7800
rect 6935 7834 7017 7842
rect 6935 7800 6959 7834
rect 6993 7800 7017 7834
rect 6935 7792 7017 7800
rect 7139 7834 7221 7842
rect 7139 7800 7163 7834
rect 7197 7800 7221 7834
rect 7139 7792 7221 7800
rect 7343 7834 7425 7842
rect 7343 7800 7367 7834
rect 7401 7800 7425 7834
rect 7343 7792 7425 7800
rect 7547 7834 7629 7842
rect 7547 7800 7571 7834
rect 7605 7800 7629 7834
rect 7547 7792 7629 7800
rect 7751 7834 7833 7842
rect 7751 7800 7775 7834
rect 7809 7800 7833 7834
rect 7751 7792 7833 7800
rect 7955 7834 8037 7842
rect 7955 7800 7979 7834
rect 8013 7800 8037 7834
rect 7955 7792 8037 7800
rect 8159 7834 8241 7842
rect 8159 7800 8183 7834
rect 8217 7800 8241 7834
rect 8159 7792 8241 7800
rect 8363 7834 8445 7842
rect 8363 7800 8387 7834
rect 8421 7800 8445 7834
rect 8363 7792 8445 7800
rect 8567 7834 8649 7842
rect 8567 7800 8591 7834
rect 8625 7800 8649 7834
rect 8567 7792 8649 7800
rect 8771 7834 8853 7842
rect 8771 7800 8795 7834
rect 8829 7800 8853 7834
rect 8771 7792 8853 7800
rect 8975 7834 9057 7842
rect 8975 7800 8999 7834
rect 9033 7800 9057 7834
rect 8975 7792 9057 7800
rect 9179 7834 9261 7842
rect 9179 7800 9203 7834
rect 9237 7800 9261 7834
rect 9179 7792 9261 7800
rect 9383 7834 9465 7842
rect 9383 7800 9407 7834
rect 9441 7800 9465 7834
rect 9383 7792 9465 7800
rect 9587 7834 9669 7842
rect 9587 7800 9611 7834
rect 9645 7800 9669 7834
rect 9587 7792 9669 7800
rect 9805 7834 9887 7842
rect 9805 7800 9829 7834
rect 9863 7800 9887 7834
rect 9805 7792 9887 7800
rect 203 6098 285 6106
rect 203 6064 227 6098
rect 261 6064 285 6098
rect 203 6056 285 6064
rect 407 6098 489 6106
rect 407 6064 431 6098
rect 465 6064 489 6098
rect 407 6056 489 6064
rect 611 6098 693 6106
rect 611 6064 635 6098
rect 669 6064 693 6098
rect 611 6056 693 6064
rect 815 6098 897 6106
rect 815 6064 839 6098
rect 873 6064 897 6098
rect 815 6056 897 6064
rect 1019 6098 1101 6106
rect 1019 6064 1043 6098
rect 1077 6064 1101 6098
rect 1019 6056 1101 6064
rect 1223 6098 1305 6106
rect 1223 6064 1247 6098
rect 1281 6064 1305 6098
rect 1223 6056 1305 6064
rect 1427 6098 1509 6106
rect 1427 6064 1451 6098
rect 1485 6064 1509 6098
rect 1427 6056 1509 6064
rect 1631 6098 1713 6106
rect 1631 6064 1655 6098
rect 1689 6064 1713 6098
rect 1631 6056 1713 6064
rect 1835 6098 1917 6106
rect 1835 6064 1859 6098
rect 1893 6064 1917 6098
rect 1835 6056 1917 6064
rect 2039 6098 2121 6106
rect 2039 6064 2063 6098
rect 2097 6064 2121 6098
rect 2039 6056 2121 6064
rect 2243 6098 2325 6106
rect 2243 6064 2267 6098
rect 2301 6064 2325 6098
rect 2243 6056 2325 6064
rect 2447 6098 2529 6106
rect 2447 6064 2471 6098
rect 2505 6064 2529 6098
rect 2447 6056 2529 6064
rect 2651 6098 2733 6106
rect 2651 6064 2675 6098
rect 2709 6064 2733 6098
rect 2651 6056 2733 6064
rect 2855 6098 2937 6106
rect 2855 6064 2879 6098
rect 2913 6064 2937 6098
rect 2855 6056 2937 6064
rect 3059 6098 3141 6106
rect 3059 6064 3083 6098
rect 3117 6064 3141 6098
rect 3059 6056 3141 6064
rect 3263 6098 3345 6106
rect 3263 6064 3287 6098
rect 3321 6064 3345 6098
rect 3263 6056 3345 6064
rect 3467 6098 3549 6106
rect 3467 6064 3491 6098
rect 3525 6064 3549 6098
rect 3467 6056 3549 6064
rect 3671 6098 3753 6106
rect 3671 6064 3695 6098
rect 3729 6064 3753 6098
rect 3671 6056 3753 6064
rect 3875 6098 3957 6106
rect 3875 6064 3899 6098
rect 3933 6064 3957 6098
rect 3875 6056 3957 6064
rect 4079 6098 4161 6106
rect 4079 6064 4103 6098
rect 4137 6064 4161 6098
rect 4079 6056 4161 6064
rect 4283 6098 4365 6106
rect 4283 6064 4307 6098
rect 4341 6064 4365 6098
rect 4283 6056 4365 6064
rect 4487 6098 4569 6106
rect 4487 6064 4511 6098
rect 4545 6064 4569 6098
rect 4487 6056 4569 6064
rect 4691 6098 4773 6106
rect 4691 6064 4715 6098
rect 4749 6064 4773 6098
rect 4691 6056 4773 6064
rect 4895 6098 4977 6106
rect 4895 6064 4919 6098
rect 4953 6064 4977 6098
rect 4895 6056 4977 6064
rect 5099 6098 5181 6106
rect 5099 6064 5123 6098
rect 5157 6064 5181 6098
rect 5099 6056 5181 6064
rect 5303 6098 5385 6106
rect 5303 6064 5327 6098
rect 5361 6064 5385 6098
rect 5303 6056 5385 6064
rect 5507 6098 5589 6106
rect 5507 6064 5531 6098
rect 5565 6064 5589 6098
rect 5507 6056 5589 6064
rect 5711 6098 5793 6106
rect 5711 6064 5735 6098
rect 5769 6064 5793 6098
rect 5711 6056 5793 6064
rect 5915 6098 5997 6106
rect 5915 6064 5939 6098
rect 5973 6064 5997 6098
rect 5915 6056 5997 6064
rect 6119 6098 6201 6106
rect 6119 6064 6143 6098
rect 6177 6064 6201 6098
rect 6119 6056 6201 6064
rect 6323 6098 6405 6106
rect 6323 6064 6347 6098
rect 6381 6064 6405 6098
rect 6323 6056 6405 6064
rect 6527 6098 6609 6106
rect 6527 6064 6551 6098
rect 6585 6064 6609 6098
rect 6527 6056 6609 6064
rect 6731 6098 6813 6106
rect 6731 6064 6755 6098
rect 6789 6064 6813 6098
rect 6731 6056 6813 6064
rect 6935 6098 7017 6106
rect 6935 6064 6959 6098
rect 6993 6064 7017 6098
rect 6935 6056 7017 6064
rect 7139 6098 7221 6106
rect 7139 6064 7163 6098
rect 7197 6064 7221 6098
rect 7139 6056 7221 6064
rect 7343 6098 7425 6106
rect 7343 6064 7367 6098
rect 7401 6064 7425 6098
rect 7343 6056 7425 6064
rect 7547 6098 7629 6106
rect 7547 6064 7571 6098
rect 7605 6064 7629 6098
rect 7547 6056 7629 6064
rect 7751 6098 7833 6106
rect 7751 6064 7775 6098
rect 7809 6064 7833 6098
rect 7751 6056 7833 6064
rect 7955 6098 8037 6106
rect 7955 6064 7979 6098
rect 8013 6064 8037 6098
rect 7955 6056 8037 6064
rect 8159 6098 8241 6106
rect 8159 6064 8183 6098
rect 8217 6064 8241 6098
rect 8159 6056 8241 6064
rect 8363 6098 8445 6106
rect 8363 6064 8387 6098
rect 8421 6064 8445 6098
rect 8363 6056 8445 6064
rect 8567 6098 8649 6106
rect 8567 6064 8591 6098
rect 8625 6064 8649 6098
rect 8567 6056 8649 6064
rect 8771 6098 8853 6106
rect 8771 6064 8795 6098
rect 8829 6064 8853 6098
rect 8771 6056 8853 6064
rect 8975 6098 9057 6106
rect 8975 6064 8999 6098
rect 9033 6064 9057 6098
rect 8975 6056 9057 6064
rect 9179 6098 9261 6106
rect 9179 6064 9203 6098
rect 9237 6064 9261 6098
rect 9179 6056 9261 6064
rect 9383 6098 9465 6106
rect 9383 6064 9407 6098
rect 9441 6064 9465 6098
rect 9383 6056 9465 6064
rect 9587 6098 9669 6106
rect 9587 6064 9611 6098
rect 9645 6064 9669 6098
rect 9587 6056 9669 6064
rect 9805 6098 9887 6106
rect 9805 6064 9829 6098
rect 9863 6064 9887 6098
rect 9805 6056 9887 6064
rect 203 4362 285 4370
rect 203 4328 227 4362
rect 261 4328 285 4362
rect 203 4320 285 4328
rect 407 4362 489 4370
rect 407 4328 431 4362
rect 465 4328 489 4362
rect 407 4320 489 4328
rect 611 4362 693 4370
rect 611 4328 635 4362
rect 669 4328 693 4362
rect 611 4320 693 4328
rect 815 4362 897 4370
rect 815 4328 839 4362
rect 873 4328 897 4362
rect 815 4320 897 4328
rect 1019 4362 1101 4370
rect 1019 4328 1043 4362
rect 1077 4328 1101 4362
rect 1019 4320 1101 4328
rect 1223 4362 1305 4370
rect 1223 4328 1247 4362
rect 1281 4328 1305 4362
rect 1223 4320 1305 4328
rect 1427 4362 1509 4370
rect 1427 4328 1451 4362
rect 1485 4328 1509 4362
rect 1427 4320 1509 4328
rect 1631 4362 1713 4370
rect 1631 4328 1655 4362
rect 1689 4328 1713 4362
rect 1631 4320 1713 4328
rect 1835 4362 1917 4370
rect 1835 4328 1859 4362
rect 1893 4328 1917 4362
rect 1835 4320 1917 4328
rect 2039 4362 2121 4370
rect 2039 4328 2063 4362
rect 2097 4328 2121 4362
rect 2039 4320 2121 4328
rect 2243 4362 2325 4370
rect 2243 4328 2267 4362
rect 2301 4328 2325 4362
rect 2243 4320 2325 4328
rect 2447 4362 2529 4370
rect 2447 4328 2471 4362
rect 2505 4328 2529 4362
rect 2447 4320 2529 4328
rect 2651 4362 2733 4370
rect 2651 4328 2675 4362
rect 2709 4328 2733 4362
rect 2651 4320 2733 4328
rect 2855 4362 2937 4370
rect 2855 4328 2879 4362
rect 2913 4328 2937 4362
rect 2855 4320 2937 4328
rect 3059 4362 3141 4370
rect 3059 4328 3083 4362
rect 3117 4328 3141 4362
rect 3059 4320 3141 4328
rect 3263 4362 3345 4370
rect 3263 4328 3287 4362
rect 3321 4328 3345 4362
rect 3263 4320 3345 4328
rect 3467 4362 3549 4370
rect 3467 4328 3491 4362
rect 3525 4328 3549 4362
rect 3467 4320 3549 4328
rect 3671 4362 3753 4370
rect 3671 4328 3695 4362
rect 3729 4328 3753 4362
rect 3671 4320 3753 4328
rect 3875 4362 3957 4370
rect 3875 4328 3899 4362
rect 3933 4328 3957 4362
rect 3875 4320 3957 4328
rect 4079 4362 4161 4370
rect 4079 4328 4103 4362
rect 4137 4328 4161 4362
rect 4079 4320 4161 4328
rect 4283 4362 4365 4370
rect 4283 4328 4307 4362
rect 4341 4328 4365 4362
rect 4283 4320 4365 4328
rect 4487 4362 4569 4370
rect 4487 4328 4511 4362
rect 4545 4328 4569 4362
rect 4487 4320 4569 4328
rect 4691 4362 4773 4370
rect 4691 4328 4715 4362
rect 4749 4328 4773 4362
rect 4691 4320 4773 4328
rect 4895 4362 4977 4370
rect 4895 4328 4919 4362
rect 4953 4328 4977 4362
rect 4895 4320 4977 4328
rect 5099 4362 5181 4370
rect 5099 4328 5123 4362
rect 5157 4328 5181 4362
rect 5099 4320 5181 4328
rect 5303 4362 5385 4370
rect 5303 4328 5327 4362
rect 5361 4328 5385 4362
rect 5303 4320 5385 4328
rect 5507 4362 5589 4370
rect 5507 4328 5531 4362
rect 5565 4328 5589 4362
rect 5507 4320 5589 4328
rect 5711 4362 5793 4370
rect 5711 4328 5735 4362
rect 5769 4328 5793 4362
rect 5711 4320 5793 4328
rect 5915 4362 5997 4370
rect 5915 4328 5939 4362
rect 5973 4328 5997 4362
rect 5915 4320 5997 4328
rect 6119 4362 6201 4370
rect 6119 4328 6143 4362
rect 6177 4328 6201 4362
rect 6119 4320 6201 4328
rect 6323 4362 6405 4370
rect 6323 4328 6347 4362
rect 6381 4328 6405 4362
rect 6323 4320 6405 4328
rect 6527 4362 6609 4370
rect 6527 4328 6551 4362
rect 6585 4328 6609 4362
rect 6527 4320 6609 4328
rect 6731 4362 6813 4370
rect 6731 4328 6755 4362
rect 6789 4328 6813 4362
rect 6731 4320 6813 4328
rect 6935 4362 7017 4370
rect 6935 4328 6959 4362
rect 6993 4328 7017 4362
rect 6935 4320 7017 4328
rect 7139 4362 7221 4370
rect 7139 4328 7163 4362
rect 7197 4328 7221 4362
rect 7139 4320 7221 4328
rect 7343 4362 7425 4370
rect 7343 4328 7367 4362
rect 7401 4328 7425 4362
rect 7343 4320 7425 4328
rect 7547 4362 7629 4370
rect 7547 4328 7571 4362
rect 7605 4328 7629 4362
rect 7547 4320 7629 4328
rect 7751 4362 7833 4370
rect 7751 4328 7775 4362
rect 7809 4328 7833 4362
rect 7751 4320 7833 4328
rect 7955 4362 8037 4370
rect 7955 4328 7979 4362
rect 8013 4328 8037 4362
rect 7955 4320 8037 4328
rect 8159 4362 8241 4370
rect 8159 4328 8183 4362
rect 8217 4328 8241 4362
rect 8159 4320 8241 4328
rect 8363 4362 8445 4370
rect 8363 4328 8387 4362
rect 8421 4328 8445 4362
rect 8363 4320 8445 4328
rect 8567 4362 8649 4370
rect 8567 4328 8591 4362
rect 8625 4328 8649 4362
rect 8567 4320 8649 4328
rect 8771 4362 8853 4370
rect 8771 4328 8795 4362
rect 8829 4328 8853 4362
rect 8771 4320 8853 4328
rect 8975 4362 9057 4370
rect 8975 4328 8999 4362
rect 9033 4328 9057 4362
rect 8975 4320 9057 4328
rect 9179 4362 9261 4370
rect 9179 4328 9203 4362
rect 9237 4328 9261 4362
rect 9179 4320 9261 4328
rect 9383 4362 9465 4370
rect 9383 4328 9407 4362
rect 9441 4328 9465 4362
rect 9383 4320 9465 4328
rect 9587 4362 9669 4370
rect 9587 4328 9611 4362
rect 9645 4328 9669 4362
rect 9587 4320 9669 4328
rect 9805 4362 9887 4370
rect 9805 4328 9829 4362
rect 9863 4328 9887 4362
rect 9805 4320 9887 4328
rect 203 2626 285 2634
rect 203 2592 227 2626
rect 261 2592 285 2626
rect 203 2584 285 2592
rect 407 2626 489 2634
rect 407 2592 431 2626
rect 465 2592 489 2626
rect 407 2584 489 2592
rect 611 2626 693 2634
rect 611 2592 635 2626
rect 669 2592 693 2626
rect 611 2584 693 2592
rect 815 2626 897 2634
rect 815 2592 839 2626
rect 873 2592 897 2626
rect 815 2584 897 2592
rect 1019 2626 1101 2634
rect 1019 2592 1043 2626
rect 1077 2592 1101 2626
rect 1019 2584 1101 2592
rect 1223 2626 1305 2634
rect 1223 2592 1247 2626
rect 1281 2592 1305 2626
rect 1223 2584 1305 2592
rect 1427 2626 1509 2634
rect 1427 2592 1451 2626
rect 1485 2592 1509 2626
rect 1427 2584 1509 2592
rect 1631 2626 1713 2634
rect 1631 2592 1655 2626
rect 1689 2592 1713 2626
rect 1631 2584 1713 2592
rect 1835 2626 1917 2634
rect 1835 2592 1859 2626
rect 1893 2592 1917 2626
rect 1835 2584 1917 2592
rect 2039 2626 2121 2634
rect 2039 2592 2063 2626
rect 2097 2592 2121 2626
rect 2039 2584 2121 2592
rect 2243 2626 2325 2634
rect 2243 2592 2267 2626
rect 2301 2592 2325 2626
rect 2243 2584 2325 2592
rect 2447 2626 2529 2634
rect 2447 2592 2471 2626
rect 2505 2592 2529 2626
rect 2447 2584 2529 2592
rect 2651 2626 2733 2634
rect 2651 2592 2675 2626
rect 2709 2592 2733 2626
rect 2651 2584 2733 2592
rect 2855 2626 2937 2634
rect 2855 2592 2879 2626
rect 2913 2592 2937 2626
rect 2855 2584 2937 2592
rect 3059 2626 3141 2634
rect 3059 2592 3083 2626
rect 3117 2592 3141 2626
rect 3059 2584 3141 2592
rect 3263 2626 3345 2634
rect 3263 2592 3287 2626
rect 3321 2592 3345 2626
rect 3263 2584 3345 2592
rect 3467 2626 3549 2634
rect 3467 2592 3491 2626
rect 3525 2592 3549 2626
rect 3467 2584 3549 2592
rect 3671 2626 3753 2634
rect 3671 2592 3695 2626
rect 3729 2592 3753 2626
rect 3671 2584 3753 2592
rect 3875 2626 3957 2634
rect 3875 2592 3899 2626
rect 3933 2592 3957 2626
rect 3875 2584 3957 2592
rect 4079 2626 4161 2634
rect 4079 2592 4103 2626
rect 4137 2592 4161 2626
rect 4079 2584 4161 2592
rect 4283 2626 4365 2634
rect 4283 2592 4307 2626
rect 4341 2592 4365 2626
rect 4283 2584 4365 2592
rect 4487 2626 4569 2634
rect 4487 2592 4511 2626
rect 4545 2592 4569 2626
rect 4487 2584 4569 2592
rect 4691 2626 4773 2634
rect 4691 2592 4715 2626
rect 4749 2592 4773 2626
rect 4691 2584 4773 2592
rect 4895 2626 4977 2634
rect 4895 2592 4919 2626
rect 4953 2592 4977 2626
rect 4895 2584 4977 2592
rect 5099 2626 5181 2634
rect 5099 2592 5123 2626
rect 5157 2592 5181 2626
rect 5099 2584 5181 2592
rect 5303 2626 5385 2634
rect 5303 2592 5327 2626
rect 5361 2592 5385 2626
rect 5303 2584 5385 2592
rect 5507 2626 5589 2634
rect 5507 2592 5531 2626
rect 5565 2592 5589 2626
rect 5507 2584 5589 2592
rect 5711 2626 5793 2634
rect 5711 2592 5735 2626
rect 5769 2592 5793 2626
rect 5711 2584 5793 2592
rect 5915 2626 5997 2634
rect 5915 2592 5939 2626
rect 5973 2592 5997 2626
rect 5915 2584 5997 2592
rect 6119 2626 6201 2634
rect 6119 2592 6143 2626
rect 6177 2592 6201 2626
rect 6119 2584 6201 2592
rect 6323 2626 6405 2634
rect 6323 2592 6347 2626
rect 6381 2592 6405 2626
rect 6323 2584 6405 2592
rect 6527 2626 6609 2634
rect 6527 2592 6551 2626
rect 6585 2592 6609 2626
rect 6527 2584 6609 2592
rect 6731 2626 6813 2634
rect 6731 2592 6755 2626
rect 6789 2592 6813 2626
rect 6731 2584 6813 2592
rect 6935 2626 7017 2634
rect 6935 2592 6959 2626
rect 6993 2592 7017 2626
rect 6935 2584 7017 2592
rect 7139 2626 7221 2634
rect 7139 2592 7163 2626
rect 7197 2592 7221 2626
rect 7139 2584 7221 2592
rect 7343 2626 7425 2634
rect 7343 2592 7367 2626
rect 7401 2592 7425 2626
rect 7343 2584 7425 2592
rect 7547 2626 7629 2634
rect 7547 2592 7571 2626
rect 7605 2592 7629 2626
rect 7547 2584 7629 2592
rect 7751 2626 7833 2634
rect 7751 2592 7775 2626
rect 7809 2592 7833 2626
rect 7751 2584 7833 2592
rect 7955 2626 8037 2634
rect 7955 2592 7979 2626
rect 8013 2592 8037 2626
rect 7955 2584 8037 2592
rect 8159 2626 8241 2634
rect 8159 2592 8183 2626
rect 8217 2592 8241 2626
rect 8159 2584 8241 2592
rect 8363 2626 8445 2634
rect 8363 2592 8387 2626
rect 8421 2592 8445 2626
rect 8363 2584 8445 2592
rect 8567 2626 8649 2634
rect 8567 2592 8591 2626
rect 8625 2592 8649 2626
rect 8567 2584 8649 2592
rect 8771 2626 8853 2634
rect 8771 2592 8795 2626
rect 8829 2592 8853 2626
rect 8771 2584 8853 2592
rect 8975 2626 9057 2634
rect 8975 2592 8999 2626
rect 9033 2592 9057 2626
rect 8975 2584 9057 2592
rect 9179 2626 9261 2634
rect 9179 2592 9203 2626
rect 9237 2592 9261 2626
rect 9179 2584 9261 2592
rect 9383 2626 9465 2634
rect 9383 2592 9407 2626
rect 9441 2592 9465 2626
rect 9383 2584 9465 2592
rect 9587 2626 9669 2634
rect 9587 2592 9611 2626
rect 9645 2592 9669 2626
rect 9587 2584 9669 2592
rect 9805 2626 9887 2634
rect 9805 2592 9829 2626
rect 9863 2592 9887 2626
rect 9805 2584 9887 2592
rect 203 890 285 898
rect 203 856 227 890
rect 261 856 285 890
rect 203 848 285 856
rect 407 890 489 898
rect 407 856 431 890
rect 465 856 489 890
rect 407 848 489 856
rect 611 890 693 898
rect 611 856 635 890
rect 669 856 693 890
rect 611 848 693 856
rect 815 890 897 898
rect 815 856 839 890
rect 873 856 897 890
rect 815 848 897 856
rect 1019 890 1101 898
rect 1019 856 1043 890
rect 1077 856 1101 890
rect 1019 848 1101 856
rect 1223 890 1305 898
rect 1223 856 1247 890
rect 1281 856 1305 890
rect 1223 848 1305 856
rect 1427 890 1509 898
rect 1427 856 1451 890
rect 1485 856 1509 890
rect 1427 848 1509 856
rect 1631 890 1713 898
rect 1631 856 1655 890
rect 1689 856 1713 890
rect 1631 848 1713 856
rect 1835 890 1917 898
rect 1835 856 1859 890
rect 1893 856 1917 890
rect 1835 848 1917 856
rect 2039 890 2121 898
rect 2039 856 2063 890
rect 2097 856 2121 890
rect 2039 848 2121 856
rect 2243 890 2325 898
rect 2243 856 2267 890
rect 2301 856 2325 890
rect 2243 848 2325 856
rect 2447 890 2529 898
rect 2447 856 2471 890
rect 2505 856 2529 890
rect 2447 848 2529 856
rect 2651 890 2733 898
rect 2651 856 2675 890
rect 2709 856 2733 890
rect 2651 848 2733 856
rect 2855 890 2937 898
rect 2855 856 2879 890
rect 2913 856 2937 890
rect 2855 848 2937 856
rect 3059 890 3141 898
rect 3059 856 3083 890
rect 3117 856 3141 890
rect 3059 848 3141 856
rect 3263 890 3345 898
rect 3263 856 3287 890
rect 3321 856 3345 890
rect 3263 848 3345 856
rect 3467 890 3549 898
rect 3467 856 3491 890
rect 3525 856 3549 890
rect 3467 848 3549 856
rect 3671 890 3753 898
rect 3671 856 3695 890
rect 3729 856 3753 890
rect 3671 848 3753 856
rect 3875 890 3957 898
rect 3875 856 3899 890
rect 3933 856 3957 890
rect 3875 848 3957 856
rect 4079 890 4161 898
rect 4079 856 4103 890
rect 4137 856 4161 890
rect 4079 848 4161 856
rect 4283 890 4365 898
rect 4283 856 4307 890
rect 4341 856 4365 890
rect 4283 848 4365 856
rect 4487 890 4569 898
rect 4487 856 4511 890
rect 4545 856 4569 890
rect 4487 848 4569 856
rect 4691 890 4773 898
rect 4691 856 4715 890
rect 4749 856 4773 890
rect 4691 848 4773 856
rect 4895 890 4977 898
rect 4895 856 4919 890
rect 4953 856 4977 890
rect 4895 848 4977 856
rect 5099 890 5181 898
rect 5099 856 5123 890
rect 5157 856 5181 890
rect 5099 848 5181 856
rect 5303 890 5385 898
rect 5303 856 5327 890
rect 5361 856 5385 890
rect 5303 848 5385 856
rect 5507 890 5589 898
rect 5507 856 5531 890
rect 5565 856 5589 890
rect 5507 848 5589 856
rect 5711 890 5793 898
rect 5711 856 5735 890
rect 5769 856 5793 890
rect 5711 848 5793 856
rect 5915 890 5997 898
rect 5915 856 5939 890
rect 5973 856 5997 890
rect 5915 848 5997 856
rect 6119 890 6201 898
rect 6119 856 6143 890
rect 6177 856 6201 890
rect 6119 848 6201 856
rect 6323 890 6405 898
rect 6323 856 6347 890
rect 6381 856 6405 890
rect 6323 848 6405 856
rect 6527 890 6609 898
rect 6527 856 6551 890
rect 6585 856 6609 890
rect 6527 848 6609 856
rect 6731 890 6813 898
rect 6731 856 6755 890
rect 6789 856 6813 890
rect 6731 848 6813 856
rect 6935 890 7017 898
rect 6935 856 6959 890
rect 6993 856 7017 890
rect 6935 848 7017 856
rect 7139 890 7221 898
rect 7139 856 7163 890
rect 7197 856 7221 890
rect 7139 848 7221 856
rect 7343 890 7425 898
rect 7343 856 7367 890
rect 7401 856 7425 890
rect 7343 848 7425 856
rect 7547 890 7629 898
rect 7547 856 7571 890
rect 7605 856 7629 890
rect 7547 848 7629 856
rect 7751 890 7833 898
rect 7751 856 7775 890
rect 7809 856 7833 890
rect 7751 848 7833 856
rect 7955 890 8037 898
rect 7955 856 7979 890
rect 8013 856 8037 890
rect 7955 848 8037 856
rect 8159 890 8241 898
rect 8159 856 8183 890
rect 8217 856 8241 890
rect 8159 848 8241 856
rect 8363 890 8445 898
rect 8363 856 8387 890
rect 8421 856 8445 890
rect 8363 848 8445 856
rect 8567 890 8649 898
rect 8567 856 8591 890
rect 8625 856 8649 890
rect 8567 848 8649 856
rect 8771 890 8853 898
rect 8771 856 8795 890
rect 8829 856 8853 890
rect 8771 848 8853 856
rect 8975 890 9057 898
rect 8975 856 8999 890
rect 9033 856 9057 890
rect 8975 848 9057 856
rect 9179 890 9261 898
rect 9179 856 9203 890
rect 9237 856 9261 890
rect 9179 848 9261 856
rect 9383 890 9465 898
rect 9383 856 9407 890
rect 9441 856 9465 890
rect 9383 848 9465 856
rect 9587 890 9669 898
rect 9587 856 9611 890
rect 9645 856 9669 890
rect 9587 848 9669 856
rect 9805 890 9887 898
rect 9805 856 9829 890
rect 9863 856 9887 890
rect 9805 848 9887 856
<< psubdiffcont >>
rect 227 9536 261 9570
rect 431 9536 465 9570
rect 635 9536 669 9570
rect 839 9536 873 9570
rect 1043 9536 1077 9570
rect 1247 9536 1281 9570
rect 1451 9536 1485 9570
rect 1655 9536 1689 9570
rect 1859 9536 1893 9570
rect 2063 9536 2097 9570
rect 2267 9536 2301 9570
rect 2471 9536 2505 9570
rect 2675 9536 2709 9570
rect 2879 9536 2913 9570
rect 3083 9536 3117 9570
rect 3287 9536 3321 9570
rect 3491 9536 3525 9570
rect 3695 9536 3729 9570
rect 3899 9536 3933 9570
rect 4103 9536 4137 9570
rect 4307 9536 4341 9570
rect 4511 9536 4545 9570
rect 4715 9536 4749 9570
rect 4919 9536 4953 9570
rect 5123 9536 5157 9570
rect 5327 9536 5361 9570
rect 5531 9536 5565 9570
rect 5735 9536 5769 9570
rect 5939 9536 5973 9570
rect 6143 9536 6177 9570
rect 6347 9536 6381 9570
rect 6551 9536 6585 9570
rect 6755 9536 6789 9570
rect 6959 9536 6993 9570
rect 7163 9536 7197 9570
rect 7367 9536 7401 9570
rect 7571 9536 7605 9570
rect 7775 9536 7809 9570
rect 7979 9536 8013 9570
rect 8183 9536 8217 9570
rect 8387 9536 8421 9570
rect 8591 9536 8625 9570
rect 8795 9536 8829 9570
rect 8999 9536 9033 9570
rect 9203 9536 9237 9570
rect 9407 9536 9441 9570
rect 9611 9536 9645 9570
rect 9829 9536 9863 9570
rect 227 7800 261 7834
rect 431 7800 465 7834
rect 635 7800 669 7834
rect 839 7800 873 7834
rect 1043 7800 1077 7834
rect 1247 7800 1281 7834
rect 1451 7800 1485 7834
rect 1655 7800 1689 7834
rect 1859 7800 1893 7834
rect 2063 7800 2097 7834
rect 2267 7800 2301 7834
rect 2471 7800 2505 7834
rect 2675 7800 2709 7834
rect 2879 7800 2913 7834
rect 3083 7800 3117 7834
rect 3287 7800 3321 7834
rect 3491 7800 3525 7834
rect 3695 7800 3729 7834
rect 3899 7800 3933 7834
rect 4103 7800 4137 7834
rect 4307 7800 4341 7834
rect 4511 7800 4545 7834
rect 4715 7800 4749 7834
rect 4919 7800 4953 7834
rect 5123 7800 5157 7834
rect 5327 7800 5361 7834
rect 5531 7800 5565 7834
rect 5735 7800 5769 7834
rect 5939 7800 5973 7834
rect 6143 7800 6177 7834
rect 6347 7800 6381 7834
rect 6551 7800 6585 7834
rect 6755 7800 6789 7834
rect 6959 7800 6993 7834
rect 7163 7800 7197 7834
rect 7367 7800 7401 7834
rect 7571 7800 7605 7834
rect 7775 7800 7809 7834
rect 7979 7800 8013 7834
rect 8183 7800 8217 7834
rect 8387 7800 8421 7834
rect 8591 7800 8625 7834
rect 8795 7800 8829 7834
rect 8999 7800 9033 7834
rect 9203 7800 9237 7834
rect 9407 7800 9441 7834
rect 9611 7800 9645 7834
rect 9829 7800 9863 7834
rect 227 6064 261 6098
rect 431 6064 465 6098
rect 635 6064 669 6098
rect 839 6064 873 6098
rect 1043 6064 1077 6098
rect 1247 6064 1281 6098
rect 1451 6064 1485 6098
rect 1655 6064 1689 6098
rect 1859 6064 1893 6098
rect 2063 6064 2097 6098
rect 2267 6064 2301 6098
rect 2471 6064 2505 6098
rect 2675 6064 2709 6098
rect 2879 6064 2913 6098
rect 3083 6064 3117 6098
rect 3287 6064 3321 6098
rect 3491 6064 3525 6098
rect 3695 6064 3729 6098
rect 3899 6064 3933 6098
rect 4103 6064 4137 6098
rect 4307 6064 4341 6098
rect 4511 6064 4545 6098
rect 4715 6064 4749 6098
rect 4919 6064 4953 6098
rect 5123 6064 5157 6098
rect 5327 6064 5361 6098
rect 5531 6064 5565 6098
rect 5735 6064 5769 6098
rect 5939 6064 5973 6098
rect 6143 6064 6177 6098
rect 6347 6064 6381 6098
rect 6551 6064 6585 6098
rect 6755 6064 6789 6098
rect 6959 6064 6993 6098
rect 7163 6064 7197 6098
rect 7367 6064 7401 6098
rect 7571 6064 7605 6098
rect 7775 6064 7809 6098
rect 7979 6064 8013 6098
rect 8183 6064 8217 6098
rect 8387 6064 8421 6098
rect 8591 6064 8625 6098
rect 8795 6064 8829 6098
rect 8999 6064 9033 6098
rect 9203 6064 9237 6098
rect 9407 6064 9441 6098
rect 9611 6064 9645 6098
rect 9829 6064 9863 6098
rect 227 4328 261 4362
rect 431 4328 465 4362
rect 635 4328 669 4362
rect 839 4328 873 4362
rect 1043 4328 1077 4362
rect 1247 4328 1281 4362
rect 1451 4328 1485 4362
rect 1655 4328 1689 4362
rect 1859 4328 1893 4362
rect 2063 4328 2097 4362
rect 2267 4328 2301 4362
rect 2471 4328 2505 4362
rect 2675 4328 2709 4362
rect 2879 4328 2913 4362
rect 3083 4328 3117 4362
rect 3287 4328 3321 4362
rect 3491 4328 3525 4362
rect 3695 4328 3729 4362
rect 3899 4328 3933 4362
rect 4103 4328 4137 4362
rect 4307 4328 4341 4362
rect 4511 4328 4545 4362
rect 4715 4328 4749 4362
rect 4919 4328 4953 4362
rect 5123 4328 5157 4362
rect 5327 4328 5361 4362
rect 5531 4328 5565 4362
rect 5735 4328 5769 4362
rect 5939 4328 5973 4362
rect 6143 4328 6177 4362
rect 6347 4328 6381 4362
rect 6551 4328 6585 4362
rect 6755 4328 6789 4362
rect 6959 4328 6993 4362
rect 7163 4328 7197 4362
rect 7367 4328 7401 4362
rect 7571 4328 7605 4362
rect 7775 4328 7809 4362
rect 7979 4328 8013 4362
rect 8183 4328 8217 4362
rect 8387 4328 8421 4362
rect 8591 4328 8625 4362
rect 8795 4328 8829 4362
rect 8999 4328 9033 4362
rect 9203 4328 9237 4362
rect 9407 4328 9441 4362
rect 9611 4328 9645 4362
rect 9829 4328 9863 4362
rect 227 2592 261 2626
rect 431 2592 465 2626
rect 635 2592 669 2626
rect 839 2592 873 2626
rect 1043 2592 1077 2626
rect 1247 2592 1281 2626
rect 1451 2592 1485 2626
rect 1655 2592 1689 2626
rect 1859 2592 1893 2626
rect 2063 2592 2097 2626
rect 2267 2592 2301 2626
rect 2471 2592 2505 2626
rect 2675 2592 2709 2626
rect 2879 2592 2913 2626
rect 3083 2592 3117 2626
rect 3287 2592 3321 2626
rect 3491 2592 3525 2626
rect 3695 2592 3729 2626
rect 3899 2592 3933 2626
rect 4103 2592 4137 2626
rect 4307 2592 4341 2626
rect 4511 2592 4545 2626
rect 4715 2592 4749 2626
rect 4919 2592 4953 2626
rect 5123 2592 5157 2626
rect 5327 2592 5361 2626
rect 5531 2592 5565 2626
rect 5735 2592 5769 2626
rect 5939 2592 5973 2626
rect 6143 2592 6177 2626
rect 6347 2592 6381 2626
rect 6551 2592 6585 2626
rect 6755 2592 6789 2626
rect 6959 2592 6993 2626
rect 7163 2592 7197 2626
rect 7367 2592 7401 2626
rect 7571 2592 7605 2626
rect 7775 2592 7809 2626
rect 7979 2592 8013 2626
rect 8183 2592 8217 2626
rect 8387 2592 8421 2626
rect 8591 2592 8625 2626
rect 8795 2592 8829 2626
rect 8999 2592 9033 2626
rect 9203 2592 9237 2626
rect 9407 2592 9441 2626
rect 9611 2592 9645 2626
rect 9829 2592 9863 2626
rect 227 856 261 890
rect 431 856 465 890
rect 635 856 669 890
rect 839 856 873 890
rect 1043 856 1077 890
rect 1247 856 1281 890
rect 1451 856 1485 890
rect 1655 856 1689 890
rect 1859 856 1893 890
rect 2063 856 2097 890
rect 2267 856 2301 890
rect 2471 856 2505 890
rect 2675 856 2709 890
rect 2879 856 2913 890
rect 3083 856 3117 890
rect 3287 856 3321 890
rect 3491 856 3525 890
rect 3695 856 3729 890
rect 3899 856 3933 890
rect 4103 856 4137 890
rect 4307 856 4341 890
rect 4511 856 4545 890
rect 4715 856 4749 890
rect 4919 856 4953 890
rect 5123 856 5157 890
rect 5327 856 5361 890
rect 5531 856 5565 890
rect 5735 856 5769 890
rect 5939 856 5973 890
rect 6143 856 6177 890
rect 6347 856 6381 890
rect 6551 856 6585 890
rect 6755 856 6789 890
rect 6959 856 6993 890
rect 7163 856 7197 890
rect 7367 856 7401 890
rect 7571 856 7605 890
rect 7775 856 7809 890
rect 7979 856 8013 890
rect 8183 856 8217 890
rect 8387 856 8421 890
rect 8591 856 8625 890
rect 8795 856 8829 890
rect 8999 856 9033 890
rect 9203 856 9237 890
rect 9407 856 9441 890
rect 9611 856 9645 890
rect 9829 856 9863 890
<< poly >>
rect 0 10132 66 10148
rect 0 10098 16 10132
rect 50 10130 66 10132
rect 1632 10132 1698 10148
rect 1632 10130 1648 10132
rect 50 10100 1648 10130
rect 50 10098 66 10100
rect 0 10082 66 10098
rect 1632 10098 1648 10100
rect 1682 10130 1698 10132
rect 3264 10132 3330 10148
rect 3264 10130 3280 10132
rect 1682 10100 3280 10130
rect 1682 10098 1698 10100
rect 1632 10082 1698 10098
rect 3264 10098 3280 10100
rect 3314 10130 3330 10132
rect 4896 10132 4962 10148
rect 4896 10130 4912 10132
rect 3314 10100 4912 10130
rect 3314 10098 3330 10100
rect 3264 10082 3330 10098
rect 4896 10098 4912 10100
rect 4946 10130 4962 10132
rect 6528 10132 6594 10148
rect 6528 10130 6544 10132
rect 4946 10100 6544 10130
rect 4946 10098 4962 10100
rect 4896 10082 4962 10098
rect 6528 10098 6544 10100
rect 6578 10130 6594 10132
rect 8160 10132 8226 10148
rect 8160 10130 8176 10132
rect 6578 10100 8176 10130
rect 6578 10098 6594 10100
rect 6528 10082 6594 10098
rect 8160 10098 8176 10100
rect 8210 10130 8226 10132
rect 9792 10132 9858 10148
rect 9792 10130 9808 10132
rect 8210 10100 9808 10130
rect 8210 10098 8226 10100
rect 8160 10082 8226 10098
rect 9792 10098 9808 10100
rect 9842 10098 9858 10132
rect 9792 10082 9858 10098
rect 0 9928 66 9944
rect 0 9894 16 9928
rect 50 9926 66 9928
rect 1632 9928 1698 9944
rect 1632 9926 1648 9928
rect 50 9896 1648 9926
rect 50 9894 66 9896
rect 0 9878 66 9894
rect 1632 9894 1648 9896
rect 1682 9926 1698 9928
rect 3264 9928 3330 9944
rect 3264 9926 3280 9928
rect 1682 9896 3280 9926
rect 1682 9894 1698 9896
rect 1632 9878 1698 9894
rect 3264 9894 3280 9896
rect 3314 9926 3330 9928
rect 4896 9928 4962 9944
rect 4896 9926 4912 9928
rect 3314 9896 4912 9926
rect 3314 9894 3330 9896
rect 3264 9878 3330 9894
rect 4896 9894 4912 9896
rect 4946 9926 4962 9928
rect 6528 9928 6594 9944
rect 6528 9926 6544 9928
rect 4946 9896 6544 9926
rect 4946 9894 4962 9896
rect 4896 9878 4962 9894
rect 6528 9894 6544 9896
rect 6578 9926 6594 9928
rect 8160 9928 8226 9944
rect 8160 9926 8176 9928
rect 6578 9896 8176 9926
rect 6578 9894 6594 9896
rect 6528 9878 6594 9894
rect 8160 9894 8176 9896
rect 8210 9926 8226 9928
rect 9792 9928 9858 9944
rect 9792 9926 9808 9928
rect 8210 9896 9808 9926
rect 8210 9894 8226 9896
rect 8160 9878 8226 9894
rect 9792 9894 9808 9896
rect 9842 9894 9858 9928
rect 9792 9878 9858 9894
rect 0 9724 66 9740
rect 0 9690 16 9724
rect 50 9722 66 9724
rect 1632 9724 1698 9740
rect 1632 9722 1648 9724
rect 50 9692 1648 9722
rect 50 9690 66 9692
rect 0 9674 66 9690
rect 1632 9690 1648 9692
rect 1682 9722 1698 9724
rect 3264 9724 3330 9740
rect 3264 9722 3280 9724
rect 1682 9692 3280 9722
rect 1682 9690 1698 9692
rect 1632 9674 1698 9690
rect 3264 9690 3280 9692
rect 3314 9722 3330 9724
rect 4896 9724 4962 9740
rect 4896 9722 4912 9724
rect 3314 9692 4912 9722
rect 3314 9690 3330 9692
rect 3264 9674 3330 9690
rect 4896 9690 4912 9692
rect 4946 9722 4962 9724
rect 6528 9724 6594 9740
rect 6528 9722 6544 9724
rect 4946 9692 6544 9722
rect 4946 9690 4962 9692
rect 4896 9674 4962 9690
rect 6528 9690 6544 9692
rect 6578 9722 6594 9724
rect 8160 9724 8226 9740
rect 8160 9722 8176 9724
rect 6578 9692 8176 9722
rect 6578 9690 6594 9692
rect 6528 9674 6594 9690
rect 8160 9690 8176 9692
rect 8210 9722 8226 9724
rect 9792 9724 9858 9740
rect 9792 9722 9808 9724
rect 8210 9692 9808 9722
rect 8210 9690 8226 9692
rect 8160 9674 8226 9690
rect 9792 9690 9808 9692
rect 9842 9690 9858 9724
rect 9792 9674 9858 9690
rect 0 9416 66 9432
rect 0 9382 16 9416
rect 50 9414 66 9416
rect 1632 9416 1698 9432
rect 1632 9414 1648 9416
rect 50 9384 1648 9414
rect 50 9382 66 9384
rect 0 9366 66 9382
rect 1632 9382 1648 9384
rect 1682 9414 1698 9416
rect 3264 9416 3330 9432
rect 3264 9414 3280 9416
rect 1682 9384 3280 9414
rect 1682 9382 1698 9384
rect 1632 9366 1698 9382
rect 3264 9382 3280 9384
rect 3314 9414 3330 9416
rect 4896 9416 4962 9432
rect 4896 9414 4912 9416
rect 3314 9384 4912 9414
rect 3314 9382 3330 9384
rect 3264 9366 3330 9382
rect 4896 9382 4912 9384
rect 4946 9414 4962 9416
rect 6528 9416 6594 9432
rect 6528 9414 6544 9416
rect 4946 9384 6544 9414
rect 4946 9382 4962 9384
rect 4896 9366 4962 9382
rect 6528 9382 6544 9384
rect 6578 9414 6594 9416
rect 8160 9416 8226 9432
rect 8160 9414 8176 9416
rect 6578 9384 8176 9414
rect 6578 9382 6594 9384
rect 6528 9366 6594 9382
rect 8160 9382 8176 9384
rect 8210 9414 8226 9416
rect 9792 9416 9858 9432
rect 9792 9414 9808 9416
rect 8210 9384 9808 9414
rect 8210 9382 8226 9384
rect 8160 9366 8226 9382
rect 9792 9382 9808 9384
rect 9842 9382 9858 9416
rect 9792 9366 9858 9382
rect 0 9212 66 9228
rect 0 9178 16 9212
rect 50 9210 66 9212
rect 1632 9212 1698 9228
rect 1632 9210 1648 9212
rect 50 9180 1648 9210
rect 50 9178 66 9180
rect 0 9162 66 9178
rect 1632 9178 1648 9180
rect 1682 9210 1698 9212
rect 3264 9212 3330 9228
rect 3264 9210 3280 9212
rect 1682 9180 3280 9210
rect 1682 9178 1698 9180
rect 1632 9162 1698 9178
rect 3264 9178 3280 9180
rect 3314 9210 3330 9212
rect 4896 9212 4962 9228
rect 4896 9210 4912 9212
rect 3314 9180 4912 9210
rect 3314 9178 3330 9180
rect 3264 9162 3330 9178
rect 4896 9178 4912 9180
rect 4946 9210 4962 9212
rect 6528 9212 6594 9228
rect 6528 9210 6544 9212
rect 4946 9180 6544 9210
rect 4946 9178 4962 9180
rect 4896 9162 4962 9178
rect 6528 9178 6544 9180
rect 6578 9210 6594 9212
rect 8160 9212 8226 9228
rect 8160 9210 8176 9212
rect 6578 9180 8176 9210
rect 6578 9178 6594 9180
rect 6528 9162 6594 9178
rect 8160 9178 8176 9180
rect 8210 9210 8226 9212
rect 9792 9212 9858 9228
rect 9792 9210 9808 9212
rect 8210 9180 9808 9210
rect 8210 9178 8226 9180
rect 8160 9162 8226 9178
rect 9792 9178 9808 9180
rect 9842 9178 9858 9212
rect 9792 9162 9858 9178
rect 0 9008 66 9024
rect 0 8974 16 9008
rect 50 9006 66 9008
rect 1632 9008 1698 9024
rect 1632 9006 1648 9008
rect 50 8976 1648 9006
rect 50 8974 66 8976
rect 0 8958 66 8974
rect 1632 8974 1648 8976
rect 1682 9006 1698 9008
rect 3264 9008 3330 9024
rect 3264 9006 3280 9008
rect 1682 8976 3280 9006
rect 1682 8974 1698 8976
rect 1632 8958 1698 8974
rect 3264 8974 3280 8976
rect 3314 9006 3330 9008
rect 4896 9008 4962 9024
rect 4896 9006 4912 9008
rect 3314 8976 4912 9006
rect 3314 8974 3330 8976
rect 3264 8958 3330 8974
rect 4896 8974 4912 8976
rect 4946 9006 4962 9008
rect 6528 9008 6594 9024
rect 6528 9006 6544 9008
rect 4946 8976 6544 9006
rect 4946 8974 4962 8976
rect 4896 8958 4962 8974
rect 6528 8974 6544 8976
rect 6578 9006 6594 9008
rect 8160 9008 8226 9024
rect 8160 9006 8176 9008
rect 6578 8976 8176 9006
rect 6578 8974 6594 8976
rect 6528 8958 6594 8974
rect 8160 8974 8176 8976
rect 8210 9006 8226 9008
rect 9792 9008 9858 9024
rect 9792 9006 9808 9008
rect 8210 8976 9808 9006
rect 8210 8974 8226 8976
rect 8160 8958 8226 8974
rect 9792 8974 9808 8976
rect 9842 8974 9858 9008
rect 9792 8958 9858 8974
rect 0 8804 66 8820
rect 0 8770 16 8804
rect 50 8802 66 8804
rect 1632 8804 1698 8820
rect 1632 8802 1648 8804
rect 50 8772 1648 8802
rect 50 8770 66 8772
rect 0 8754 66 8770
rect 1632 8770 1648 8772
rect 1682 8802 1698 8804
rect 3264 8804 3330 8820
rect 3264 8802 3280 8804
rect 1682 8772 3280 8802
rect 1682 8770 1698 8772
rect 1632 8754 1698 8770
rect 3264 8770 3280 8772
rect 3314 8802 3330 8804
rect 4896 8804 4962 8820
rect 4896 8802 4912 8804
rect 3314 8772 4912 8802
rect 3314 8770 3330 8772
rect 3264 8754 3330 8770
rect 4896 8770 4912 8772
rect 4946 8802 4962 8804
rect 6528 8804 6594 8820
rect 6528 8802 6544 8804
rect 4946 8772 6544 8802
rect 4946 8770 4962 8772
rect 4896 8754 4962 8770
rect 6528 8770 6544 8772
rect 6578 8802 6594 8804
rect 8160 8804 8226 8820
rect 8160 8802 8176 8804
rect 6578 8772 8176 8802
rect 6578 8770 6594 8772
rect 6528 8754 6594 8770
rect 8160 8770 8176 8772
rect 8210 8802 8226 8804
rect 9792 8804 9858 8820
rect 9792 8802 9808 8804
rect 8210 8772 9808 8802
rect 8210 8770 8226 8772
rect 8160 8754 8226 8770
rect 9792 8770 9808 8772
rect 9842 8770 9858 8804
rect 9792 8754 9858 8770
rect 0 8600 66 8616
rect 0 8566 16 8600
rect 50 8598 66 8600
rect 1632 8600 1698 8616
rect 1632 8598 1648 8600
rect 50 8568 1648 8598
rect 50 8566 66 8568
rect 0 8550 66 8566
rect 1632 8566 1648 8568
rect 1682 8598 1698 8600
rect 3264 8600 3330 8616
rect 3264 8598 3280 8600
rect 1682 8568 3280 8598
rect 1682 8566 1698 8568
rect 1632 8550 1698 8566
rect 3264 8566 3280 8568
rect 3314 8598 3330 8600
rect 4896 8600 4962 8616
rect 4896 8598 4912 8600
rect 3314 8568 4912 8598
rect 3314 8566 3330 8568
rect 3264 8550 3330 8566
rect 4896 8566 4912 8568
rect 4946 8598 4962 8600
rect 6528 8600 6594 8616
rect 6528 8598 6544 8600
rect 4946 8568 6544 8598
rect 4946 8566 4962 8568
rect 4896 8550 4962 8566
rect 6528 8566 6544 8568
rect 6578 8598 6594 8600
rect 8160 8600 8226 8616
rect 8160 8598 8176 8600
rect 6578 8568 8176 8598
rect 6578 8566 6594 8568
rect 6528 8550 6594 8566
rect 8160 8566 8176 8568
rect 8210 8598 8226 8600
rect 9792 8600 9858 8616
rect 9792 8598 9808 8600
rect 8210 8568 9808 8598
rect 8210 8566 8226 8568
rect 8160 8550 8226 8566
rect 9792 8566 9808 8568
rect 9842 8566 9858 8600
rect 9792 8550 9858 8566
rect 0 8396 66 8412
rect 0 8362 16 8396
rect 50 8394 66 8396
rect 1632 8396 1698 8412
rect 1632 8394 1648 8396
rect 50 8364 1648 8394
rect 50 8362 66 8364
rect 0 8346 66 8362
rect 1632 8362 1648 8364
rect 1682 8394 1698 8396
rect 3264 8396 3330 8412
rect 3264 8394 3280 8396
rect 1682 8364 3280 8394
rect 1682 8362 1698 8364
rect 1632 8346 1698 8362
rect 3264 8362 3280 8364
rect 3314 8394 3330 8396
rect 4896 8396 4962 8412
rect 4896 8394 4912 8396
rect 3314 8364 4912 8394
rect 3314 8362 3330 8364
rect 3264 8346 3330 8362
rect 4896 8362 4912 8364
rect 4946 8394 4962 8396
rect 6528 8396 6594 8412
rect 6528 8394 6544 8396
rect 4946 8364 6544 8394
rect 4946 8362 4962 8364
rect 4896 8346 4962 8362
rect 6528 8362 6544 8364
rect 6578 8394 6594 8396
rect 8160 8396 8226 8412
rect 8160 8394 8176 8396
rect 6578 8364 8176 8394
rect 6578 8362 6594 8364
rect 6528 8346 6594 8362
rect 8160 8362 8176 8364
rect 8210 8394 8226 8396
rect 9792 8396 9858 8412
rect 9792 8394 9808 8396
rect 8210 8364 9808 8394
rect 8210 8362 8226 8364
rect 8160 8346 8226 8362
rect 9792 8362 9808 8364
rect 9842 8362 9858 8396
rect 9792 8346 9858 8362
rect 0 8192 66 8208
rect 0 8158 16 8192
rect 50 8190 66 8192
rect 1632 8192 1698 8208
rect 1632 8190 1648 8192
rect 50 8160 1648 8190
rect 50 8158 66 8160
rect 0 8142 66 8158
rect 1632 8158 1648 8160
rect 1682 8190 1698 8192
rect 3264 8192 3330 8208
rect 3264 8190 3280 8192
rect 1682 8160 3280 8190
rect 1682 8158 1698 8160
rect 1632 8142 1698 8158
rect 3264 8158 3280 8160
rect 3314 8190 3330 8192
rect 4896 8192 4962 8208
rect 4896 8190 4912 8192
rect 3314 8160 4912 8190
rect 3314 8158 3330 8160
rect 3264 8142 3330 8158
rect 4896 8158 4912 8160
rect 4946 8190 4962 8192
rect 6528 8192 6594 8208
rect 6528 8190 6544 8192
rect 4946 8160 6544 8190
rect 4946 8158 4962 8160
rect 4896 8142 4962 8158
rect 6528 8158 6544 8160
rect 6578 8190 6594 8192
rect 8160 8192 8226 8208
rect 8160 8190 8176 8192
rect 6578 8160 8176 8190
rect 6578 8158 6594 8160
rect 6528 8142 6594 8158
rect 8160 8158 8176 8160
rect 8210 8190 8226 8192
rect 9792 8192 9858 8208
rect 9792 8190 9808 8192
rect 8210 8160 9808 8190
rect 8210 8158 8226 8160
rect 8160 8142 8226 8158
rect 9792 8158 9808 8160
rect 9842 8158 9858 8192
rect 9792 8142 9858 8158
rect 0 7988 66 8004
rect 0 7954 16 7988
rect 50 7986 66 7988
rect 1632 7988 1698 8004
rect 1632 7986 1648 7988
rect 50 7956 1648 7986
rect 50 7954 66 7956
rect 0 7938 66 7954
rect 1632 7954 1648 7956
rect 1682 7986 1698 7988
rect 3264 7988 3330 8004
rect 3264 7986 3280 7988
rect 1682 7956 3280 7986
rect 1682 7954 1698 7956
rect 1632 7938 1698 7954
rect 3264 7954 3280 7956
rect 3314 7986 3330 7988
rect 4896 7988 4962 8004
rect 4896 7986 4912 7988
rect 3314 7956 4912 7986
rect 3314 7954 3330 7956
rect 3264 7938 3330 7954
rect 4896 7954 4912 7956
rect 4946 7986 4962 7988
rect 6528 7988 6594 8004
rect 6528 7986 6544 7988
rect 4946 7956 6544 7986
rect 4946 7954 4962 7956
rect 4896 7938 4962 7954
rect 6528 7954 6544 7956
rect 6578 7986 6594 7988
rect 8160 7988 8226 8004
rect 8160 7986 8176 7988
rect 6578 7956 8176 7986
rect 6578 7954 6594 7956
rect 6528 7938 6594 7954
rect 8160 7954 8176 7956
rect 8210 7986 8226 7988
rect 9792 7988 9858 8004
rect 9792 7986 9808 7988
rect 8210 7956 9808 7986
rect 8210 7954 8226 7956
rect 8160 7938 8226 7954
rect 9792 7954 9808 7956
rect 9842 7954 9858 7988
rect 9792 7938 9858 7954
rect 0 7680 66 7696
rect 0 7646 16 7680
rect 50 7678 66 7680
rect 1632 7680 1698 7696
rect 1632 7678 1648 7680
rect 50 7648 1648 7678
rect 50 7646 66 7648
rect 0 7630 66 7646
rect 1632 7646 1648 7648
rect 1682 7678 1698 7680
rect 3264 7680 3330 7696
rect 3264 7678 3280 7680
rect 1682 7648 3280 7678
rect 1682 7646 1698 7648
rect 1632 7630 1698 7646
rect 3264 7646 3280 7648
rect 3314 7678 3330 7680
rect 4896 7680 4962 7696
rect 4896 7678 4912 7680
rect 3314 7648 4912 7678
rect 3314 7646 3330 7648
rect 3264 7630 3330 7646
rect 4896 7646 4912 7648
rect 4946 7678 4962 7680
rect 6528 7680 6594 7696
rect 6528 7678 6544 7680
rect 4946 7648 6544 7678
rect 4946 7646 4962 7648
rect 4896 7630 4962 7646
rect 6528 7646 6544 7648
rect 6578 7678 6594 7680
rect 8160 7680 8226 7696
rect 8160 7678 8176 7680
rect 6578 7648 8176 7678
rect 6578 7646 6594 7648
rect 6528 7630 6594 7646
rect 8160 7646 8176 7648
rect 8210 7678 8226 7680
rect 9792 7680 9858 7696
rect 9792 7678 9808 7680
rect 8210 7648 9808 7678
rect 8210 7646 8226 7648
rect 8160 7630 8226 7646
rect 9792 7646 9808 7648
rect 9842 7646 9858 7680
rect 9792 7630 9858 7646
rect 0 7476 66 7492
rect 0 7442 16 7476
rect 50 7474 66 7476
rect 1632 7476 1698 7492
rect 1632 7474 1648 7476
rect 50 7444 1648 7474
rect 50 7442 66 7444
rect 0 7426 66 7442
rect 1632 7442 1648 7444
rect 1682 7474 1698 7476
rect 3264 7476 3330 7492
rect 3264 7474 3280 7476
rect 1682 7444 3280 7474
rect 1682 7442 1698 7444
rect 1632 7426 1698 7442
rect 3264 7442 3280 7444
rect 3314 7474 3330 7476
rect 4896 7476 4962 7492
rect 4896 7474 4912 7476
rect 3314 7444 4912 7474
rect 3314 7442 3330 7444
rect 3264 7426 3330 7442
rect 4896 7442 4912 7444
rect 4946 7474 4962 7476
rect 6528 7476 6594 7492
rect 6528 7474 6544 7476
rect 4946 7444 6544 7474
rect 4946 7442 4962 7444
rect 4896 7426 4962 7442
rect 6528 7442 6544 7444
rect 6578 7474 6594 7476
rect 8160 7476 8226 7492
rect 8160 7474 8176 7476
rect 6578 7444 8176 7474
rect 6578 7442 6594 7444
rect 6528 7426 6594 7442
rect 8160 7442 8176 7444
rect 8210 7474 8226 7476
rect 9792 7476 9858 7492
rect 9792 7474 9808 7476
rect 8210 7444 9808 7474
rect 8210 7442 8226 7444
rect 8160 7426 8226 7442
rect 9792 7442 9808 7444
rect 9842 7442 9858 7476
rect 9792 7426 9858 7442
rect 0 7272 66 7288
rect 0 7238 16 7272
rect 50 7270 66 7272
rect 1632 7272 1698 7288
rect 1632 7270 1648 7272
rect 50 7240 1648 7270
rect 50 7238 66 7240
rect 0 7222 66 7238
rect 1632 7238 1648 7240
rect 1682 7270 1698 7272
rect 3264 7272 3330 7288
rect 3264 7270 3280 7272
rect 1682 7240 3280 7270
rect 1682 7238 1698 7240
rect 1632 7222 1698 7238
rect 3264 7238 3280 7240
rect 3314 7270 3330 7272
rect 4896 7272 4962 7288
rect 4896 7270 4912 7272
rect 3314 7240 4912 7270
rect 3314 7238 3330 7240
rect 3264 7222 3330 7238
rect 4896 7238 4912 7240
rect 4946 7270 4962 7272
rect 6528 7272 6594 7288
rect 6528 7270 6544 7272
rect 4946 7240 6544 7270
rect 4946 7238 4962 7240
rect 4896 7222 4962 7238
rect 6528 7238 6544 7240
rect 6578 7270 6594 7272
rect 8160 7272 8226 7288
rect 8160 7270 8176 7272
rect 6578 7240 8176 7270
rect 6578 7238 6594 7240
rect 6528 7222 6594 7238
rect 8160 7238 8176 7240
rect 8210 7270 8226 7272
rect 9792 7272 9858 7288
rect 9792 7270 9808 7272
rect 8210 7240 9808 7270
rect 8210 7238 8226 7240
rect 8160 7222 8226 7238
rect 9792 7238 9808 7240
rect 9842 7238 9858 7272
rect 9792 7222 9858 7238
rect 0 7068 66 7084
rect 0 7034 16 7068
rect 50 7066 66 7068
rect 1632 7068 1698 7084
rect 1632 7066 1648 7068
rect 50 7036 1648 7066
rect 50 7034 66 7036
rect 0 7018 66 7034
rect 1632 7034 1648 7036
rect 1682 7066 1698 7068
rect 3264 7068 3330 7084
rect 3264 7066 3280 7068
rect 1682 7036 3280 7066
rect 1682 7034 1698 7036
rect 1632 7018 1698 7034
rect 3264 7034 3280 7036
rect 3314 7066 3330 7068
rect 4896 7068 4962 7084
rect 4896 7066 4912 7068
rect 3314 7036 4912 7066
rect 3314 7034 3330 7036
rect 3264 7018 3330 7034
rect 4896 7034 4912 7036
rect 4946 7066 4962 7068
rect 6528 7068 6594 7084
rect 6528 7066 6544 7068
rect 4946 7036 6544 7066
rect 4946 7034 4962 7036
rect 4896 7018 4962 7034
rect 6528 7034 6544 7036
rect 6578 7066 6594 7068
rect 8160 7068 8226 7084
rect 8160 7066 8176 7068
rect 6578 7036 8176 7066
rect 6578 7034 6594 7036
rect 6528 7018 6594 7034
rect 8160 7034 8176 7036
rect 8210 7066 8226 7068
rect 9792 7068 9858 7084
rect 9792 7066 9808 7068
rect 8210 7036 9808 7066
rect 8210 7034 8226 7036
rect 8160 7018 8226 7034
rect 9792 7034 9808 7036
rect 9842 7034 9858 7068
rect 9792 7018 9858 7034
rect 0 6864 66 6880
rect 0 6830 16 6864
rect 50 6862 66 6864
rect 1632 6864 1698 6880
rect 1632 6862 1648 6864
rect 50 6832 1648 6862
rect 50 6830 66 6832
rect 0 6814 66 6830
rect 1632 6830 1648 6832
rect 1682 6862 1698 6864
rect 3264 6864 3330 6880
rect 3264 6862 3280 6864
rect 1682 6832 3280 6862
rect 1682 6830 1698 6832
rect 1632 6814 1698 6830
rect 3264 6830 3280 6832
rect 3314 6862 3330 6864
rect 4896 6864 4962 6880
rect 4896 6862 4912 6864
rect 3314 6832 4912 6862
rect 3314 6830 3330 6832
rect 3264 6814 3330 6830
rect 4896 6830 4912 6832
rect 4946 6862 4962 6864
rect 6528 6864 6594 6880
rect 6528 6862 6544 6864
rect 4946 6832 6544 6862
rect 4946 6830 4962 6832
rect 4896 6814 4962 6830
rect 6528 6830 6544 6832
rect 6578 6862 6594 6864
rect 8160 6864 8226 6880
rect 8160 6862 8176 6864
rect 6578 6832 8176 6862
rect 6578 6830 6594 6832
rect 6528 6814 6594 6830
rect 8160 6830 8176 6832
rect 8210 6862 8226 6864
rect 9792 6864 9858 6880
rect 9792 6862 9808 6864
rect 8210 6832 9808 6862
rect 8210 6830 8226 6832
rect 8160 6814 8226 6830
rect 9792 6830 9808 6832
rect 9842 6830 9858 6864
rect 9792 6814 9858 6830
rect 0 6660 66 6676
rect 0 6626 16 6660
rect 50 6658 66 6660
rect 1632 6660 1698 6676
rect 1632 6658 1648 6660
rect 50 6628 1648 6658
rect 50 6626 66 6628
rect 0 6610 66 6626
rect 1632 6626 1648 6628
rect 1682 6658 1698 6660
rect 3264 6660 3330 6676
rect 3264 6658 3280 6660
rect 1682 6628 3280 6658
rect 1682 6626 1698 6628
rect 1632 6610 1698 6626
rect 3264 6626 3280 6628
rect 3314 6658 3330 6660
rect 4896 6660 4962 6676
rect 4896 6658 4912 6660
rect 3314 6628 4912 6658
rect 3314 6626 3330 6628
rect 3264 6610 3330 6626
rect 4896 6626 4912 6628
rect 4946 6658 4962 6660
rect 6528 6660 6594 6676
rect 6528 6658 6544 6660
rect 4946 6628 6544 6658
rect 4946 6626 4962 6628
rect 4896 6610 4962 6626
rect 6528 6626 6544 6628
rect 6578 6658 6594 6660
rect 8160 6660 8226 6676
rect 8160 6658 8176 6660
rect 6578 6628 8176 6658
rect 6578 6626 6594 6628
rect 6528 6610 6594 6626
rect 8160 6626 8176 6628
rect 8210 6658 8226 6660
rect 9792 6660 9858 6676
rect 9792 6658 9808 6660
rect 8210 6628 9808 6658
rect 8210 6626 8226 6628
rect 8160 6610 8226 6626
rect 9792 6626 9808 6628
rect 9842 6626 9858 6660
rect 9792 6610 9858 6626
rect 0 6456 66 6472
rect 0 6422 16 6456
rect 50 6454 66 6456
rect 1632 6456 1698 6472
rect 1632 6454 1648 6456
rect 50 6424 1648 6454
rect 50 6422 66 6424
rect 0 6406 66 6422
rect 1632 6422 1648 6424
rect 1682 6454 1698 6456
rect 3264 6456 3330 6472
rect 3264 6454 3280 6456
rect 1682 6424 3280 6454
rect 1682 6422 1698 6424
rect 1632 6406 1698 6422
rect 3264 6422 3280 6424
rect 3314 6454 3330 6456
rect 4896 6456 4962 6472
rect 4896 6454 4912 6456
rect 3314 6424 4912 6454
rect 3314 6422 3330 6424
rect 3264 6406 3330 6422
rect 4896 6422 4912 6424
rect 4946 6454 4962 6456
rect 6528 6456 6594 6472
rect 6528 6454 6544 6456
rect 4946 6424 6544 6454
rect 4946 6422 4962 6424
rect 4896 6406 4962 6422
rect 6528 6422 6544 6424
rect 6578 6454 6594 6456
rect 8160 6456 8226 6472
rect 8160 6454 8176 6456
rect 6578 6424 8176 6454
rect 6578 6422 6594 6424
rect 6528 6406 6594 6422
rect 8160 6422 8176 6424
rect 8210 6454 8226 6456
rect 9792 6456 9858 6472
rect 9792 6454 9808 6456
rect 8210 6424 9808 6454
rect 8210 6422 8226 6424
rect 8160 6406 8226 6422
rect 9792 6422 9808 6424
rect 9842 6422 9858 6456
rect 9792 6406 9858 6422
rect 0 6252 66 6268
rect 0 6218 16 6252
rect 50 6250 66 6252
rect 1632 6252 1698 6268
rect 1632 6250 1648 6252
rect 50 6220 1648 6250
rect 50 6218 66 6220
rect 0 6202 66 6218
rect 1632 6218 1648 6220
rect 1682 6250 1698 6252
rect 3264 6252 3330 6268
rect 3264 6250 3280 6252
rect 1682 6220 3280 6250
rect 1682 6218 1698 6220
rect 1632 6202 1698 6218
rect 3264 6218 3280 6220
rect 3314 6250 3330 6252
rect 4896 6252 4962 6268
rect 4896 6250 4912 6252
rect 3314 6220 4912 6250
rect 3314 6218 3330 6220
rect 3264 6202 3330 6218
rect 4896 6218 4912 6220
rect 4946 6250 4962 6252
rect 6528 6252 6594 6268
rect 6528 6250 6544 6252
rect 4946 6220 6544 6250
rect 4946 6218 4962 6220
rect 4896 6202 4962 6218
rect 6528 6218 6544 6220
rect 6578 6250 6594 6252
rect 8160 6252 8226 6268
rect 8160 6250 8176 6252
rect 6578 6220 8176 6250
rect 6578 6218 6594 6220
rect 6528 6202 6594 6218
rect 8160 6218 8176 6220
rect 8210 6250 8226 6252
rect 9792 6252 9858 6268
rect 9792 6250 9808 6252
rect 8210 6220 9808 6250
rect 8210 6218 8226 6220
rect 8160 6202 8226 6218
rect 9792 6218 9808 6220
rect 9842 6218 9858 6252
rect 9792 6202 9858 6218
rect 0 5944 66 5960
rect 0 5910 16 5944
rect 50 5942 66 5944
rect 1632 5944 1698 5960
rect 1632 5942 1648 5944
rect 50 5912 1648 5942
rect 50 5910 66 5912
rect 0 5894 66 5910
rect 1632 5910 1648 5912
rect 1682 5942 1698 5944
rect 3264 5944 3330 5960
rect 3264 5942 3280 5944
rect 1682 5912 3280 5942
rect 1682 5910 1698 5912
rect 1632 5894 1698 5910
rect 3264 5910 3280 5912
rect 3314 5942 3330 5944
rect 4896 5944 4962 5960
rect 4896 5942 4912 5944
rect 3314 5912 4912 5942
rect 3314 5910 3330 5912
rect 3264 5894 3330 5910
rect 4896 5910 4912 5912
rect 4946 5942 4962 5944
rect 6528 5944 6594 5960
rect 6528 5942 6544 5944
rect 4946 5912 6544 5942
rect 4946 5910 4962 5912
rect 4896 5894 4962 5910
rect 6528 5910 6544 5912
rect 6578 5942 6594 5944
rect 8160 5944 8226 5960
rect 8160 5942 8176 5944
rect 6578 5912 8176 5942
rect 6578 5910 6594 5912
rect 6528 5894 6594 5910
rect 8160 5910 8176 5912
rect 8210 5942 8226 5944
rect 9792 5944 9858 5960
rect 9792 5942 9808 5944
rect 8210 5912 9808 5942
rect 8210 5910 8226 5912
rect 8160 5894 8226 5910
rect 9792 5910 9808 5912
rect 9842 5910 9858 5944
rect 9792 5894 9858 5910
rect 0 5740 66 5756
rect 0 5706 16 5740
rect 50 5738 66 5740
rect 1632 5740 1698 5756
rect 1632 5738 1648 5740
rect 50 5708 1648 5738
rect 50 5706 66 5708
rect 0 5690 66 5706
rect 1632 5706 1648 5708
rect 1682 5738 1698 5740
rect 3264 5740 3330 5756
rect 3264 5738 3280 5740
rect 1682 5708 3280 5738
rect 1682 5706 1698 5708
rect 1632 5690 1698 5706
rect 3264 5706 3280 5708
rect 3314 5738 3330 5740
rect 4896 5740 4962 5756
rect 4896 5738 4912 5740
rect 3314 5708 4912 5738
rect 3314 5706 3330 5708
rect 3264 5690 3330 5706
rect 4896 5706 4912 5708
rect 4946 5738 4962 5740
rect 6528 5740 6594 5756
rect 6528 5738 6544 5740
rect 4946 5708 6544 5738
rect 4946 5706 4962 5708
rect 4896 5690 4962 5706
rect 6528 5706 6544 5708
rect 6578 5738 6594 5740
rect 8160 5740 8226 5756
rect 8160 5738 8176 5740
rect 6578 5708 8176 5738
rect 6578 5706 6594 5708
rect 6528 5690 6594 5706
rect 8160 5706 8176 5708
rect 8210 5738 8226 5740
rect 9792 5740 9858 5756
rect 9792 5738 9808 5740
rect 8210 5708 9808 5738
rect 8210 5706 8226 5708
rect 8160 5690 8226 5706
rect 9792 5706 9808 5708
rect 9842 5706 9858 5740
rect 9792 5690 9858 5706
rect 0 5536 66 5552
rect 0 5502 16 5536
rect 50 5534 66 5536
rect 1632 5536 1698 5552
rect 1632 5534 1648 5536
rect 50 5504 1648 5534
rect 50 5502 66 5504
rect 0 5486 66 5502
rect 1632 5502 1648 5504
rect 1682 5534 1698 5536
rect 3264 5536 3330 5552
rect 3264 5534 3280 5536
rect 1682 5504 3280 5534
rect 1682 5502 1698 5504
rect 1632 5486 1698 5502
rect 3264 5502 3280 5504
rect 3314 5534 3330 5536
rect 4896 5536 4962 5552
rect 4896 5534 4912 5536
rect 3314 5504 4912 5534
rect 3314 5502 3330 5504
rect 3264 5486 3330 5502
rect 4896 5502 4912 5504
rect 4946 5534 4962 5536
rect 6528 5536 6594 5552
rect 6528 5534 6544 5536
rect 4946 5504 6544 5534
rect 4946 5502 4962 5504
rect 4896 5486 4962 5502
rect 6528 5502 6544 5504
rect 6578 5534 6594 5536
rect 8160 5536 8226 5552
rect 8160 5534 8176 5536
rect 6578 5504 8176 5534
rect 6578 5502 6594 5504
rect 6528 5486 6594 5502
rect 8160 5502 8176 5504
rect 8210 5534 8226 5536
rect 9792 5536 9858 5552
rect 9792 5534 9808 5536
rect 8210 5504 9808 5534
rect 8210 5502 8226 5504
rect 8160 5486 8226 5502
rect 9792 5502 9808 5504
rect 9842 5502 9858 5536
rect 9792 5486 9858 5502
rect 0 5332 66 5348
rect 0 5298 16 5332
rect 50 5330 66 5332
rect 1632 5332 1698 5348
rect 1632 5330 1648 5332
rect 50 5300 1648 5330
rect 50 5298 66 5300
rect 0 5282 66 5298
rect 1632 5298 1648 5300
rect 1682 5330 1698 5332
rect 3264 5332 3330 5348
rect 3264 5330 3280 5332
rect 1682 5300 3280 5330
rect 1682 5298 1698 5300
rect 1632 5282 1698 5298
rect 3264 5298 3280 5300
rect 3314 5330 3330 5332
rect 4896 5332 4962 5348
rect 4896 5330 4912 5332
rect 3314 5300 4912 5330
rect 3314 5298 3330 5300
rect 3264 5282 3330 5298
rect 4896 5298 4912 5300
rect 4946 5330 4962 5332
rect 6528 5332 6594 5348
rect 6528 5330 6544 5332
rect 4946 5300 6544 5330
rect 4946 5298 4962 5300
rect 4896 5282 4962 5298
rect 6528 5298 6544 5300
rect 6578 5330 6594 5332
rect 8160 5332 8226 5348
rect 8160 5330 8176 5332
rect 6578 5300 8176 5330
rect 6578 5298 6594 5300
rect 6528 5282 6594 5298
rect 8160 5298 8176 5300
rect 8210 5330 8226 5332
rect 9792 5332 9858 5348
rect 9792 5330 9808 5332
rect 8210 5300 9808 5330
rect 8210 5298 8226 5300
rect 8160 5282 8226 5298
rect 9792 5298 9808 5300
rect 9842 5298 9858 5332
rect 9792 5282 9858 5298
rect 0 5128 66 5144
rect 0 5094 16 5128
rect 50 5126 66 5128
rect 1632 5128 1698 5144
rect 1632 5126 1648 5128
rect 50 5096 1648 5126
rect 50 5094 66 5096
rect 0 5078 66 5094
rect 1632 5094 1648 5096
rect 1682 5126 1698 5128
rect 3264 5128 3330 5144
rect 3264 5126 3280 5128
rect 1682 5096 3280 5126
rect 1682 5094 1698 5096
rect 1632 5078 1698 5094
rect 3264 5094 3280 5096
rect 3314 5126 3330 5128
rect 4896 5128 4962 5144
rect 4896 5126 4912 5128
rect 3314 5096 4912 5126
rect 3314 5094 3330 5096
rect 3264 5078 3330 5094
rect 4896 5094 4912 5096
rect 4946 5126 4962 5128
rect 6528 5128 6594 5144
rect 6528 5126 6544 5128
rect 4946 5096 6544 5126
rect 4946 5094 4962 5096
rect 4896 5078 4962 5094
rect 6528 5094 6544 5096
rect 6578 5126 6594 5128
rect 8160 5128 8226 5144
rect 8160 5126 8176 5128
rect 6578 5096 8176 5126
rect 6578 5094 6594 5096
rect 6528 5078 6594 5094
rect 8160 5094 8176 5096
rect 8210 5126 8226 5128
rect 9792 5128 9858 5144
rect 9792 5126 9808 5128
rect 8210 5096 9808 5126
rect 8210 5094 8226 5096
rect 8160 5078 8226 5094
rect 9792 5094 9808 5096
rect 9842 5094 9858 5128
rect 9792 5078 9858 5094
rect 0 4924 66 4940
rect 0 4890 16 4924
rect 50 4922 66 4924
rect 1632 4924 1698 4940
rect 1632 4922 1648 4924
rect 50 4892 1648 4922
rect 50 4890 66 4892
rect 0 4874 66 4890
rect 1632 4890 1648 4892
rect 1682 4922 1698 4924
rect 3264 4924 3330 4940
rect 3264 4922 3280 4924
rect 1682 4892 3280 4922
rect 1682 4890 1698 4892
rect 1632 4874 1698 4890
rect 3264 4890 3280 4892
rect 3314 4922 3330 4924
rect 4896 4924 4962 4940
rect 4896 4922 4912 4924
rect 3314 4892 4912 4922
rect 3314 4890 3330 4892
rect 3264 4874 3330 4890
rect 4896 4890 4912 4892
rect 4946 4922 4962 4924
rect 6528 4924 6594 4940
rect 6528 4922 6544 4924
rect 4946 4892 6544 4922
rect 4946 4890 4962 4892
rect 4896 4874 4962 4890
rect 6528 4890 6544 4892
rect 6578 4922 6594 4924
rect 8160 4924 8226 4940
rect 8160 4922 8176 4924
rect 6578 4892 8176 4922
rect 6578 4890 6594 4892
rect 6528 4874 6594 4890
rect 8160 4890 8176 4892
rect 8210 4922 8226 4924
rect 9792 4924 9858 4940
rect 9792 4922 9808 4924
rect 8210 4892 9808 4922
rect 8210 4890 8226 4892
rect 8160 4874 8226 4890
rect 9792 4890 9808 4892
rect 9842 4890 9858 4924
rect 9792 4874 9858 4890
rect 0 4720 66 4736
rect 0 4686 16 4720
rect 50 4718 66 4720
rect 1632 4720 1698 4736
rect 1632 4718 1648 4720
rect 50 4688 1648 4718
rect 50 4686 66 4688
rect 0 4670 66 4686
rect 1632 4686 1648 4688
rect 1682 4718 1698 4720
rect 3264 4720 3330 4736
rect 3264 4718 3280 4720
rect 1682 4688 3280 4718
rect 1682 4686 1698 4688
rect 1632 4670 1698 4686
rect 3264 4686 3280 4688
rect 3314 4718 3330 4720
rect 4896 4720 4962 4736
rect 4896 4718 4912 4720
rect 3314 4688 4912 4718
rect 3314 4686 3330 4688
rect 3264 4670 3330 4686
rect 4896 4686 4912 4688
rect 4946 4718 4962 4720
rect 6528 4720 6594 4736
rect 6528 4718 6544 4720
rect 4946 4688 6544 4718
rect 4946 4686 4962 4688
rect 4896 4670 4962 4686
rect 6528 4686 6544 4688
rect 6578 4718 6594 4720
rect 8160 4720 8226 4736
rect 8160 4718 8176 4720
rect 6578 4688 8176 4718
rect 6578 4686 6594 4688
rect 6528 4670 6594 4686
rect 8160 4686 8176 4688
rect 8210 4718 8226 4720
rect 9792 4720 9858 4736
rect 9792 4718 9808 4720
rect 8210 4688 9808 4718
rect 8210 4686 8226 4688
rect 8160 4670 8226 4686
rect 9792 4686 9808 4688
rect 9842 4686 9858 4720
rect 9792 4670 9858 4686
rect 0 4516 66 4532
rect 0 4482 16 4516
rect 50 4514 66 4516
rect 1632 4516 1698 4532
rect 1632 4514 1648 4516
rect 50 4484 1648 4514
rect 50 4482 66 4484
rect 0 4466 66 4482
rect 1632 4482 1648 4484
rect 1682 4514 1698 4516
rect 3264 4516 3330 4532
rect 3264 4514 3280 4516
rect 1682 4484 3280 4514
rect 1682 4482 1698 4484
rect 1632 4466 1698 4482
rect 3264 4482 3280 4484
rect 3314 4514 3330 4516
rect 4896 4516 4962 4532
rect 4896 4514 4912 4516
rect 3314 4484 4912 4514
rect 3314 4482 3330 4484
rect 3264 4466 3330 4482
rect 4896 4482 4912 4484
rect 4946 4514 4962 4516
rect 6528 4516 6594 4532
rect 6528 4514 6544 4516
rect 4946 4484 6544 4514
rect 4946 4482 4962 4484
rect 4896 4466 4962 4482
rect 6528 4482 6544 4484
rect 6578 4514 6594 4516
rect 8160 4516 8226 4532
rect 8160 4514 8176 4516
rect 6578 4484 8176 4514
rect 6578 4482 6594 4484
rect 6528 4466 6594 4482
rect 8160 4482 8176 4484
rect 8210 4514 8226 4516
rect 9792 4516 9858 4532
rect 9792 4514 9808 4516
rect 8210 4484 9808 4514
rect 8210 4482 8226 4484
rect 8160 4466 8226 4482
rect 9792 4482 9808 4484
rect 9842 4482 9858 4516
rect 9792 4466 9858 4482
rect 0 4208 66 4224
rect 0 4174 16 4208
rect 50 4206 66 4208
rect 1632 4208 1698 4224
rect 1632 4206 1648 4208
rect 50 4176 1648 4206
rect 50 4174 66 4176
rect 0 4158 66 4174
rect 1632 4174 1648 4176
rect 1682 4206 1698 4208
rect 3264 4208 3330 4224
rect 3264 4206 3280 4208
rect 1682 4176 3280 4206
rect 1682 4174 1698 4176
rect 1632 4158 1698 4174
rect 3264 4174 3280 4176
rect 3314 4206 3330 4208
rect 4896 4208 4962 4224
rect 4896 4206 4912 4208
rect 3314 4176 4912 4206
rect 3314 4174 3330 4176
rect 3264 4158 3330 4174
rect 4896 4174 4912 4176
rect 4946 4206 4962 4208
rect 6528 4208 6594 4224
rect 6528 4206 6544 4208
rect 4946 4176 6544 4206
rect 4946 4174 4962 4176
rect 4896 4158 4962 4174
rect 6528 4174 6544 4176
rect 6578 4206 6594 4208
rect 8160 4208 8226 4224
rect 8160 4206 8176 4208
rect 6578 4176 8176 4206
rect 6578 4174 6594 4176
rect 6528 4158 6594 4174
rect 8160 4174 8176 4176
rect 8210 4206 8226 4208
rect 9792 4208 9858 4224
rect 9792 4206 9808 4208
rect 8210 4176 9808 4206
rect 8210 4174 8226 4176
rect 8160 4158 8226 4174
rect 9792 4174 9808 4176
rect 9842 4174 9858 4208
rect 9792 4158 9858 4174
rect 0 4004 66 4020
rect 0 3970 16 4004
rect 50 4002 66 4004
rect 1632 4004 1698 4020
rect 1632 4002 1648 4004
rect 50 3972 1648 4002
rect 50 3970 66 3972
rect 0 3954 66 3970
rect 1632 3970 1648 3972
rect 1682 4002 1698 4004
rect 3264 4004 3330 4020
rect 3264 4002 3280 4004
rect 1682 3972 3280 4002
rect 1682 3970 1698 3972
rect 1632 3954 1698 3970
rect 3264 3970 3280 3972
rect 3314 4002 3330 4004
rect 4896 4004 4962 4020
rect 4896 4002 4912 4004
rect 3314 3972 4912 4002
rect 3314 3970 3330 3972
rect 3264 3954 3330 3970
rect 4896 3970 4912 3972
rect 4946 4002 4962 4004
rect 6528 4004 6594 4020
rect 6528 4002 6544 4004
rect 4946 3972 6544 4002
rect 4946 3970 4962 3972
rect 4896 3954 4962 3970
rect 6528 3970 6544 3972
rect 6578 4002 6594 4004
rect 8160 4004 8226 4020
rect 8160 4002 8176 4004
rect 6578 3972 8176 4002
rect 6578 3970 6594 3972
rect 6528 3954 6594 3970
rect 8160 3970 8176 3972
rect 8210 4002 8226 4004
rect 9792 4004 9858 4020
rect 9792 4002 9808 4004
rect 8210 3972 9808 4002
rect 8210 3970 8226 3972
rect 8160 3954 8226 3970
rect 9792 3970 9808 3972
rect 9842 3970 9858 4004
rect 9792 3954 9858 3970
rect 0 3800 66 3816
rect 0 3766 16 3800
rect 50 3798 66 3800
rect 1632 3800 1698 3816
rect 1632 3798 1648 3800
rect 50 3768 1648 3798
rect 50 3766 66 3768
rect 0 3750 66 3766
rect 1632 3766 1648 3768
rect 1682 3798 1698 3800
rect 3264 3800 3330 3816
rect 3264 3798 3280 3800
rect 1682 3768 3280 3798
rect 1682 3766 1698 3768
rect 1632 3750 1698 3766
rect 3264 3766 3280 3768
rect 3314 3798 3330 3800
rect 4896 3800 4962 3816
rect 4896 3798 4912 3800
rect 3314 3768 4912 3798
rect 3314 3766 3330 3768
rect 3264 3750 3330 3766
rect 4896 3766 4912 3768
rect 4946 3798 4962 3800
rect 6528 3800 6594 3816
rect 6528 3798 6544 3800
rect 4946 3768 6544 3798
rect 4946 3766 4962 3768
rect 4896 3750 4962 3766
rect 6528 3766 6544 3768
rect 6578 3798 6594 3800
rect 8160 3800 8226 3816
rect 8160 3798 8176 3800
rect 6578 3768 8176 3798
rect 6578 3766 6594 3768
rect 6528 3750 6594 3766
rect 8160 3766 8176 3768
rect 8210 3798 8226 3800
rect 9792 3800 9858 3816
rect 9792 3798 9808 3800
rect 8210 3768 9808 3798
rect 8210 3766 8226 3768
rect 8160 3750 8226 3766
rect 9792 3766 9808 3768
rect 9842 3766 9858 3800
rect 9792 3750 9858 3766
rect 0 3596 66 3612
rect 0 3562 16 3596
rect 50 3594 66 3596
rect 1632 3596 1698 3612
rect 1632 3594 1648 3596
rect 50 3564 1648 3594
rect 50 3562 66 3564
rect 0 3546 66 3562
rect 1632 3562 1648 3564
rect 1682 3594 1698 3596
rect 3264 3596 3330 3612
rect 3264 3594 3280 3596
rect 1682 3564 3280 3594
rect 1682 3562 1698 3564
rect 1632 3546 1698 3562
rect 3264 3562 3280 3564
rect 3314 3594 3330 3596
rect 4896 3596 4962 3612
rect 4896 3594 4912 3596
rect 3314 3564 4912 3594
rect 3314 3562 3330 3564
rect 3264 3546 3330 3562
rect 4896 3562 4912 3564
rect 4946 3594 4962 3596
rect 6528 3596 6594 3612
rect 6528 3594 6544 3596
rect 4946 3564 6544 3594
rect 4946 3562 4962 3564
rect 4896 3546 4962 3562
rect 6528 3562 6544 3564
rect 6578 3594 6594 3596
rect 8160 3596 8226 3612
rect 8160 3594 8176 3596
rect 6578 3564 8176 3594
rect 6578 3562 6594 3564
rect 6528 3546 6594 3562
rect 8160 3562 8176 3564
rect 8210 3594 8226 3596
rect 9792 3596 9858 3612
rect 9792 3594 9808 3596
rect 8210 3564 9808 3594
rect 8210 3562 8226 3564
rect 8160 3546 8226 3562
rect 9792 3562 9808 3564
rect 9842 3562 9858 3596
rect 9792 3546 9858 3562
rect 0 3392 66 3408
rect 0 3358 16 3392
rect 50 3390 66 3392
rect 1632 3392 1698 3408
rect 1632 3390 1648 3392
rect 50 3360 1648 3390
rect 50 3358 66 3360
rect 0 3342 66 3358
rect 1632 3358 1648 3360
rect 1682 3390 1698 3392
rect 3264 3392 3330 3408
rect 3264 3390 3280 3392
rect 1682 3360 3280 3390
rect 1682 3358 1698 3360
rect 1632 3342 1698 3358
rect 3264 3358 3280 3360
rect 3314 3390 3330 3392
rect 4896 3392 4962 3408
rect 4896 3390 4912 3392
rect 3314 3360 4912 3390
rect 3314 3358 3330 3360
rect 3264 3342 3330 3358
rect 4896 3358 4912 3360
rect 4946 3390 4962 3392
rect 6528 3392 6594 3408
rect 6528 3390 6544 3392
rect 4946 3360 6544 3390
rect 4946 3358 4962 3360
rect 4896 3342 4962 3358
rect 6528 3358 6544 3360
rect 6578 3390 6594 3392
rect 8160 3392 8226 3408
rect 8160 3390 8176 3392
rect 6578 3360 8176 3390
rect 6578 3358 6594 3360
rect 6528 3342 6594 3358
rect 8160 3358 8176 3360
rect 8210 3390 8226 3392
rect 9792 3392 9858 3408
rect 9792 3390 9808 3392
rect 8210 3360 9808 3390
rect 8210 3358 8226 3360
rect 8160 3342 8226 3358
rect 9792 3358 9808 3360
rect 9842 3358 9858 3392
rect 9792 3342 9858 3358
rect 0 3188 66 3204
rect 0 3154 16 3188
rect 50 3186 66 3188
rect 1632 3188 1698 3204
rect 1632 3186 1648 3188
rect 50 3156 1648 3186
rect 50 3154 66 3156
rect 0 3138 66 3154
rect 1632 3154 1648 3156
rect 1682 3186 1698 3188
rect 3264 3188 3330 3204
rect 3264 3186 3280 3188
rect 1682 3156 3280 3186
rect 1682 3154 1698 3156
rect 1632 3138 1698 3154
rect 3264 3154 3280 3156
rect 3314 3186 3330 3188
rect 4896 3188 4962 3204
rect 4896 3186 4912 3188
rect 3314 3156 4912 3186
rect 3314 3154 3330 3156
rect 3264 3138 3330 3154
rect 4896 3154 4912 3156
rect 4946 3186 4962 3188
rect 6528 3188 6594 3204
rect 6528 3186 6544 3188
rect 4946 3156 6544 3186
rect 4946 3154 4962 3156
rect 4896 3138 4962 3154
rect 6528 3154 6544 3156
rect 6578 3186 6594 3188
rect 8160 3188 8226 3204
rect 8160 3186 8176 3188
rect 6578 3156 8176 3186
rect 6578 3154 6594 3156
rect 6528 3138 6594 3154
rect 8160 3154 8176 3156
rect 8210 3186 8226 3188
rect 9792 3188 9858 3204
rect 9792 3186 9808 3188
rect 8210 3156 9808 3186
rect 8210 3154 8226 3156
rect 8160 3138 8226 3154
rect 9792 3154 9808 3156
rect 9842 3154 9858 3188
rect 9792 3138 9858 3154
rect 0 2984 66 3000
rect 0 2950 16 2984
rect 50 2982 66 2984
rect 1632 2984 1698 3000
rect 1632 2982 1648 2984
rect 50 2952 1648 2982
rect 50 2950 66 2952
rect 0 2934 66 2950
rect 1632 2950 1648 2952
rect 1682 2982 1698 2984
rect 3264 2984 3330 3000
rect 3264 2982 3280 2984
rect 1682 2952 3280 2982
rect 1682 2950 1698 2952
rect 1632 2934 1698 2950
rect 3264 2950 3280 2952
rect 3314 2982 3330 2984
rect 4896 2984 4962 3000
rect 4896 2982 4912 2984
rect 3314 2952 4912 2982
rect 3314 2950 3330 2952
rect 3264 2934 3330 2950
rect 4896 2950 4912 2952
rect 4946 2982 4962 2984
rect 6528 2984 6594 3000
rect 6528 2982 6544 2984
rect 4946 2952 6544 2982
rect 4946 2950 4962 2952
rect 4896 2934 4962 2950
rect 6528 2950 6544 2952
rect 6578 2982 6594 2984
rect 8160 2984 8226 3000
rect 8160 2982 8176 2984
rect 6578 2952 8176 2982
rect 6578 2950 6594 2952
rect 6528 2934 6594 2950
rect 8160 2950 8176 2952
rect 8210 2982 8226 2984
rect 9792 2984 9858 3000
rect 9792 2982 9808 2984
rect 8210 2952 9808 2982
rect 8210 2950 8226 2952
rect 8160 2934 8226 2950
rect 9792 2950 9808 2952
rect 9842 2950 9858 2984
rect 9792 2934 9858 2950
rect 0 2780 66 2796
rect 0 2746 16 2780
rect 50 2778 66 2780
rect 1632 2780 1698 2796
rect 1632 2778 1648 2780
rect 50 2748 1648 2778
rect 50 2746 66 2748
rect 0 2730 66 2746
rect 1632 2746 1648 2748
rect 1682 2778 1698 2780
rect 3264 2780 3330 2796
rect 3264 2778 3280 2780
rect 1682 2748 3280 2778
rect 1682 2746 1698 2748
rect 1632 2730 1698 2746
rect 3264 2746 3280 2748
rect 3314 2778 3330 2780
rect 4896 2780 4962 2796
rect 4896 2778 4912 2780
rect 3314 2748 4912 2778
rect 3314 2746 3330 2748
rect 3264 2730 3330 2746
rect 4896 2746 4912 2748
rect 4946 2778 4962 2780
rect 6528 2780 6594 2796
rect 6528 2778 6544 2780
rect 4946 2748 6544 2778
rect 4946 2746 4962 2748
rect 4896 2730 4962 2746
rect 6528 2746 6544 2748
rect 6578 2778 6594 2780
rect 8160 2780 8226 2796
rect 8160 2778 8176 2780
rect 6578 2748 8176 2778
rect 6578 2746 6594 2748
rect 6528 2730 6594 2746
rect 8160 2746 8176 2748
rect 8210 2778 8226 2780
rect 9792 2780 9858 2796
rect 9792 2778 9808 2780
rect 8210 2748 9808 2778
rect 8210 2746 8226 2748
rect 8160 2730 8226 2746
rect 9792 2746 9808 2748
rect 9842 2746 9858 2780
rect 9792 2730 9858 2746
rect 0 2472 66 2488
rect 0 2438 16 2472
rect 50 2470 66 2472
rect 1632 2472 1698 2488
rect 1632 2470 1648 2472
rect 50 2440 1648 2470
rect 50 2438 66 2440
rect 0 2422 66 2438
rect 1632 2438 1648 2440
rect 1682 2470 1698 2472
rect 3264 2472 3330 2488
rect 3264 2470 3280 2472
rect 1682 2440 3280 2470
rect 1682 2438 1698 2440
rect 1632 2422 1698 2438
rect 3264 2438 3280 2440
rect 3314 2470 3330 2472
rect 4896 2472 4962 2488
rect 4896 2470 4912 2472
rect 3314 2440 4912 2470
rect 3314 2438 3330 2440
rect 3264 2422 3330 2438
rect 4896 2438 4912 2440
rect 4946 2470 4962 2472
rect 6528 2472 6594 2488
rect 6528 2470 6544 2472
rect 4946 2440 6544 2470
rect 4946 2438 4962 2440
rect 4896 2422 4962 2438
rect 6528 2438 6544 2440
rect 6578 2470 6594 2472
rect 8160 2472 8226 2488
rect 8160 2470 8176 2472
rect 6578 2440 8176 2470
rect 6578 2438 6594 2440
rect 6528 2422 6594 2438
rect 8160 2438 8176 2440
rect 8210 2470 8226 2472
rect 9792 2472 9858 2488
rect 9792 2470 9808 2472
rect 8210 2440 9808 2470
rect 8210 2438 8226 2440
rect 8160 2422 8226 2438
rect 9792 2438 9808 2440
rect 9842 2438 9858 2472
rect 9792 2422 9858 2438
rect 0 2268 66 2284
rect 0 2234 16 2268
rect 50 2266 66 2268
rect 1632 2268 1698 2284
rect 1632 2266 1648 2268
rect 50 2236 1648 2266
rect 50 2234 66 2236
rect 0 2218 66 2234
rect 1632 2234 1648 2236
rect 1682 2266 1698 2268
rect 3264 2268 3330 2284
rect 3264 2266 3280 2268
rect 1682 2236 3280 2266
rect 1682 2234 1698 2236
rect 1632 2218 1698 2234
rect 3264 2234 3280 2236
rect 3314 2266 3330 2268
rect 4896 2268 4962 2284
rect 4896 2266 4912 2268
rect 3314 2236 4912 2266
rect 3314 2234 3330 2236
rect 3264 2218 3330 2234
rect 4896 2234 4912 2236
rect 4946 2266 4962 2268
rect 6528 2268 6594 2284
rect 6528 2266 6544 2268
rect 4946 2236 6544 2266
rect 4946 2234 4962 2236
rect 4896 2218 4962 2234
rect 6528 2234 6544 2236
rect 6578 2266 6594 2268
rect 8160 2268 8226 2284
rect 8160 2266 8176 2268
rect 6578 2236 8176 2266
rect 6578 2234 6594 2236
rect 6528 2218 6594 2234
rect 8160 2234 8176 2236
rect 8210 2266 8226 2268
rect 9792 2268 9858 2284
rect 9792 2266 9808 2268
rect 8210 2236 9808 2266
rect 8210 2234 8226 2236
rect 8160 2218 8226 2234
rect 9792 2234 9808 2236
rect 9842 2234 9858 2268
rect 9792 2218 9858 2234
rect 0 2064 66 2080
rect 0 2030 16 2064
rect 50 2062 66 2064
rect 1632 2064 1698 2080
rect 1632 2062 1648 2064
rect 50 2032 1648 2062
rect 50 2030 66 2032
rect 0 2014 66 2030
rect 1632 2030 1648 2032
rect 1682 2062 1698 2064
rect 3264 2064 3330 2080
rect 3264 2062 3280 2064
rect 1682 2032 3280 2062
rect 1682 2030 1698 2032
rect 1632 2014 1698 2030
rect 3264 2030 3280 2032
rect 3314 2062 3330 2064
rect 4896 2064 4962 2080
rect 4896 2062 4912 2064
rect 3314 2032 4912 2062
rect 3314 2030 3330 2032
rect 3264 2014 3330 2030
rect 4896 2030 4912 2032
rect 4946 2062 4962 2064
rect 6528 2064 6594 2080
rect 6528 2062 6544 2064
rect 4946 2032 6544 2062
rect 4946 2030 4962 2032
rect 4896 2014 4962 2030
rect 6528 2030 6544 2032
rect 6578 2062 6594 2064
rect 8160 2064 8226 2080
rect 8160 2062 8176 2064
rect 6578 2032 8176 2062
rect 6578 2030 6594 2032
rect 6528 2014 6594 2030
rect 8160 2030 8176 2032
rect 8210 2062 8226 2064
rect 9792 2064 9858 2080
rect 9792 2062 9808 2064
rect 8210 2032 9808 2062
rect 8210 2030 8226 2032
rect 8160 2014 8226 2030
rect 9792 2030 9808 2032
rect 9842 2030 9858 2064
rect 9792 2014 9858 2030
rect 0 1860 66 1876
rect 0 1826 16 1860
rect 50 1858 66 1860
rect 1632 1860 1698 1876
rect 1632 1858 1648 1860
rect 50 1828 1648 1858
rect 50 1826 66 1828
rect 0 1810 66 1826
rect 1632 1826 1648 1828
rect 1682 1858 1698 1860
rect 3264 1860 3330 1876
rect 3264 1858 3280 1860
rect 1682 1828 3280 1858
rect 1682 1826 1698 1828
rect 1632 1810 1698 1826
rect 3264 1826 3280 1828
rect 3314 1858 3330 1860
rect 4896 1860 4962 1876
rect 4896 1858 4912 1860
rect 3314 1828 4912 1858
rect 3314 1826 3330 1828
rect 3264 1810 3330 1826
rect 4896 1826 4912 1828
rect 4946 1858 4962 1860
rect 6528 1860 6594 1876
rect 6528 1858 6544 1860
rect 4946 1828 6544 1858
rect 4946 1826 4962 1828
rect 4896 1810 4962 1826
rect 6528 1826 6544 1828
rect 6578 1858 6594 1860
rect 8160 1860 8226 1876
rect 8160 1858 8176 1860
rect 6578 1828 8176 1858
rect 6578 1826 6594 1828
rect 6528 1810 6594 1826
rect 8160 1826 8176 1828
rect 8210 1858 8226 1860
rect 9792 1860 9858 1876
rect 9792 1858 9808 1860
rect 8210 1828 9808 1858
rect 8210 1826 8226 1828
rect 8160 1810 8226 1826
rect 9792 1826 9808 1828
rect 9842 1826 9858 1860
rect 9792 1810 9858 1826
rect 0 1656 66 1672
rect 0 1622 16 1656
rect 50 1654 66 1656
rect 1632 1656 1698 1672
rect 1632 1654 1648 1656
rect 50 1624 1648 1654
rect 50 1622 66 1624
rect 0 1606 66 1622
rect 1632 1622 1648 1624
rect 1682 1654 1698 1656
rect 3264 1656 3330 1672
rect 3264 1654 3280 1656
rect 1682 1624 3280 1654
rect 1682 1622 1698 1624
rect 1632 1606 1698 1622
rect 3264 1622 3280 1624
rect 3314 1654 3330 1656
rect 4896 1656 4962 1672
rect 4896 1654 4912 1656
rect 3314 1624 4912 1654
rect 3314 1622 3330 1624
rect 3264 1606 3330 1622
rect 4896 1622 4912 1624
rect 4946 1654 4962 1656
rect 6528 1656 6594 1672
rect 6528 1654 6544 1656
rect 4946 1624 6544 1654
rect 4946 1622 4962 1624
rect 4896 1606 4962 1622
rect 6528 1622 6544 1624
rect 6578 1654 6594 1656
rect 8160 1656 8226 1672
rect 8160 1654 8176 1656
rect 6578 1624 8176 1654
rect 6578 1622 6594 1624
rect 6528 1606 6594 1622
rect 8160 1622 8176 1624
rect 8210 1654 8226 1656
rect 9792 1656 9858 1672
rect 9792 1654 9808 1656
rect 8210 1624 9808 1654
rect 8210 1622 8226 1624
rect 8160 1606 8226 1622
rect 9792 1622 9808 1624
rect 9842 1622 9858 1656
rect 9792 1606 9858 1622
rect 0 1452 66 1468
rect 0 1418 16 1452
rect 50 1450 66 1452
rect 1632 1452 1698 1468
rect 1632 1450 1648 1452
rect 50 1420 1648 1450
rect 50 1418 66 1420
rect 0 1402 66 1418
rect 1632 1418 1648 1420
rect 1682 1450 1698 1452
rect 3264 1452 3330 1468
rect 3264 1450 3280 1452
rect 1682 1420 3280 1450
rect 1682 1418 1698 1420
rect 1632 1402 1698 1418
rect 3264 1418 3280 1420
rect 3314 1450 3330 1452
rect 4896 1452 4962 1468
rect 4896 1450 4912 1452
rect 3314 1420 4912 1450
rect 3314 1418 3330 1420
rect 3264 1402 3330 1418
rect 4896 1418 4912 1420
rect 4946 1450 4962 1452
rect 6528 1452 6594 1468
rect 6528 1450 6544 1452
rect 4946 1420 6544 1450
rect 4946 1418 4962 1420
rect 4896 1402 4962 1418
rect 6528 1418 6544 1420
rect 6578 1450 6594 1452
rect 8160 1452 8226 1468
rect 8160 1450 8176 1452
rect 6578 1420 8176 1450
rect 6578 1418 6594 1420
rect 6528 1402 6594 1418
rect 8160 1418 8176 1420
rect 8210 1450 8226 1452
rect 9792 1452 9858 1468
rect 9792 1450 9808 1452
rect 8210 1420 9808 1450
rect 8210 1418 8226 1420
rect 8160 1402 8226 1418
rect 9792 1418 9808 1420
rect 9842 1418 9858 1452
rect 9792 1402 9858 1418
rect 0 1248 66 1264
rect 0 1214 16 1248
rect 50 1246 66 1248
rect 1632 1248 1698 1264
rect 1632 1246 1648 1248
rect 50 1216 1648 1246
rect 50 1214 66 1216
rect 0 1198 66 1214
rect 1632 1214 1648 1216
rect 1682 1246 1698 1248
rect 3264 1248 3330 1264
rect 3264 1246 3280 1248
rect 1682 1216 3280 1246
rect 1682 1214 1698 1216
rect 1632 1198 1698 1214
rect 3264 1214 3280 1216
rect 3314 1246 3330 1248
rect 4896 1248 4962 1264
rect 4896 1246 4912 1248
rect 3314 1216 4912 1246
rect 3314 1214 3330 1216
rect 3264 1198 3330 1214
rect 4896 1214 4912 1216
rect 4946 1246 4962 1248
rect 6528 1248 6594 1264
rect 6528 1246 6544 1248
rect 4946 1216 6544 1246
rect 4946 1214 4962 1216
rect 4896 1198 4962 1214
rect 6528 1214 6544 1216
rect 6578 1246 6594 1248
rect 8160 1248 8226 1264
rect 8160 1246 8176 1248
rect 6578 1216 8176 1246
rect 6578 1214 6594 1216
rect 6528 1198 6594 1214
rect 8160 1214 8176 1216
rect 8210 1246 8226 1248
rect 9792 1248 9858 1264
rect 9792 1246 9808 1248
rect 8210 1216 9808 1246
rect 8210 1214 8226 1216
rect 8160 1198 8226 1214
rect 9792 1214 9808 1216
rect 9842 1214 9858 1248
rect 9792 1198 9858 1214
rect 0 1044 66 1060
rect 0 1010 16 1044
rect 50 1042 66 1044
rect 1632 1044 1698 1060
rect 1632 1042 1648 1044
rect 50 1012 1648 1042
rect 50 1010 66 1012
rect 0 994 66 1010
rect 1632 1010 1648 1012
rect 1682 1042 1698 1044
rect 3264 1044 3330 1060
rect 3264 1042 3280 1044
rect 1682 1012 3280 1042
rect 1682 1010 1698 1012
rect 1632 994 1698 1010
rect 3264 1010 3280 1012
rect 3314 1042 3330 1044
rect 4896 1044 4962 1060
rect 4896 1042 4912 1044
rect 3314 1012 4912 1042
rect 3314 1010 3330 1012
rect 3264 994 3330 1010
rect 4896 1010 4912 1012
rect 4946 1042 4962 1044
rect 6528 1044 6594 1060
rect 6528 1042 6544 1044
rect 4946 1012 6544 1042
rect 4946 1010 4962 1012
rect 4896 994 4962 1010
rect 6528 1010 6544 1012
rect 6578 1042 6594 1044
rect 8160 1044 8226 1060
rect 8160 1042 8176 1044
rect 6578 1012 8176 1042
rect 6578 1010 6594 1012
rect 6528 994 6594 1010
rect 8160 1010 8176 1012
rect 8210 1042 8226 1044
rect 9792 1044 9858 1060
rect 9792 1042 9808 1044
rect 8210 1012 9808 1042
rect 8210 1010 8226 1012
rect 8160 994 8226 1010
rect 9792 1010 9808 1012
rect 9842 1010 9858 1044
rect 9792 994 9858 1010
<< polycont >>
rect 16 10098 50 10132
rect 1648 10098 1682 10132
rect 3280 10098 3314 10132
rect 4912 10098 4946 10132
rect 6544 10098 6578 10132
rect 8176 10098 8210 10132
rect 9808 10098 9842 10132
rect 16 9894 50 9928
rect 1648 9894 1682 9928
rect 3280 9894 3314 9928
rect 4912 9894 4946 9928
rect 6544 9894 6578 9928
rect 8176 9894 8210 9928
rect 9808 9894 9842 9928
rect 16 9690 50 9724
rect 1648 9690 1682 9724
rect 3280 9690 3314 9724
rect 4912 9690 4946 9724
rect 6544 9690 6578 9724
rect 8176 9690 8210 9724
rect 9808 9690 9842 9724
rect 16 9382 50 9416
rect 1648 9382 1682 9416
rect 3280 9382 3314 9416
rect 4912 9382 4946 9416
rect 6544 9382 6578 9416
rect 8176 9382 8210 9416
rect 9808 9382 9842 9416
rect 16 9178 50 9212
rect 1648 9178 1682 9212
rect 3280 9178 3314 9212
rect 4912 9178 4946 9212
rect 6544 9178 6578 9212
rect 8176 9178 8210 9212
rect 9808 9178 9842 9212
rect 16 8974 50 9008
rect 1648 8974 1682 9008
rect 3280 8974 3314 9008
rect 4912 8974 4946 9008
rect 6544 8974 6578 9008
rect 8176 8974 8210 9008
rect 9808 8974 9842 9008
rect 16 8770 50 8804
rect 1648 8770 1682 8804
rect 3280 8770 3314 8804
rect 4912 8770 4946 8804
rect 6544 8770 6578 8804
rect 8176 8770 8210 8804
rect 9808 8770 9842 8804
rect 16 8566 50 8600
rect 1648 8566 1682 8600
rect 3280 8566 3314 8600
rect 4912 8566 4946 8600
rect 6544 8566 6578 8600
rect 8176 8566 8210 8600
rect 9808 8566 9842 8600
rect 16 8362 50 8396
rect 1648 8362 1682 8396
rect 3280 8362 3314 8396
rect 4912 8362 4946 8396
rect 6544 8362 6578 8396
rect 8176 8362 8210 8396
rect 9808 8362 9842 8396
rect 16 8158 50 8192
rect 1648 8158 1682 8192
rect 3280 8158 3314 8192
rect 4912 8158 4946 8192
rect 6544 8158 6578 8192
rect 8176 8158 8210 8192
rect 9808 8158 9842 8192
rect 16 7954 50 7988
rect 1648 7954 1682 7988
rect 3280 7954 3314 7988
rect 4912 7954 4946 7988
rect 6544 7954 6578 7988
rect 8176 7954 8210 7988
rect 9808 7954 9842 7988
rect 16 7646 50 7680
rect 1648 7646 1682 7680
rect 3280 7646 3314 7680
rect 4912 7646 4946 7680
rect 6544 7646 6578 7680
rect 8176 7646 8210 7680
rect 9808 7646 9842 7680
rect 16 7442 50 7476
rect 1648 7442 1682 7476
rect 3280 7442 3314 7476
rect 4912 7442 4946 7476
rect 6544 7442 6578 7476
rect 8176 7442 8210 7476
rect 9808 7442 9842 7476
rect 16 7238 50 7272
rect 1648 7238 1682 7272
rect 3280 7238 3314 7272
rect 4912 7238 4946 7272
rect 6544 7238 6578 7272
rect 8176 7238 8210 7272
rect 9808 7238 9842 7272
rect 16 7034 50 7068
rect 1648 7034 1682 7068
rect 3280 7034 3314 7068
rect 4912 7034 4946 7068
rect 6544 7034 6578 7068
rect 8176 7034 8210 7068
rect 9808 7034 9842 7068
rect 16 6830 50 6864
rect 1648 6830 1682 6864
rect 3280 6830 3314 6864
rect 4912 6830 4946 6864
rect 6544 6830 6578 6864
rect 8176 6830 8210 6864
rect 9808 6830 9842 6864
rect 16 6626 50 6660
rect 1648 6626 1682 6660
rect 3280 6626 3314 6660
rect 4912 6626 4946 6660
rect 6544 6626 6578 6660
rect 8176 6626 8210 6660
rect 9808 6626 9842 6660
rect 16 6422 50 6456
rect 1648 6422 1682 6456
rect 3280 6422 3314 6456
rect 4912 6422 4946 6456
rect 6544 6422 6578 6456
rect 8176 6422 8210 6456
rect 9808 6422 9842 6456
rect 16 6218 50 6252
rect 1648 6218 1682 6252
rect 3280 6218 3314 6252
rect 4912 6218 4946 6252
rect 6544 6218 6578 6252
rect 8176 6218 8210 6252
rect 9808 6218 9842 6252
rect 16 5910 50 5944
rect 1648 5910 1682 5944
rect 3280 5910 3314 5944
rect 4912 5910 4946 5944
rect 6544 5910 6578 5944
rect 8176 5910 8210 5944
rect 9808 5910 9842 5944
rect 16 5706 50 5740
rect 1648 5706 1682 5740
rect 3280 5706 3314 5740
rect 4912 5706 4946 5740
rect 6544 5706 6578 5740
rect 8176 5706 8210 5740
rect 9808 5706 9842 5740
rect 16 5502 50 5536
rect 1648 5502 1682 5536
rect 3280 5502 3314 5536
rect 4912 5502 4946 5536
rect 6544 5502 6578 5536
rect 8176 5502 8210 5536
rect 9808 5502 9842 5536
rect 16 5298 50 5332
rect 1648 5298 1682 5332
rect 3280 5298 3314 5332
rect 4912 5298 4946 5332
rect 6544 5298 6578 5332
rect 8176 5298 8210 5332
rect 9808 5298 9842 5332
rect 16 5094 50 5128
rect 1648 5094 1682 5128
rect 3280 5094 3314 5128
rect 4912 5094 4946 5128
rect 6544 5094 6578 5128
rect 8176 5094 8210 5128
rect 9808 5094 9842 5128
rect 16 4890 50 4924
rect 1648 4890 1682 4924
rect 3280 4890 3314 4924
rect 4912 4890 4946 4924
rect 6544 4890 6578 4924
rect 8176 4890 8210 4924
rect 9808 4890 9842 4924
rect 16 4686 50 4720
rect 1648 4686 1682 4720
rect 3280 4686 3314 4720
rect 4912 4686 4946 4720
rect 6544 4686 6578 4720
rect 8176 4686 8210 4720
rect 9808 4686 9842 4720
rect 16 4482 50 4516
rect 1648 4482 1682 4516
rect 3280 4482 3314 4516
rect 4912 4482 4946 4516
rect 6544 4482 6578 4516
rect 8176 4482 8210 4516
rect 9808 4482 9842 4516
rect 16 4174 50 4208
rect 1648 4174 1682 4208
rect 3280 4174 3314 4208
rect 4912 4174 4946 4208
rect 6544 4174 6578 4208
rect 8176 4174 8210 4208
rect 9808 4174 9842 4208
rect 16 3970 50 4004
rect 1648 3970 1682 4004
rect 3280 3970 3314 4004
rect 4912 3970 4946 4004
rect 6544 3970 6578 4004
rect 8176 3970 8210 4004
rect 9808 3970 9842 4004
rect 16 3766 50 3800
rect 1648 3766 1682 3800
rect 3280 3766 3314 3800
rect 4912 3766 4946 3800
rect 6544 3766 6578 3800
rect 8176 3766 8210 3800
rect 9808 3766 9842 3800
rect 16 3562 50 3596
rect 1648 3562 1682 3596
rect 3280 3562 3314 3596
rect 4912 3562 4946 3596
rect 6544 3562 6578 3596
rect 8176 3562 8210 3596
rect 9808 3562 9842 3596
rect 16 3358 50 3392
rect 1648 3358 1682 3392
rect 3280 3358 3314 3392
rect 4912 3358 4946 3392
rect 6544 3358 6578 3392
rect 8176 3358 8210 3392
rect 9808 3358 9842 3392
rect 16 3154 50 3188
rect 1648 3154 1682 3188
rect 3280 3154 3314 3188
rect 4912 3154 4946 3188
rect 6544 3154 6578 3188
rect 8176 3154 8210 3188
rect 9808 3154 9842 3188
rect 16 2950 50 2984
rect 1648 2950 1682 2984
rect 3280 2950 3314 2984
rect 4912 2950 4946 2984
rect 6544 2950 6578 2984
rect 8176 2950 8210 2984
rect 9808 2950 9842 2984
rect 16 2746 50 2780
rect 1648 2746 1682 2780
rect 3280 2746 3314 2780
rect 4912 2746 4946 2780
rect 6544 2746 6578 2780
rect 8176 2746 8210 2780
rect 9808 2746 9842 2780
rect 16 2438 50 2472
rect 1648 2438 1682 2472
rect 3280 2438 3314 2472
rect 4912 2438 4946 2472
rect 6544 2438 6578 2472
rect 8176 2438 8210 2472
rect 9808 2438 9842 2472
rect 16 2234 50 2268
rect 1648 2234 1682 2268
rect 3280 2234 3314 2268
rect 4912 2234 4946 2268
rect 6544 2234 6578 2268
rect 8176 2234 8210 2268
rect 9808 2234 9842 2268
rect 16 2030 50 2064
rect 1648 2030 1682 2064
rect 3280 2030 3314 2064
rect 4912 2030 4946 2064
rect 6544 2030 6578 2064
rect 8176 2030 8210 2064
rect 9808 2030 9842 2064
rect 16 1826 50 1860
rect 1648 1826 1682 1860
rect 3280 1826 3314 1860
rect 4912 1826 4946 1860
rect 6544 1826 6578 1860
rect 8176 1826 8210 1860
rect 9808 1826 9842 1860
rect 16 1622 50 1656
rect 1648 1622 1682 1656
rect 3280 1622 3314 1656
rect 4912 1622 4946 1656
rect 6544 1622 6578 1656
rect 8176 1622 8210 1656
rect 9808 1622 9842 1656
rect 16 1418 50 1452
rect 1648 1418 1682 1452
rect 3280 1418 3314 1452
rect 4912 1418 4946 1452
rect 6544 1418 6578 1452
rect 8176 1418 8210 1452
rect 9808 1418 9842 1452
rect 16 1214 50 1248
rect 1648 1214 1682 1248
rect 3280 1214 3314 1248
rect 4912 1214 4946 1248
rect 6544 1214 6578 1248
rect 8176 1214 8210 1248
rect 9808 1214 9842 1248
rect 16 1010 50 1044
rect 1648 1010 1682 1044
rect 3280 1010 3314 1044
rect 4912 1010 4946 1044
rect 6544 1010 6578 1044
rect 8176 1010 8210 1044
rect 9808 1010 9842 1044
<< locali >>
rect 16 10132 50 10148
rect 16 10082 50 10098
rect 1648 10132 1682 10148
rect 1648 10082 1682 10098
rect 3280 10132 3314 10148
rect 3280 10082 3314 10098
rect 4912 10132 4946 10148
rect 4912 10082 4946 10098
rect 6544 10132 6578 10148
rect 6544 10082 6578 10098
rect 8176 10132 8210 10148
rect 8176 10082 8210 10098
rect 9808 10132 9842 10148
rect 9808 10082 9842 10098
rect 16 9928 50 9944
rect 16 9878 50 9894
rect 1648 9928 1682 9944
rect 1648 9878 1682 9894
rect 3280 9928 3314 9944
rect 3280 9878 3314 9894
rect 4912 9928 4946 9944
rect 4912 9878 4946 9894
rect 6544 9928 6578 9944
rect 6544 9878 6578 9894
rect 8176 9928 8210 9944
rect 8176 9878 8210 9894
rect 9808 9928 9842 9944
rect 9808 9878 9842 9894
rect 16 9724 50 9740
rect 16 9674 50 9690
rect 1648 9724 1682 9740
rect 1648 9674 1682 9690
rect 3280 9724 3314 9740
rect 3280 9674 3314 9690
rect 4912 9724 4946 9740
rect 4912 9674 4946 9690
rect 6544 9724 6578 9740
rect 6544 9674 6578 9690
rect 8176 9724 8210 9740
rect 8176 9674 8210 9690
rect 9808 9724 9842 9740
rect 9808 9674 9842 9690
rect 211 9536 227 9570
rect 261 9536 277 9570
rect 415 9536 431 9570
rect 465 9536 481 9570
rect 619 9536 635 9570
rect 669 9536 685 9570
rect 823 9536 839 9570
rect 873 9536 889 9570
rect 1027 9536 1043 9570
rect 1077 9536 1093 9570
rect 1231 9536 1247 9570
rect 1281 9536 1297 9570
rect 1435 9536 1451 9570
rect 1485 9536 1501 9570
rect 1639 9536 1655 9570
rect 1689 9536 1705 9570
rect 1843 9536 1859 9570
rect 1893 9536 1909 9570
rect 2047 9536 2063 9570
rect 2097 9536 2113 9570
rect 2251 9536 2267 9570
rect 2301 9536 2317 9570
rect 2455 9536 2471 9570
rect 2505 9536 2521 9570
rect 2659 9536 2675 9570
rect 2709 9536 2725 9570
rect 2863 9536 2879 9570
rect 2913 9536 2929 9570
rect 3067 9536 3083 9570
rect 3117 9536 3133 9570
rect 3271 9536 3287 9570
rect 3321 9536 3337 9570
rect 3475 9536 3491 9570
rect 3525 9536 3541 9570
rect 3679 9536 3695 9570
rect 3729 9536 3745 9570
rect 3883 9536 3899 9570
rect 3933 9536 3949 9570
rect 4087 9536 4103 9570
rect 4137 9536 4153 9570
rect 4291 9536 4307 9570
rect 4341 9536 4357 9570
rect 4495 9536 4511 9570
rect 4545 9536 4561 9570
rect 4699 9536 4715 9570
rect 4749 9536 4765 9570
rect 4903 9536 4919 9570
rect 4953 9536 4969 9570
rect 5107 9536 5123 9570
rect 5157 9536 5173 9570
rect 5311 9536 5327 9570
rect 5361 9536 5377 9570
rect 5515 9536 5531 9570
rect 5565 9536 5581 9570
rect 5719 9536 5735 9570
rect 5769 9536 5785 9570
rect 5923 9536 5939 9570
rect 5973 9536 5989 9570
rect 6127 9536 6143 9570
rect 6177 9536 6193 9570
rect 6331 9536 6347 9570
rect 6381 9536 6397 9570
rect 6535 9536 6551 9570
rect 6585 9536 6601 9570
rect 6739 9536 6755 9570
rect 6789 9536 6805 9570
rect 6943 9536 6959 9570
rect 6993 9536 7009 9570
rect 7147 9536 7163 9570
rect 7197 9536 7213 9570
rect 7351 9536 7367 9570
rect 7401 9536 7417 9570
rect 7555 9536 7571 9570
rect 7605 9536 7621 9570
rect 7759 9536 7775 9570
rect 7809 9536 7825 9570
rect 7963 9536 7979 9570
rect 8013 9536 8029 9570
rect 8167 9536 8183 9570
rect 8217 9536 8233 9570
rect 8371 9536 8387 9570
rect 8421 9536 8437 9570
rect 8575 9536 8591 9570
rect 8625 9536 8641 9570
rect 8779 9536 8795 9570
rect 8829 9536 8845 9570
rect 8983 9536 8999 9570
rect 9033 9536 9049 9570
rect 9187 9536 9203 9570
rect 9237 9536 9253 9570
rect 9391 9536 9407 9570
rect 9441 9536 9457 9570
rect 9595 9536 9611 9570
rect 9645 9536 9661 9570
rect 9813 9536 9829 9570
rect 9863 9536 9879 9570
rect 16 9416 50 9432
rect 16 9366 50 9382
rect 1648 9416 1682 9432
rect 1648 9366 1682 9382
rect 3280 9416 3314 9432
rect 3280 9366 3314 9382
rect 4912 9416 4946 9432
rect 4912 9366 4946 9382
rect 6544 9416 6578 9432
rect 6544 9366 6578 9382
rect 8176 9416 8210 9432
rect 8176 9366 8210 9382
rect 9808 9416 9842 9432
rect 9808 9366 9842 9382
rect 16 9212 50 9228
rect 16 9162 50 9178
rect 1648 9212 1682 9228
rect 1648 9162 1682 9178
rect 3280 9212 3314 9228
rect 3280 9162 3314 9178
rect 4912 9212 4946 9228
rect 4912 9162 4946 9178
rect 6544 9212 6578 9228
rect 6544 9162 6578 9178
rect 8176 9212 8210 9228
rect 8176 9162 8210 9178
rect 9808 9212 9842 9228
rect 9808 9162 9842 9178
rect 16 9008 50 9024
rect 16 8958 50 8974
rect 1648 9008 1682 9024
rect 1648 8958 1682 8974
rect 3280 9008 3314 9024
rect 3280 8958 3314 8974
rect 4912 9008 4946 9024
rect 4912 8958 4946 8974
rect 6544 9008 6578 9024
rect 6544 8958 6578 8974
rect 8176 9008 8210 9024
rect 8176 8958 8210 8974
rect 9808 9008 9842 9024
rect 9808 8958 9842 8974
rect 16 8804 50 8820
rect 16 8754 50 8770
rect 1648 8804 1682 8820
rect 1648 8754 1682 8770
rect 3280 8804 3314 8820
rect 3280 8754 3314 8770
rect 4912 8804 4946 8820
rect 4912 8754 4946 8770
rect 6544 8804 6578 8820
rect 6544 8754 6578 8770
rect 8176 8804 8210 8820
rect 8176 8754 8210 8770
rect 9808 8804 9842 8820
rect 9808 8754 9842 8770
rect 16 8600 50 8616
rect 16 8550 50 8566
rect 1648 8600 1682 8616
rect 1648 8550 1682 8566
rect 3280 8600 3314 8616
rect 3280 8550 3314 8566
rect 4912 8600 4946 8616
rect 4912 8550 4946 8566
rect 6544 8600 6578 8616
rect 6544 8550 6578 8566
rect 8176 8600 8210 8616
rect 8176 8550 8210 8566
rect 9808 8600 9842 8616
rect 9808 8550 9842 8566
rect 16 8396 50 8412
rect 16 8346 50 8362
rect 1648 8396 1682 8412
rect 1648 8346 1682 8362
rect 3280 8396 3314 8412
rect 3280 8346 3314 8362
rect 4912 8396 4946 8412
rect 4912 8346 4946 8362
rect 6544 8396 6578 8412
rect 6544 8346 6578 8362
rect 8176 8396 8210 8412
rect 8176 8346 8210 8362
rect 9808 8396 9842 8412
rect 9808 8346 9842 8362
rect 16 8192 50 8208
rect 16 8142 50 8158
rect 1648 8192 1682 8208
rect 1648 8142 1682 8158
rect 3280 8192 3314 8208
rect 3280 8142 3314 8158
rect 4912 8192 4946 8208
rect 4912 8142 4946 8158
rect 6544 8192 6578 8208
rect 6544 8142 6578 8158
rect 8176 8192 8210 8208
rect 8176 8142 8210 8158
rect 9808 8192 9842 8208
rect 9808 8142 9842 8158
rect 16 7988 50 8004
rect 16 7938 50 7954
rect 1648 7988 1682 8004
rect 1648 7938 1682 7954
rect 3280 7988 3314 8004
rect 3280 7938 3314 7954
rect 4912 7988 4946 8004
rect 4912 7938 4946 7954
rect 6544 7988 6578 8004
rect 6544 7938 6578 7954
rect 8176 7988 8210 8004
rect 8176 7938 8210 7954
rect 9808 7988 9842 8004
rect 9808 7938 9842 7954
rect 211 7800 227 7834
rect 261 7800 277 7834
rect 415 7800 431 7834
rect 465 7800 481 7834
rect 619 7800 635 7834
rect 669 7800 685 7834
rect 823 7800 839 7834
rect 873 7800 889 7834
rect 1027 7800 1043 7834
rect 1077 7800 1093 7834
rect 1231 7800 1247 7834
rect 1281 7800 1297 7834
rect 1435 7800 1451 7834
rect 1485 7800 1501 7834
rect 1639 7800 1655 7834
rect 1689 7800 1705 7834
rect 1843 7800 1859 7834
rect 1893 7800 1909 7834
rect 2047 7800 2063 7834
rect 2097 7800 2113 7834
rect 2251 7800 2267 7834
rect 2301 7800 2317 7834
rect 2455 7800 2471 7834
rect 2505 7800 2521 7834
rect 2659 7800 2675 7834
rect 2709 7800 2725 7834
rect 2863 7800 2879 7834
rect 2913 7800 2929 7834
rect 3067 7800 3083 7834
rect 3117 7800 3133 7834
rect 3271 7800 3287 7834
rect 3321 7800 3337 7834
rect 3475 7800 3491 7834
rect 3525 7800 3541 7834
rect 3679 7800 3695 7834
rect 3729 7800 3745 7834
rect 3883 7800 3899 7834
rect 3933 7800 3949 7834
rect 4087 7800 4103 7834
rect 4137 7800 4153 7834
rect 4291 7800 4307 7834
rect 4341 7800 4357 7834
rect 4495 7800 4511 7834
rect 4545 7800 4561 7834
rect 4699 7800 4715 7834
rect 4749 7800 4765 7834
rect 4903 7800 4919 7834
rect 4953 7800 4969 7834
rect 5107 7800 5123 7834
rect 5157 7800 5173 7834
rect 5311 7800 5327 7834
rect 5361 7800 5377 7834
rect 5515 7800 5531 7834
rect 5565 7800 5581 7834
rect 5719 7800 5735 7834
rect 5769 7800 5785 7834
rect 5923 7800 5939 7834
rect 5973 7800 5989 7834
rect 6127 7800 6143 7834
rect 6177 7800 6193 7834
rect 6331 7800 6347 7834
rect 6381 7800 6397 7834
rect 6535 7800 6551 7834
rect 6585 7800 6601 7834
rect 6739 7800 6755 7834
rect 6789 7800 6805 7834
rect 6943 7800 6959 7834
rect 6993 7800 7009 7834
rect 7147 7800 7163 7834
rect 7197 7800 7213 7834
rect 7351 7800 7367 7834
rect 7401 7800 7417 7834
rect 7555 7800 7571 7834
rect 7605 7800 7621 7834
rect 7759 7800 7775 7834
rect 7809 7800 7825 7834
rect 7963 7800 7979 7834
rect 8013 7800 8029 7834
rect 8167 7800 8183 7834
rect 8217 7800 8233 7834
rect 8371 7800 8387 7834
rect 8421 7800 8437 7834
rect 8575 7800 8591 7834
rect 8625 7800 8641 7834
rect 8779 7800 8795 7834
rect 8829 7800 8845 7834
rect 8983 7800 8999 7834
rect 9033 7800 9049 7834
rect 9187 7800 9203 7834
rect 9237 7800 9253 7834
rect 9391 7800 9407 7834
rect 9441 7800 9457 7834
rect 9595 7800 9611 7834
rect 9645 7800 9661 7834
rect 9813 7800 9829 7834
rect 9863 7800 9879 7834
rect 16 7680 50 7696
rect 16 7630 50 7646
rect 1648 7680 1682 7696
rect 1648 7630 1682 7646
rect 3280 7680 3314 7696
rect 3280 7630 3314 7646
rect 4912 7680 4946 7696
rect 4912 7630 4946 7646
rect 6544 7680 6578 7696
rect 6544 7630 6578 7646
rect 8176 7680 8210 7696
rect 8176 7630 8210 7646
rect 9808 7680 9842 7696
rect 9808 7630 9842 7646
rect 16 7476 50 7492
rect 16 7426 50 7442
rect 1648 7476 1682 7492
rect 1648 7426 1682 7442
rect 3280 7476 3314 7492
rect 3280 7426 3314 7442
rect 4912 7476 4946 7492
rect 4912 7426 4946 7442
rect 6544 7476 6578 7492
rect 6544 7426 6578 7442
rect 8176 7476 8210 7492
rect 8176 7426 8210 7442
rect 9808 7476 9842 7492
rect 9808 7426 9842 7442
rect 16 7272 50 7288
rect 16 7222 50 7238
rect 1648 7272 1682 7288
rect 1648 7222 1682 7238
rect 3280 7272 3314 7288
rect 3280 7222 3314 7238
rect 4912 7272 4946 7288
rect 4912 7222 4946 7238
rect 6544 7272 6578 7288
rect 6544 7222 6578 7238
rect 8176 7272 8210 7288
rect 8176 7222 8210 7238
rect 9808 7272 9842 7288
rect 9808 7222 9842 7238
rect 16 7068 50 7084
rect 16 7018 50 7034
rect 1648 7068 1682 7084
rect 1648 7018 1682 7034
rect 3280 7068 3314 7084
rect 3280 7018 3314 7034
rect 4912 7068 4946 7084
rect 4912 7018 4946 7034
rect 6544 7068 6578 7084
rect 6544 7018 6578 7034
rect 8176 7068 8210 7084
rect 8176 7018 8210 7034
rect 9808 7068 9842 7084
rect 9808 7018 9842 7034
rect 16 6864 50 6880
rect 16 6814 50 6830
rect 1648 6864 1682 6880
rect 1648 6814 1682 6830
rect 3280 6864 3314 6880
rect 3280 6814 3314 6830
rect 4912 6864 4946 6880
rect 4912 6814 4946 6830
rect 6544 6864 6578 6880
rect 6544 6814 6578 6830
rect 8176 6864 8210 6880
rect 8176 6814 8210 6830
rect 9808 6864 9842 6880
rect 9808 6814 9842 6830
rect 16 6660 50 6676
rect 16 6610 50 6626
rect 1648 6660 1682 6676
rect 1648 6610 1682 6626
rect 3280 6660 3314 6676
rect 3280 6610 3314 6626
rect 4912 6660 4946 6676
rect 4912 6610 4946 6626
rect 6544 6660 6578 6676
rect 6544 6610 6578 6626
rect 8176 6660 8210 6676
rect 8176 6610 8210 6626
rect 9808 6660 9842 6676
rect 9808 6610 9842 6626
rect 16 6456 50 6472
rect 16 6406 50 6422
rect 1648 6456 1682 6472
rect 1648 6406 1682 6422
rect 3280 6456 3314 6472
rect 3280 6406 3314 6422
rect 4912 6456 4946 6472
rect 4912 6406 4946 6422
rect 6544 6456 6578 6472
rect 6544 6406 6578 6422
rect 8176 6456 8210 6472
rect 8176 6406 8210 6422
rect 9808 6456 9842 6472
rect 9808 6406 9842 6422
rect 16 6252 50 6268
rect 16 6202 50 6218
rect 1648 6252 1682 6268
rect 1648 6202 1682 6218
rect 3280 6252 3314 6268
rect 3280 6202 3314 6218
rect 4912 6252 4946 6268
rect 4912 6202 4946 6218
rect 6544 6252 6578 6268
rect 6544 6202 6578 6218
rect 8176 6252 8210 6268
rect 8176 6202 8210 6218
rect 9808 6252 9842 6268
rect 9808 6202 9842 6218
rect 211 6064 227 6098
rect 261 6064 277 6098
rect 415 6064 431 6098
rect 465 6064 481 6098
rect 619 6064 635 6098
rect 669 6064 685 6098
rect 823 6064 839 6098
rect 873 6064 889 6098
rect 1027 6064 1043 6098
rect 1077 6064 1093 6098
rect 1231 6064 1247 6098
rect 1281 6064 1297 6098
rect 1435 6064 1451 6098
rect 1485 6064 1501 6098
rect 1639 6064 1655 6098
rect 1689 6064 1705 6098
rect 1843 6064 1859 6098
rect 1893 6064 1909 6098
rect 2047 6064 2063 6098
rect 2097 6064 2113 6098
rect 2251 6064 2267 6098
rect 2301 6064 2317 6098
rect 2455 6064 2471 6098
rect 2505 6064 2521 6098
rect 2659 6064 2675 6098
rect 2709 6064 2725 6098
rect 2863 6064 2879 6098
rect 2913 6064 2929 6098
rect 3067 6064 3083 6098
rect 3117 6064 3133 6098
rect 3271 6064 3287 6098
rect 3321 6064 3337 6098
rect 3475 6064 3491 6098
rect 3525 6064 3541 6098
rect 3679 6064 3695 6098
rect 3729 6064 3745 6098
rect 3883 6064 3899 6098
rect 3933 6064 3949 6098
rect 4087 6064 4103 6098
rect 4137 6064 4153 6098
rect 4291 6064 4307 6098
rect 4341 6064 4357 6098
rect 4495 6064 4511 6098
rect 4545 6064 4561 6098
rect 4699 6064 4715 6098
rect 4749 6064 4765 6098
rect 4903 6064 4919 6098
rect 4953 6064 4969 6098
rect 5107 6064 5123 6098
rect 5157 6064 5173 6098
rect 5311 6064 5327 6098
rect 5361 6064 5377 6098
rect 5515 6064 5531 6098
rect 5565 6064 5581 6098
rect 5719 6064 5735 6098
rect 5769 6064 5785 6098
rect 5923 6064 5939 6098
rect 5973 6064 5989 6098
rect 6127 6064 6143 6098
rect 6177 6064 6193 6098
rect 6331 6064 6347 6098
rect 6381 6064 6397 6098
rect 6535 6064 6551 6098
rect 6585 6064 6601 6098
rect 6739 6064 6755 6098
rect 6789 6064 6805 6098
rect 6943 6064 6959 6098
rect 6993 6064 7009 6098
rect 7147 6064 7163 6098
rect 7197 6064 7213 6098
rect 7351 6064 7367 6098
rect 7401 6064 7417 6098
rect 7555 6064 7571 6098
rect 7605 6064 7621 6098
rect 7759 6064 7775 6098
rect 7809 6064 7825 6098
rect 7963 6064 7979 6098
rect 8013 6064 8029 6098
rect 8167 6064 8183 6098
rect 8217 6064 8233 6098
rect 8371 6064 8387 6098
rect 8421 6064 8437 6098
rect 8575 6064 8591 6098
rect 8625 6064 8641 6098
rect 8779 6064 8795 6098
rect 8829 6064 8845 6098
rect 8983 6064 8999 6098
rect 9033 6064 9049 6098
rect 9187 6064 9203 6098
rect 9237 6064 9253 6098
rect 9391 6064 9407 6098
rect 9441 6064 9457 6098
rect 9595 6064 9611 6098
rect 9645 6064 9661 6098
rect 9813 6064 9829 6098
rect 9863 6064 9879 6098
rect 16 5944 50 5960
rect 16 5894 50 5910
rect 1648 5944 1682 5960
rect 1648 5894 1682 5910
rect 3280 5944 3314 5960
rect 3280 5894 3314 5910
rect 4912 5944 4946 5960
rect 4912 5894 4946 5910
rect 6544 5944 6578 5960
rect 6544 5894 6578 5910
rect 8176 5944 8210 5960
rect 8176 5894 8210 5910
rect 9808 5944 9842 5960
rect 9808 5894 9842 5910
rect 16 5740 50 5756
rect 16 5690 50 5706
rect 1648 5740 1682 5756
rect 1648 5690 1682 5706
rect 3280 5740 3314 5756
rect 3280 5690 3314 5706
rect 4912 5740 4946 5756
rect 4912 5690 4946 5706
rect 6544 5740 6578 5756
rect 6544 5690 6578 5706
rect 8176 5740 8210 5756
rect 8176 5690 8210 5706
rect 9808 5740 9842 5756
rect 9808 5690 9842 5706
rect 16 5536 50 5552
rect 16 5486 50 5502
rect 1648 5536 1682 5552
rect 1648 5486 1682 5502
rect 3280 5536 3314 5552
rect 3280 5486 3314 5502
rect 4912 5536 4946 5552
rect 4912 5486 4946 5502
rect 6544 5536 6578 5552
rect 6544 5486 6578 5502
rect 8176 5536 8210 5552
rect 8176 5486 8210 5502
rect 9808 5536 9842 5552
rect 9808 5486 9842 5502
rect 16 5332 50 5348
rect 16 5282 50 5298
rect 1648 5332 1682 5348
rect 1648 5282 1682 5298
rect 3280 5332 3314 5348
rect 3280 5282 3314 5298
rect 4912 5332 4946 5348
rect 4912 5282 4946 5298
rect 6544 5332 6578 5348
rect 6544 5282 6578 5298
rect 8176 5332 8210 5348
rect 8176 5282 8210 5298
rect 9808 5332 9842 5348
rect 9808 5282 9842 5298
rect 16 5128 50 5144
rect 16 5078 50 5094
rect 1648 5128 1682 5144
rect 1648 5078 1682 5094
rect 3280 5128 3314 5144
rect 3280 5078 3314 5094
rect 4912 5128 4946 5144
rect 4912 5078 4946 5094
rect 6544 5128 6578 5144
rect 6544 5078 6578 5094
rect 8176 5128 8210 5144
rect 8176 5078 8210 5094
rect 9808 5128 9842 5144
rect 9808 5078 9842 5094
rect 16 4924 50 4940
rect 16 4874 50 4890
rect 1648 4924 1682 4940
rect 1648 4874 1682 4890
rect 3280 4924 3314 4940
rect 3280 4874 3314 4890
rect 4912 4924 4946 4940
rect 4912 4874 4946 4890
rect 6544 4924 6578 4940
rect 6544 4874 6578 4890
rect 8176 4924 8210 4940
rect 8176 4874 8210 4890
rect 9808 4924 9842 4940
rect 9808 4874 9842 4890
rect 16 4720 50 4736
rect 16 4670 50 4686
rect 1648 4720 1682 4736
rect 1648 4670 1682 4686
rect 3280 4720 3314 4736
rect 3280 4670 3314 4686
rect 4912 4720 4946 4736
rect 4912 4670 4946 4686
rect 6544 4720 6578 4736
rect 6544 4670 6578 4686
rect 8176 4720 8210 4736
rect 8176 4670 8210 4686
rect 9808 4720 9842 4736
rect 9808 4670 9842 4686
rect 16 4516 50 4532
rect 16 4466 50 4482
rect 1648 4516 1682 4532
rect 1648 4466 1682 4482
rect 3280 4516 3314 4532
rect 3280 4466 3314 4482
rect 4912 4516 4946 4532
rect 4912 4466 4946 4482
rect 6544 4516 6578 4532
rect 6544 4466 6578 4482
rect 8176 4516 8210 4532
rect 8176 4466 8210 4482
rect 9808 4516 9842 4532
rect 9808 4466 9842 4482
rect 211 4328 227 4362
rect 261 4328 277 4362
rect 415 4328 431 4362
rect 465 4328 481 4362
rect 619 4328 635 4362
rect 669 4328 685 4362
rect 823 4328 839 4362
rect 873 4328 889 4362
rect 1027 4328 1043 4362
rect 1077 4328 1093 4362
rect 1231 4328 1247 4362
rect 1281 4328 1297 4362
rect 1435 4328 1451 4362
rect 1485 4328 1501 4362
rect 1639 4328 1655 4362
rect 1689 4328 1705 4362
rect 1843 4328 1859 4362
rect 1893 4328 1909 4362
rect 2047 4328 2063 4362
rect 2097 4328 2113 4362
rect 2251 4328 2267 4362
rect 2301 4328 2317 4362
rect 2455 4328 2471 4362
rect 2505 4328 2521 4362
rect 2659 4328 2675 4362
rect 2709 4328 2725 4362
rect 2863 4328 2879 4362
rect 2913 4328 2929 4362
rect 3067 4328 3083 4362
rect 3117 4328 3133 4362
rect 3271 4328 3287 4362
rect 3321 4328 3337 4362
rect 3475 4328 3491 4362
rect 3525 4328 3541 4362
rect 3679 4328 3695 4362
rect 3729 4328 3745 4362
rect 3883 4328 3899 4362
rect 3933 4328 3949 4362
rect 4087 4328 4103 4362
rect 4137 4328 4153 4362
rect 4291 4328 4307 4362
rect 4341 4328 4357 4362
rect 4495 4328 4511 4362
rect 4545 4328 4561 4362
rect 4699 4328 4715 4362
rect 4749 4328 4765 4362
rect 4903 4328 4919 4362
rect 4953 4328 4969 4362
rect 5107 4328 5123 4362
rect 5157 4328 5173 4362
rect 5311 4328 5327 4362
rect 5361 4328 5377 4362
rect 5515 4328 5531 4362
rect 5565 4328 5581 4362
rect 5719 4328 5735 4362
rect 5769 4328 5785 4362
rect 5923 4328 5939 4362
rect 5973 4328 5989 4362
rect 6127 4328 6143 4362
rect 6177 4328 6193 4362
rect 6331 4328 6347 4362
rect 6381 4328 6397 4362
rect 6535 4328 6551 4362
rect 6585 4328 6601 4362
rect 6739 4328 6755 4362
rect 6789 4328 6805 4362
rect 6943 4328 6959 4362
rect 6993 4328 7009 4362
rect 7147 4328 7163 4362
rect 7197 4328 7213 4362
rect 7351 4328 7367 4362
rect 7401 4328 7417 4362
rect 7555 4328 7571 4362
rect 7605 4328 7621 4362
rect 7759 4328 7775 4362
rect 7809 4328 7825 4362
rect 7963 4328 7979 4362
rect 8013 4328 8029 4362
rect 8167 4328 8183 4362
rect 8217 4328 8233 4362
rect 8371 4328 8387 4362
rect 8421 4328 8437 4362
rect 8575 4328 8591 4362
rect 8625 4328 8641 4362
rect 8779 4328 8795 4362
rect 8829 4328 8845 4362
rect 8983 4328 8999 4362
rect 9033 4328 9049 4362
rect 9187 4328 9203 4362
rect 9237 4328 9253 4362
rect 9391 4328 9407 4362
rect 9441 4328 9457 4362
rect 9595 4328 9611 4362
rect 9645 4328 9661 4362
rect 9813 4328 9829 4362
rect 9863 4328 9879 4362
rect 16 4208 50 4224
rect 16 4158 50 4174
rect 1648 4208 1682 4224
rect 1648 4158 1682 4174
rect 3280 4208 3314 4224
rect 3280 4158 3314 4174
rect 4912 4208 4946 4224
rect 4912 4158 4946 4174
rect 6544 4208 6578 4224
rect 6544 4158 6578 4174
rect 8176 4208 8210 4224
rect 8176 4158 8210 4174
rect 9808 4208 9842 4224
rect 9808 4158 9842 4174
rect 16 4004 50 4020
rect 16 3954 50 3970
rect 1648 4004 1682 4020
rect 1648 3954 1682 3970
rect 3280 4004 3314 4020
rect 3280 3954 3314 3970
rect 4912 4004 4946 4020
rect 4912 3954 4946 3970
rect 6544 4004 6578 4020
rect 6544 3954 6578 3970
rect 8176 4004 8210 4020
rect 8176 3954 8210 3970
rect 9808 4004 9842 4020
rect 9808 3954 9842 3970
rect 16 3800 50 3816
rect 16 3750 50 3766
rect 1648 3800 1682 3816
rect 1648 3750 1682 3766
rect 3280 3800 3314 3816
rect 3280 3750 3314 3766
rect 4912 3800 4946 3816
rect 4912 3750 4946 3766
rect 6544 3800 6578 3816
rect 6544 3750 6578 3766
rect 8176 3800 8210 3816
rect 8176 3750 8210 3766
rect 9808 3800 9842 3816
rect 9808 3750 9842 3766
rect 16 3596 50 3612
rect 16 3546 50 3562
rect 1648 3596 1682 3612
rect 1648 3546 1682 3562
rect 3280 3596 3314 3612
rect 3280 3546 3314 3562
rect 4912 3596 4946 3612
rect 4912 3546 4946 3562
rect 6544 3596 6578 3612
rect 6544 3546 6578 3562
rect 8176 3596 8210 3612
rect 8176 3546 8210 3562
rect 9808 3596 9842 3612
rect 9808 3546 9842 3562
rect 16 3392 50 3408
rect 16 3342 50 3358
rect 1648 3392 1682 3408
rect 1648 3342 1682 3358
rect 3280 3392 3314 3408
rect 3280 3342 3314 3358
rect 4912 3392 4946 3408
rect 4912 3342 4946 3358
rect 6544 3392 6578 3408
rect 6544 3342 6578 3358
rect 8176 3392 8210 3408
rect 8176 3342 8210 3358
rect 9808 3392 9842 3408
rect 9808 3342 9842 3358
rect 16 3188 50 3204
rect 16 3138 50 3154
rect 1648 3188 1682 3204
rect 1648 3138 1682 3154
rect 3280 3188 3314 3204
rect 3280 3138 3314 3154
rect 4912 3188 4946 3204
rect 4912 3138 4946 3154
rect 6544 3188 6578 3204
rect 6544 3138 6578 3154
rect 8176 3188 8210 3204
rect 8176 3138 8210 3154
rect 9808 3188 9842 3204
rect 9808 3138 9842 3154
rect 16 2984 50 3000
rect 16 2934 50 2950
rect 1648 2984 1682 3000
rect 1648 2934 1682 2950
rect 3280 2984 3314 3000
rect 3280 2934 3314 2950
rect 4912 2984 4946 3000
rect 4912 2934 4946 2950
rect 6544 2984 6578 3000
rect 6544 2934 6578 2950
rect 8176 2984 8210 3000
rect 8176 2934 8210 2950
rect 9808 2984 9842 3000
rect 9808 2934 9842 2950
rect 16 2780 50 2796
rect 16 2730 50 2746
rect 1648 2780 1682 2796
rect 1648 2730 1682 2746
rect 3280 2780 3314 2796
rect 3280 2730 3314 2746
rect 4912 2780 4946 2796
rect 4912 2730 4946 2746
rect 6544 2780 6578 2796
rect 6544 2730 6578 2746
rect 8176 2780 8210 2796
rect 8176 2730 8210 2746
rect 9808 2780 9842 2796
rect 9808 2730 9842 2746
rect 211 2592 227 2626
rect 261 2592 277 2626
rect 415 2592 431 2626
rect 465 2592 481 2626
rect 619 2592 635 2626
rect 669 2592 685 2626
rect 823 2592 839 2626
rect 873 2592 889 2626
rect 1027 2592 1043 2626
rect 1077 2592 1093 2626
rect 1231 2592 1247 2626
rect 1281 2592 1297 2626
rect 1435 2592 1451 2626
rect 1485 2592 1501 2626
rect 1639 2592 1655 2626
rect 1689 2592 1705 2626
rect 1843 2592 1859 2626
rect 1893 2592 1909 2626
rect 2047 2592 2063 2626
rect 2097 2592 2113 2626
rect 2251 2592 2267 2626
rect 2301 2592 2317 2626
rect 2455 2592 2471 2626
rect 2505 2592 2521 2626
rect 2659 2592 2675 2626
rect 2709 2592 2725 2626
rect 2863 2592 2879 2626
rect 2913 2592 2929 2626
rect 3067 2592 3083 2626
rect 3117 2592 3133 2626
rect 3271 2592 3287 2626
rect 3321 2592 3337 2626
rect 3475 2592 3491 2626
rect 3525 2592 3541 2626
rect 3679 2592 3695 2626
rect 3729 2592 3745 2626
rect 3883 2592 3899 2626
rect 3933 2592 3949 2626
rect 4087 2592 4103 2626
rect 4137 2592 4153 2626
rect 4291 2592 4307 2626
rect 4341 2592 4357 2626
rect 4495 2592 4511 2626
rect 4545 2592 4561 2626
rect 4699 2592 4715 2626
rect 4749 2592 4765 2626
rect 4903 2592 4919 2626
rect 4953 2592 4969 2626
rect 5107 2592 5123 2626
rect 5157 2592 5173 2626
rect 5311 2592 5327 2626
rect 5361 2592 5377 2626
rect 5515 2592 5531 2626
rect 5565 2592 5581 2626
rect 5719 2592 5735 2626
rect 5769 2592 5785 2626
rect 5923 2592 5939 2626
rect 5973 2592 5989 2626
rect 6127 2592 6143 2626
rect 6177 2592 6193 2626
rect 6331 2592 6347 2626
rect 6381 2592 6397 2626
rect 6535 2592 6551 2626
rect 6585 2592 6601 2626
rect 6739 2592 6755 2626
rect 6789 2592 6805 2626
rect 6943 2592 6959 2626
rect 6993 2592 7009 2626
rect 7147 2592 7163 2626
rect 7197 2592 7213 2626
rect 7351 2592 7367 2626
rect 7401 2592 7417 2626
rect 7555 2592 7571 2626
rect 7605 2592 7621 2626
rect 7759 2592 7775 2626
rect 7809 2592 7825 2626
rect 7963 2592 7979 2626
rect 8013 2592 8029 2626
rect 8167 2592 8183 2626
rect 8217 2592 8233 2626
rect 8371 2592 8387 2626
rect 8421 2592 8437 2626
rect 8575 2592 8591 2626
rect 8625 2592 8641 2626
rect 8779 2592 8795 2626
rect 8829 2592 8845 2626
rect 8983 2592 8999 2626
rect 9033 2592 9049 2626
rect 9187 2592 9203 2626
rect 9237 2592 9253 2626
rect 9391 2592 9407 2626
rect 9441 2592 9457 2626
rect 9595 2592 9611 2626
rect 9645 2592 9661 2626
rect 9813 2592 9829 2626
rect 9863 2592 9879 2626
rect 16 2472 50 2488
rect 16 2422 50 2438
rect 1648 2472 1682 2488
rect 1648 2422 1682 2438
rect 3280 2472 3314 2488
rect 3280 2422 3314 2438
rect 4912 2472 4946 2488
rect 4912 2422 4946 2438
rect 6544 2472 6578 2488
rect 6544 2422 6578 2438
rect 8176 2472 8210 2488
rect 8176 2422 8210 2438
rect 9808 2472 9842 2488
rect 9808 2422 9842 2438
rect 16 2268 50 2284
rect 16 2218 50 2234
rect 1648 2268 1682 2284
rect 1648 2218 1682 2234
rect 3280 2268 3314 2284
rect 3280 2218 3314 2234
rect 4912 2268 4946 2284
rect 4912 2218 4946 2234
rect 6544 2268 6578 2284
rect 6544 2218 6578 2234
rect 8176 2268 8210 2284
rect 8176 2218 8210 2234
rect 9808 2268 9842 2284
rect 9808 2218 9842 2234
rect 16 2064 50 2080
rect 16 2014 50 2030
rect 1648 2064 1682 2080
rect 1648 2014 1682 2030
rect 3280 2064 3314 2080
rect 3280 2014 3314 2030
rect 4912 2064 4946 2080
rect 4912 2014 4946 2030
rect 6544 2064 6578 2080
rect 6544 2014 6578 2030
rect 8176 2064 8210 2080
rect 8176 2014 8210 2030
rect 9808 2064 9842 2080
rect 9808 2014 9842 2030
rect 16 1860 50 1876
rect 16 1810 50 1826
rect 1648 1860 1682 1876
rect 1648 1810 1682 1826
rect 3280 1860 3314 1876
rect 3280 1810 3314 1826
rect 4912 1860 4946 1876
rect 4912 1810 4946 1826
rect 6544 1860 6578 1876
rect 6544 1810 6578 1826
rect 8176 1860 8210 1876
rect 8176 1810 8210 1826
rect 9808 1860 9842 1876
rect 9808 1810 9842 1826
rect 16 1656 50 1672
rect 16 1606 50 1622
rect 1648 1656 1682 1672
rect 1648 1606 1682 1622
rect 3280 1656 3314 1672
rect 3280 1606 3314 1622
rect 4912 1656 4946 1672
rect 4912 1606 4946 1622
rect 6544 1656 6578 1672
rect 6544 1606 6578 1622
rect 8176 1656 8210 1672
rect 8176 1606 8210 1622
rect 9808 1656 9842 1672
rect 9808 1606 9842 1622
rect 16 1452 50 1468
rect 16 1402 50 1418
rect 1648 1452 1682 1468
rect 1648 1402 1682 1418
rect 3280 1452 3314 1468
rect 3280 1402 3314 1418
rect 4912 1452 4946 1468
rect 4912 1402 4946 1418
rect 6544 1452 6578 1468
rect 6544 1402 6578 1418
rect 8176 1452 8210 1468
rect 8176 1402 8210 1418
rect 9808 1452 9842 1468
rect 9808 1402 9842 1418
rect 16 1248 50 1264
rect 16 1198 50 1214
rect 1648 1248 1682 1264
rect 1648 1198 1682 1214
rect 3280 1248 3314 1264
rect 3280 1198 3314 1214
rect 4912 1248 4946 1264
rect 4912 1198 4946 1214
rect 6544 1248 6578 1264
rect 6544 1198 6578 1214
rect 8176 1248 8210 1264
rect 8176 1198 8210 1214
rect 9808 1248 9842 1264
rect 9808 1198 9842 1214
rect 16 1044 50 1060
rect 16 994 50 1010
rect 1648 1044 1682 1060
rect 1648 994 1682 1010
rect 3280 1044 3314 1060
rect 3280 994 3314 1010
rect 4912 1044 4946 1060
rect 4912 994 4946 1010
rect 6544 1044 6578 1060
rect 6544 994 6578 1010
rect 8176 1044 8210 1060
rect 8176 994 8210 1010
rect 9808 1044 9842 1060
rect 9808 994 9842 1010
rect 211 856 227 890
rect 261 856 277 890
rect 415 856 431 890
rect 465 856 481 890
rect 619 856 635 890
rect 669 856 685 890
rect 823 856 839 890
rect 873 856 889 890
rect 1027 856 1043 890
rect 1077 856 1093 890
rect 1231 856 1247 890
rect 1281 856 1297 890
rect 1435 856 1451 890
rect 1485 856 1501 890
rect 1639 856 1655 890
rect 1689 856 1705 890
rect 1843 856 1859 890
rect 1893 856 1909 890
rect 2047 856 2063 890
rect 2097 856 2113 890
rect 2251 856 2267 890
rect 2301 856 2317 890
rect 2455 856 2471 890
rect 2505 856 2521 890
rect 2659 856 2675 890
rect 2709 856 2725 890
rect 2863 856 2879 890
rect 2913 856 2929 890
rect 3067 856 3083 890
rect 3117 856 3133 890
rect 3271 856 3287 890
rect 3321 856 3337 890
rect 3475 856 3491 890
rect 3525 856 3541 890
rect 3679 856 3695 890
rect 3729 856 3745 890
rect 3883 856 3899 890
rect 3933 856 3949 890
rect 4087 856 4103 890
rect 4137 856 4153 890
rect 4291 856 4307 890
rect 4341 856 4357 890
rect 4495 856 4511 890
rect 4545 856 4561 890
rect 4699 856 4715 890
rect 4749 856 4765 890
rect 4903 856 4919 890
rect 4953 856 4969 890
rect 5107 856 5123 890
rect 5157 856 5173 890
rect 5311 856 5327 890
rect 5361 856 5377 890
rect 5515 856 5531 890
rect 5565 856 5581 890
rect 5719 856 5735 890
rect 5769 856 5785 890
rect 5923 856 5939 890
rect 5973 856 5989 890
rect 6127 856 6143 890
rect 6177 856 6193 890
rect 6331 856 6347 890
rect 6381 856 6397 890
rect 6535 856 6551 890
rect 6585 856 6601 890
rect 6739 856 6755 890
rect 6789 856 6805 890
rect 6943 856 6959 890
rect 6993 856 7009 890
rect 7147 856 7163 890
rect 7197 856 7213 890
rect 7351 856 7367 890
rect 7401 856 7417 890
rect 7555 856 7571 890
rect 7605 856 7621 890
rect 7759 856 7775 890
rect 7809 856 7825 890
rect 7963 856 7979 890
rect 8013 856 8029 890
rect 8167 856 8183 890
rect 8217 856 8233 890
rect 8371 856 8387 890
rect 8421 856 8437 890
rect 8575 856 8591 890
rect 8625 856 8641 890
rect 8779 856 8795 890
rect 8829 856 8845 890
rect 8983 856 8999 890
rect 9033 856 9049 890
rect 9187 856 9203 890
rect 9237 856 9253 890
rect 9391 856 9407 890
rect 9441 856 9457 890
rect 9595 856 9611 890
rect 9645 856 9661 890
rect 9813 856 9829 890
rect 9863 856 9879 890
<< viali >>
rect 16 10098 50 10132
rect 1648 10098 1682 10132
rect 3280 10098 3314 10132
rect 4912 10098 4946 10132
rect 6544 10098 6578 10132
rect 8176 10098 8210 10132
rect 9808 10098 9842 10132
rect 16 9894 50 9928
rect 1648 9894 1682 9928
rect 3280 9894 3314 9928
rect 4912 9894 4946 9928
rect 6544 9894 6578 9928
rect 8176 9894 8210 9928
rect 9808 9894 9842 9928
rect 16 9690 50 9724
rect 1648 9690 1682 9724
rect 3280 9690 3314 9724
rect 4912 9690 4946 9724
rect 6544 9690 6578 9724
rect 8176 9690 8210 9724
rect 9808 9690 9842 9724
rect 227 9536 261 9570
rect 431 9536 465 9570
rect 635 9536 669 9570
rect 839 9536 873 9570
rect 1043 9536 1077 9570
rect 1247 9536 1281 9570
rect 1451 9536 1485 9570
rect 1655 9536 1689 9570
rect 1859 9536 1893 9570
rect 2063 9536 2097 9570
rect 2267 9536 2301 9570
rect 2471 9536 2505 9570
rect 2675 9536 2709 9570
rect 2879 9536 2913 9570
rect 3083 9536 3117 9570
rect 3287 9536 3321 9570
rect 3491 9536 3525 9570
rect 3695 9536 3729 9570
rect 3899 9536 3933 9570
rect 4103 9536 4137 9570
rect 4307 9536 4341 9570
rect 4511 9536 4545 9570
rect 4715 9536 4749 9570
rect 4919 9536 4953 9570
rect 5123 9536 5157 9570
rect 5327 9536 5361 9570
rect 5531 9536 5565 9570
rect 5735 9536 5769 9570
rect 5939 9536 5973 9570
rect 6143 9536 6177 9570
rect 6347 9536 6381 9570
rect 6551 9536 6585 9570
rect 6755 9536 6789 9570
rect 6959 9536 6993 9570
rect 7163 9536 7197 9570
rect 7367 9536 7401 9570
rect 7571 9536 7605 9570
rect 7775 9536 7809 9570
rect 7979 9536 8013 9570
rect 8183 9536 8217 9570
rect 8387 9536 8421 9570
rect 8591 9536 8625 9570
rect 8795 9536 8829 9570
rect 8999 9536 9033 9570
rect 9203 9536 9237 9570
rect 9407 9536 9441 9570
rect 9611 9536 9645 9570
rect 9829 9536 9863 9570
rect 16 9382 50 9416
rect 1648 9382 1682 9416
rect 3280 9382 3314 9416
rect 4912 9382 4946 9416
rect 6544 9382 6578 9416
rect 8176 9382 8210 9416
rect 9808 9382 9842 9416
rect 16 9178 50 9212
rect 1648 9178 1682 9212
rect 3280 9178 3314 9212
rect 4912 9178 4946 9212
rect 6544 9178 6578 9212
rect 8176 9178 8210 9212
rect 9808 9178 9842 9212
rect 16 8974 50 9008
rect 1648 8974 1682 9008
rect 3280 8974 3314 9008
rect 4912 8974 4946 9008
rect 6544 8974 6578 9008
rect 8176 8974 8210 9008
rect 9808 8974 9842 9008
rect 16 8770 50 8804
rect 1648 8770 1682 8804
rect 3280 8770 3314 8804
rect 4912 8770 4946 8804
rect 6544 8770 6578 8804
rect 8176 8770 8210 8804
rect 9808 8770 9842 8804
rect 16 8566 50 8600
rect 1648 8566 1682 8600
rect 3280 8566 3314 8600
rect 4912 8566 4946 8600
rect 6544 8566 6578 8600
rect 8176 8566 8210 8600
rect 9808 8566 9842 8600
rect 16 8362 50 8396
rect 1648 8362 1682 8396
rect 3280 8362 3314 8396
rect 4912 8362 4946 8396
rect 6544 8362 6578 8396
rect 8176 8362 8210 8396
rect 9808 8362 9842 8396
rect 16 8158 50 8192
rect 1648 8158 1682 8192
rect 3280 8158 3314 8192
rect 4912 8158 4946 8192
rect 6544 8158 6578 8192
rect 8176 8158 8210 8192
rect 9808 8158 9842 8192
rect 16 7954 50 7988
rect 1648 7954 1682 7988
rect 3280 7954 3314 7988
rect 4912 7954 4946 7988
rect 6544 7954 6578 7988
rect 8176 7954 8210 7988
rect 9808 7954 9842 7988
rect 227 7800 261 7834
rect 431 7800 465 7834
rect 635 7800 669 7834
rect 839 7800 873 7834
rect 1043 7800 1077 7834
rect 1247 7800 1281 7834
rect 1451 7800 1485 7834
rect 1655 7800 1689 7834
rect 1859 7800 1893 7834
rect 2063 7800 2097 7834
rect 2267 7800 2301 7834
rect 2471 7800 2505 7834
rect 2675 7800 2709 7834
rect 2879 7800 2913 7834
rect 3083 7800 3117 7834
rect 3287 7800 3321 7834
rect 3491 7800 3525 7834
rect 3695 7800 3729 7834
rect 3899 7800 3933 7834
rect 4103 7800 4137 7834
rect 4307 7800 4341 7834
rect 4511 7800 4545 7834
rect 4715 7800 4749 7834
rect 4919 7800 4953 7834
rect 5123 7800 5157 7834
rect 5327 7800 5361 7834
rect 5531 7800 5565 7834
rect 5735 7800 5769 7834
rect 5939 7800 5973 7834
rect 6143 7800 6177 7834
rect 6347 7800 6381 7834
rect 6551 7800 6585 7834
rect 6755 7800 6789 7834
rect 6959 7800 6993 7834
rect 7163 7800 7197 7834
rect 7367 7800 7401 7834
rect 7571 7800 7605 7834
rect 7775 7800 7809 7834
rect 7979 7800 8013 7834
rect 8183 7800 8217 7834
rect 8387 7800 8421 7834
rect 8591 7800 8625 7834
rect 8795 7800 8829 7834
rect 8999 7800 9033 7834
rect 9203 7800 9237 7834
rect 9407 7800 9441 7834
rect 9611 7800 9645 7834
rect 9829 7800 9863 7834
rect 16 7646 50 7680
rect 1648 7646 1682 7680
rect 3280 7646 3314 7680
rect 4912 7646 4946 7680
rect 6544 7646 6578 7680
rect 8176 7646 8210 7680
rect 9808 7646 9842 7680
rect 16 7442 50 7476
rect 1648 7442 1682 7476
rect 3280 7442 3314 7476
rect 4912 7442 4946 7476
rect 6544 7442 6578 7476
rect 8176 7442 8210 7476
rect 9808 7442 9842 7476
rect 16 7238 50 7272
rect 1648 7238 1682 7272
rect 3280 7238 3314 7272
rect 4912 7238 4946 7272
rect 6544 7238 6578 7272
rect 8176 7238 8210 7272
rect 9808 7238 9842 7272
rect 16 7034 50 7068
rect 1648 7034 1682 7068
rect 3280 7034 3314 7068
rect 4912 7034 4946 7068
rect 6544 7034 6578 7068
rect 8176 7034 8210 7068
rect 9808 7034 9842 7068
rect 16 6830 50 6864
rect 1648 6830 1682 6864
rect 3280 6830 3314 6864
rect 4912 6830 4946 6864
rect 6544 6830 6578 6864
rect 8176 6830 8210 6864
rect 9808 6830 9842 6864
rect 16 6626 50 6660
rect 1648 6626 1682 6660
rect 3280 6626 3314 6660
rect 4912 6626 4946 6660
rect 6544 6626 6578 6660
rect 8176 6626 8210 6660
rect 9808 6626 9842 6660
rect 16 6422 50 6456
rect 1648 6422 1682 6456
rect 3280 6422 3314 6456
rect 4912 6422 4946 6456
rect 6544 6422 6578 6456
rect 8176 6422 8210 6456
rect 9808 6422 9842 6456
rect 16 6218 50 6252
rect 1648 6218 1682 6252
rect 3280 6218 3314 6252
rect 4912 6218 4946 6252
rect 6544 6218 6578 6252
rect 8176 6218 8210 6252
rect 9808 6218 9842 6252
rect 227 6064 261 6098
rect 431 6064 465 6098
rect 635 6064 669 6098
rect 839 6064 873 6098
rect 1043 6064 1077 6098
rect 1247 6064 1281 6098
rect 1451 6064 1485 6098
rect 1655 6064 1689 6098
rect 1859 6064 1893 6098
rect 2063 6064 2097 6098
rect 2267 6064 2301 6098
rect 2471 6064 2505 6098
rect 2675 6064 2709 6098
rect 2879 6064 2913 6098
rect 3083 6064 3117 6098
rect 3287 6064 3321 6098
rect 3491 6064 3525 6098
rect 3695 6064 3729 6098
rect 3899 6064 3933 6098
rect 4103 6064 4137 6098
rect 4307 6064 4341 6098
rect 4511 6064 4545 6098
rect 4715 6064 4749 6098
rect 4919 6064 4953 6098
rect 5123 6064 5157 6098
rect 5327 6064 5361 6098
rect 5531 6064 5565 6098
rect 5735 6064 5769 6098
rect 5939 6064 5973 6098
rect 6143 6064 6177 6098
rect 6347 6064 6381 6098
rect 6551 6064 6585 6098
rect 6755 6064 6789 6098
rect 6959 6064 6993 6098
rect 7163 6064 7197 6098
rect 7367 6064 7401 6098
rect 7571 6064 7605 6098
rect 7775 6064 7809 6098
rect 7979 6064 8013 6098
rect 8183 6064 8217 6098
rect 8387 6064 8421 6098
rect 8591 6064 8625 6098
rect 8795 6064 8829 6098
rect 8999 6064 9033 6098
rect 9203 6064 9237 6098
rect 9407 6064 9441 6098
rect 9611 6064 9645 6098
rect 9829 6064 9863 6098
rect 16 5910 50 5944
rect 1648 5910 1682 5944
rect 3280 5910 3314 5944
rect 4912 5910 4946 5944
rect 6544 5910 6578 5944
rect 8176 5910 8210 5944
rect 9808 5910 9842 5944
rect 16 5706 50 5740
rect 1648 5706 1682 5740
rect 3280 5706 3314 5740
rect 4912 5706 4946 5740
rect 6544 5706 6578 5740
rect 8176 5706 8210 5740
rect 9808 5706 9842 5740
rect 16 5502 50 5536
rect 1648 5502 1682 5536
rect 3280 5502 3314 5536
rect 4912 5502 4946 5536
rect 6544 5502 6578 5536
rect 8176 5502 8210 5536
rect 9808 5502 9842 5536
rect 16 5298 50 5332
rect 1648 5298 1682 5332
rect 3280 5298 3314 5332
rect 4912 5298 4946 5332
rect 6544 5298 6578 5332
rect 8176 5298 8210 5332
rect 9808 5298 9842 5332
rect 16 5094 50 5128
rect 1648 5094 1682 5128
rect 3280 5094 3314 5128
rect 4912 5094 4946 5128
rect 6544 5094 6578 5128
rect 8176 5094 8210 5128
rect 9808 5094 9842 5128
rect 16 4890 50 4924
rect 1648 4890 1682 4924
rect 3280 4890 3314 4924
rect 4912 4890 4946 4924
rect 6544 4890 6578 4924
rect 8176 4890 8210 4924
rect 9808 4890 9842 4924
rect 16 4686 50 4720
rect 1648 4686 1682 4720
rect 3280 4686 3314 4720
rect 4912 4686 4946 4720
rect 6544 4686 6578 4720
rect 8176 4686 8210 4720
rect 9808 4686 9842 4720
rect 16 4482 50 4516
rect 1648 4482 1682 4516
rect 3280 4482 3314 4516
rect 4912 4482 4946 4516
rect 6544 4482 6578 4516
rect 8176 4482 8210 4516
rect 9808 4482 9842 4516
rect 227 4328 261 4362
rect 431 4328 465 4362
rect 635 4328 669 4362
rect 839 4328 873 4362
rect 1043 4328 1077 4362
rect 1247 4328 1281 4362
rect 1451 4328 1485 4362
rect 1655 4328 1689 4362
rect 1859 4328 1893 4362
rect 2063 4328 2097 4362
rect 2267 4328 2301 4362
rect 2471 4328 2505 4362
rect 2675 4328 2709 4362
rect 2879 4328 2913 4362
rect 3083 4328 3117 4362
rect 3287 4328 3321 4362
rect 3491 4328 3525 4362
rect 3695 4328 3729 4362
rect 3899 4328 3933 4362
rect 4103 4328 4137 4362
rect 4307 4328 4341 4362
rect 4511 4328 4545 4362
rect 4715 4328 4749 4362
rect 4919 4328 4953 4362
rect 5123 4328 5157 4362
rect 5327 4328 5361 4362
rect 5531 4328 5565 4362
rect 5735 4328 5769 4362
rect 5939 4328 5973 4362
rect 6143 4328 6177 4362
rect 6347 4328 6381 4362
rect 6551 4328 6585 4362
rect 6755 4328 6789 4362
rect 6959 4328 6993 4362
rect 7163 4328 7197 4362
rect 7367 4328 7401 4362
rect 7571 4328 7605 4362
rect 7775 4328 7809 4362
rect 7979 4328 8013 4362
rect 8183 4328 8217 4362
rect 8387 4328 8421 4362
rect 8591 4328 8625 4362
rect 8795 4328 8829 4362
rect 8999 4328 9033 4362
rect 9203 4328 9237 4362
rect 9407 4328 9441 4362
rect 9611 4328 9645 4362
rect 9829 4328 9863 4362
rect 16 4174 50 4208
rect 1648 4174 1682 4208
rect 3280 4174 3314 4208
rect 4912 4174 4946 4208
rect 6544 4174 6578 4208
rect 8176 4174 8210 4208
rect 9808 4174 9842 4208
rect 16 3970 50 4004
rect 1648 3970 1682 4004
rect 3280 3970 3314 4004
rect 4912 3970 4946 4004
rect 6544 3970 6578 4004
rect 8176 3970 8210 4004
rect 9808 3970 9842 4004
rect 16 3766 50 3800
rect 1648 3766 1682 3800
rect 3280 3766 3314 3800
rect 4912 3766 4946 3800
rect 6544 3766 6578 3800
rect 8176 3766 8210 3800
rect 9808 3766 9842 3800
rect 16 3562 50 3596
rect 1648 3562 1682 3596
rect 3280 3562 3314 3596
rect 4912 3562 4946 3596
rect 6544 3562 6578 3596
rect 8176 3562 8210 3596
rect 9808 3562 9842 3596
rect 16 3358 50 3392
rect 1648 3358 1682 3392
rect 3280 3358 3314 3392
rect 4912 3358 4946 3392
rect 6544 3358 6578 3392
rect 8176 3358 8210 3392
rect 9808 3358 9842 3392
rect 16 3154 50 3188
rect 1648 3154 1682 3188
rect 3280 3154 3314 3188
rect 4912 3154 4946 3188
rect 6544 3154 6578 3188
rect 8176 3154 8210 3188
rect 9808 3154 9842 3188
rect 16 2950 50 2984
rect 1648 2950 1682 2984
rect 3280 2950 3314 2984
rect 4912 2950 4946 2984
rect 6544 2950 6578 2984
rect 8176 2950 8210 2984
rect 9808 2950 9842 2984
rect 16 2746 50 2780
rect 1648 2746 1682 2780
rect 3280 2746 3314 2780
rect 4912 2746 4946 2780
rect 6544 2746 6578 2780
rect 8176 2746 8210 2780
rect 9808 2746 9842 2780
rect 227 2592 261 2626
rect 431 2592 465 2626
rect 635 2592 669 2626
rect 839 2592 873 2626
rect 1043 2592 1077 2626
rect 1247 2592 1281 2626
rect 1451 2592 1485 2626
rect 1655 2592 1689 2626
rect 1859 2592 1893 2626
rect 2063 2592 2097 2626
rect 2267 2592 2301 2626
rect 2471 2592 2505 2626
rect 2675 2592 2709 2626
rect 2879 2592 2913 2626
rect 3083 2592 3117 2626
rect 3287 2592 3321 2626
rect 3491 2592 3525 2626
rect 3695 2592 3729 2626
rect 3899 2592 3933 2626
rect 4103 2592 4137 2626
rect 4307 2592 4341 2626
rect 4511 2592 4545 2626
rect 4715 2592 4749 2626
rect 4919 2592 4953 2626
rect 5123 2592 5157 2626
rect 5327 2592 5361 2626
rect 5531 2592 5565 2626
rect 5735 2592 5769 2626
rect 5939 2592 5973 2626
rect 6143 2592 6177 2626
rect 6347 2592 6381 2626
rect 6551 2592 6585 2626
rect 6755 2592 6789 2626
rect 6959 2592 6993 2626
rect 7163 2592 7197 2626
rect 7367 2592 7401 2626
rect 7571 2592 7605 2626
rect 7775 2592 7809 2626
rect 7979 2592 8013 2626
rect 8183 2592 8217 2626
rect 8387 2592 8421 2626
rect 8591 2592 8625 2626
rect 8795 2592 8829 2626
rect 8999 2592 9033 2626
rect 9203 2592 9237 2626
rect 9407 2592 9441 2626
rect 9611 2592 9645 2626
rect 9829 2592 9863 2626
rect 16 2438 50 2472
rect 1648 2438 1682 2472
rect 3280 2438 3314 2472
rect 4912 2438 4946 2472
rect 6544 2438 6578 2472
rect 8176 2438 8210 2472
rect 9808 2438 9842 2472
rect 16 2234 50 2268
rect 1648 2234 1682 2268
rect 3280 2234 3314 2268
rect 4912 2234 4946 2268
rect 6544 2234 6578 2268
rect 8176 2234 8210 2268
rect 9808 2234 9842 2268
rect 16 2030 50 2064
rect 1648 2030 1682 2064
rect 3280 2030 3314 2064
rect 4912 2030 4946 2064
rect 6544 2030 6578 2064
rect 8176 2030 8210 2064
rect 9808 2030 9842 2064
rect 16 1826 50 1860
rect 1648 1826 1682 1860
rect 3280 1826 3314 1860
rect 4912 1826 4946 1860
rect 6544 1826 6578 1860
rect 8176 1826 8210 1860
rect 9808 1826 9842 1860
rect 16 1622 50 1656
rect 1648 1622 1682 1656
rect 3280 1622 3314 1656
rect 4912 1622 4946 1656
rect 6544 1622 6578 1656
rect 8176 1622 8210 1656
rect 9808 1622 9842 1656
rect 16 1418 50 1452
rect 1648 1418 1682 1452
rect 3280 1418 3314 1452
rect 4912 1418 4946 1452
rect 6544 1418 6578 1452
rect 8176 1418 8210 1452
rect 9808 1418 9842 1452
rect 16 1214 50 1248
rect 1648 1214 1682 1248
rect 3280 1214 3314 1248
rect 4912 1214 4946 1248
rect 6544 1214 6578 1248
rect 8176 1214 8210 1248
rect 9808 1214 9842 1248
rect 16 1010 50 1044
rect 1648 1010 1682 1044
rect 3280 1010 3314 1044
rect 4912 1010 4946 1044
rect 6544 1010 6578 1044
rect 8176 1010 8210 1044
rect 9808 1010 9842 1044
rect 227 856 261 890
rect 431 856 465 890
rect 635 856 669 890
rect 839 856 873 890
rect 1043 856 1077 890
rect 1247 856 1281 890
rect 1451 856 1485 890
rect 1655 856 1689 890
rect 1859 856 1893 890
rect 2063 856 2097 890
rect 2267 856 2301 890
rect 2471 856 2505 890
rect 2675 856 2709 890
rect 2879 856 2913 890
rect 3083 856 3117 890
rect 3287 856 3321 890
rect 3491 856 3525 890
rect 3695 856 3729 890
rect 3899 856 3933 890
rect 4103 856 4137 890
rect 4307 856 4341 890
rect 4511 856 4545 890
rect 4715 856 4749 890
rect 4919 856 4953 890
rect 5123 856 5157 890
rect 5327 856 5361 890
rect 5531 856 5565 890
rect 5735 856 5769 890
rect 5939 856 5973 890
rect 6143 856 6177 890
rect 6347 856 6381 890
rect 6551 856 6585 890
rect 6755 856 6789 890
rect 6959 856 6993 890
rect 7163 856 7197 890
rect 7367 856 7401 890
rect 7571 856 7605 890
rect 7775 856 7809 890
rect 7979 856 8013 890
rect 8183 856 8217 890
rect 8387 856 8421 890
rect 8591 856 8625 890
rect 8795 856 8829 890
rect 8999 856 9033 890
rect 9203 856 9237 890
rect 9407 856 9441 890
rect 9611 856 9645 890
rect 9829 856 9863 890
<< metal1 >>
rect 114 10228 9758 10256
rect 8 10141 59 10148
rect 1640 10141 1691 10148
rect 3272 10141 3323 10148
rect 4904 10141 4955 10148
rect 6536 10141 6587 10148
rect 8168 10141 8219 10148
rect 9800 10141 9851 10148
rect 1 10089 7 10141
rect 59 10089 65 10141
rect 1633 10089 1639 10141
rect 1691 10089 1697 10141
rect 3265 10089 3271 10141
rect 3323 10089 3329 10141
rect 4897 10089 4903 10141
rect 4955 10089 4961 10141
rect 6529 10089 6535 10141
rect 6587 10089 6593 10141
rect 8161 10089 8167 10141
rect 8219 10089 8225 10141
rect 9793 10089 9799 10141
rect 9851 10129 9857 10141
rect 9851 10101 10041 10129
rect 9851 10089 9857 10101
rect 8 10082 59 10089
rect 1640 10082 1691 10089
rect 3272 10082 3323 10089
rect 4904 10082 4955 10089
rect 6536 10082 6587 10089
rect 8168 10082 8219 10089
rect 9800 10082 9851 10089
rect 8 9937 59 9944
rect 1640 9937 1691 9944
rect 3272 9937 3323 9944
rect 4904 9937 4955 9944
rect 6536 9937 6587 9944
rect 8168 9937 8219 9944
rect 9800 9937 9851 9944
rect 1 9885 7 9937
rect 59 9885 65 9937
rect 1633 9885 1639 9937
rect 1691 9885 1697 9937
rect 3265 9885 3271 9937
rect 3323 9885 3329 9937
rect 4897 9885 4903 9937
rect 4955 9885 4961 9937
rect 6529 9885 6535 9937
rect 6587 9885 6593 9937
rect 8161 9885 8167 9937
rect 8219 9885 8225 9937
rect 9793 9885 9799 9937
rect 9851 9885 9857 9937
rect 8 9878 59 9885
rect 1640 9878 1691 9885
rect 3272 9878 3323 9885
rect 4904 9878 4955 9885
rect 6536 9878 6587 9885
rect 8168 9878 8219 9885
rect 9800 9878 9851 9885
rect 8 9733 59 9740
rect 1640 9733 1691 9740
rect 3272 9733 3323 9740
rect 4904 9733 4955 9740
rect 6536 9733 6587 9740
rect 8168 9733 8219 9740
rect 9800 9733 9851 9740
rect 1 9681 7 9733
rect 59 9681 65 9733
rect 1633 9681 1639 9733
rect 1691 9681 1697 9733
rect 3265 9681 3271 9733
rect 3323 9681 3329 9733
rect 4897 9681 4903 9733
rect 4955 9681 4961 9733
rect 6529 9681 6535 9733
rect 6587 9681 6593 9733
rect 8161 9681 8167 9733
rect 8219 9681 8225 9733
rect 9793 9681 9799 9733
rect 9851 9681 9857 9733
rect 8 9674 59 9681
rect 1640 9674 1691 9681
rect 3272 9674 3323 9681
rect 4904 9674 4955 9681
rect 6536 9674 6587 9681
rect 8168 9674 8219 9681
rect 9800 9674 9851 9681
rect 128 9449 156 9657
rect 218 9579 270 9585
rect 218 9521 270 9527
rect 332 9449 360 9657
rect 422 9579 474 9585
rect 422 9521 474 9527
rect 536 9449 564 9657
rect 626 9579 678 9585
rect 626 9521 678 9527
rect 740 9449 768 9657
rect 830 9579 882 9585
rect 830 9521 882 9527
rect 944 9449 972 9657
rect 1034 9579 1086 9585
rect 1034 9521 1086 9527
rect 1148 9449 1176 9657
rect 1238 9579 1290 9585
rect 1238 9521 1290 9527
rect 1352 9449 1380 9657
rect 1442 9579 1494 9585
rect 1442 9521 1494 9527
rect 1556 9449 1584 9657
rect 1646 9579 1698 9585
rect 1646 9521 1698 9527
rect 1760 9449 1788 9657
rect 1850 9579 1902 9585
rect 1850 9521 1902 9527
rect 1964 9449 1992 9657
rect 2054 9579 2106 9585
rect 2054 9521 2106 9527
rect 2168 9449 2196 9657
rect 2258 9579 2310 9585
rect 2258 9521 2310 9527
rect 2372 9449 2400 9657
rect 2462 9579 2514 9585
rect 2462 9521 2514 9527
rect 2576 9449 2604 9657
rect 2666 9579 2718 9585
rect 2666 9521 2718 9527
rect 2780 9449 2808 9657
rect 2870 9579 2922 9585
rect 2870 9521 2922 9527
rect 2984 9449 3012 9657
rect 3074 9579 3126 9585
rect 3074 9521 3126 9527
rect 3188 9449 3216 9657
rect 3278 9579 3330 9585
rect 3278 9521 3330 9527
rect 3392 9449 3420 9657
rect 3482 9579 3534 9585
rect 3482 9521 3534 9527
rect 3596 9449 3624 9657
rect 3686 9579 3738 9585
rect 3686 9521 3738 9527
rect 3800 9449 3828 9657
rect 3890 9579 3942 9585
rect 3890 9521 3942 9527
rect 4004 9449 4032 9657
rect 4094 9579 4146 9585
rect 4094 9521 4146 9527
rect 4208 9449 4236 9657
rect 4298 9579 4350 9585
rect 4298 9521 4350 9527
rect 4412 9449 4440 9657
rect 4502 9579 4554 9585
rect 4502 9521 4554 9527
rect 4616 9449 4644 9657
rect 4706 9579 4758 9585
rect 4706 9521 4758 9527
rect 4820 9449 4848 9657
rect 4910 9579 4962 9585
rect 4910 9521 4962 9527
rect 5024 9449 5052 9657
rect 5114 9579 5166 9585
rect 5114 9521 5166 9527
rect 5228 9449 5256 9657
rect 5318 9579 5370 9585
rect 5318 9521 5370 9527
rect 5432 9449 5460 9657
rect 5522 9579 5574 9585
rect 5522 9521 5574 9527
rect 5636 9449 5664 9657
rect 5726 9579 5778 9585
rect 5726 9521 5778 9527
rect 5840 9449 5868 9657
rect 5930 9579 5982 9585
rect 5930 9521 5982 9527
rect 6044 9449 6072 9657
rect 6134 9579 6186 9585
rect 6134 9521 6186 9527
rect 6248 9449 6276 9657
rect 6338 9579 6390 9585
rect 6338 9521 6390 9527
rect 6452 9449 6480 9657
rect 6542 9579 6594 9585
rect 6542 9521 6594 9527
rect 6656 9449 6684 9657
rect 6746 9579 6798 9585
rect 6746 9521 6798 9527
rect 6860 9449 6888 9657
rect 6950 9579 7002 9585
rect 6950 9521 7002 9527
rect 7064 9449 7092 9657
rect 7154 9579 7206 9585
rect 7154 9521 7206 9527
rect 7268 9449 7296 9657
rect 7358 9579 7410 9585
rect 7358 9521 7410 9527
rect 7472 9449 7500 9657
rect 7562 9579 7614 9585
rect 7562 9521 7614 9527
rect 7676 9449 7704 9657
rect 7766 9579 7818 9585
rect 7766 9521 7818 9527
rect 7880 9449 7908 9657
rect 7970 9579 8022 9585
rect 7970 9521 8022 9527
rect 8084 9449 8112 9657
rect 8174 9579 8226 9585
rect 8174 9521 8226 9527
rect 8288 9449 8316 9657
rect 8378 9579 8430 9585
rect 8378 9521 8430 9527
rect 8492 9449 8520 9657
rect 8582 9579 8634 9585
rect 8582 9521 8634 9527
rect 8696 9449 8724 9657
rect 8786 9579 8838 9585
rect 8786 9521 8838 9527
rect 8900 9449 8928 9657
rect 8990 9579 9042 9585
rect 8990 9521 9042 9527
rect 9104 9449 9132 9657
rect 9194 9579 9246 9585
rect 9194 9521 9246 9527
rect 9308 9449 9336 9657
rect 9398 9579 9450 9585
rect 9398 9521 9450 9527
rect 9512 9449 9540 9657
rect 9602 9579 9654 9585
rect 9602 9521 9654 9527
rect 9716 9449 9744 9657
rect 9820 9579 9872 9585
rect 9820 9521 9872 9527
rect 8 9425 59 9432
rect 1640 9425 1691 9432
rect 3272 9425 3323 9432
rect 4904 9425 4955 9432
rect 6536 9425 6587 9432
rect 8168 9425 8219 9432
rect 9800 9425 9851 9432
rect 1 9373 7 9425
rect 59 9373 65 9425
rect 1633 9373 1639 9425
rect 1691 9373 1697 9425
rect 3265 9373 3271 9425
rect 3323 9373 3329 9425
rect 4897 9373 4903 9425
rect 4955 9373 4961 9425
rect 6529 9373 6535 9425
rect 6587 9373 6593 9425
rect 8161 9373 8167 9425
rect 8219 9373 8225 9425
rect 9793 9373 9799 9425
rect 9851 9373 9857 9425
rect 8 9366 59 9373
rect 1640 9366 1691 9373
rect 3272 9366 3323 9373
rect 4904 9366 4955 9373
rect 6536 9366 6587 9373
rect 8168 9366 8219 9373
rect 9800 9366 9851 9373
rect 8 9221 59 9228
rect 1640 9221 1691 9228
rect 3272 9221 3323 9228
rect 4904 9221 4955 9228
rect 6536 9221 6587 9228
rect 8168 9221 8219 9228
rect 9800 9221 9851 9228
rect 1 9169 7 9221
rect 59 9169 65 9221
rect 1633 9169 1639 9221
rect 1691 9169 1697 9221
rect 3265 9169 3271 9221
rect 3323 9169 3329 9221
rect 4897 9169 4903 9221
rect 4955 9169 4961 9221
rect 6529 9169 6535 9221
rect 6587 9169 6593 9221
rect 8161 9169 8167 9221
rect 8219 9169 8225 9221
rect 9793 9169 9799 9221
rect 9851 9169 9857 9221
rect 8 9162 59 9169
rect 1640 9162 1691 9169
rect 3272 9162 3323 9169
rect 4904 9162 4955 9169
rect 6536 9162 6587 9169
rect 8168 9162 8219 9169
rect 9800 9162 9851 9169
rect 8 9017 59 9024
rect 1640 9017 1691 9024
rect 3272 9017 3323 9024
rect 4904 9017 4955 9024
rect 6536 9017 6587 9024
rect 8168 9017 8219 9024
rect 9800 9017 9851 9024
rect 1 8965 7 9017
rect 59 8965 65 9017
rect 1633 8965 1639 9017
rect 1691 8965 1697 9017
rect 3265 8965 3271 9017
rect 3323 8965 3329 9017
rect 4897 8965 4903 9017
rect 4955 8965 4961 9017
rect 6529 8965 6535 9017
rect 6587 8965 6593 9017
rect 8161 8965 8167 9017
rect 8219 8965 8225 9017
rect 9793 8965 9799 9017
rect 9851 8965 9857 9017
rect 8 8958 59 8965
rect 1640 8958 1691 8965
rect 3272 8958 3323 8965
rect 4904 8958 4955 8965
rect 6536 8958 6587 8965
rect 8168 8958 8219 8965
rect 9800 8958 9851 8965
rect 8 8813 59 8820
rect 1640 8813 1691 8820
rect 3272 8813 3323 8820
rect 4904 8813 4955 8820
rect 6536 8813 6587 8820
rect 8168 8813 8219 8820
rect 9800 8813 9851 8820
rect 1 8761 7 8813
rect 59 8761 65 8813
rect 1633 8761 1639 8813
rect 1691 8761 1697 8813
rect 3265 8761 3271 8813
rect 3323 8761 3329 8813
rect 4897 8761 4903 8813
rect 4955 8761 4961 8813
rect 6529 8761 6535 8813
rect 6587 8761 6593 8813
rect 8161 8761 8167 8813
rect 8219 8761 8225 8813
rect 9793 8761 9799 8813
rect 9851 8761 9857 8813
rect 8 8754 59 8761
rect 1640 8754 1691 8761
rect 3272 8754 3323 8761
rect 4904 8754 4955 8761
rect 6536 8754 6587 8761
rect 8168 8754 8219 8761
rect 9800 8754 9851 8761
rect 8 8609 59 8616
rect 1640 8609 1691 8616
rect 3272 8609 3323 8616
rect 4904 8609 4955 8616
rect 6536 8609 6587 8616
rect 8168 8609 8219 8616
rect 9800 8609 9851 8616
rect 1 8557 7 8609
rect 59 8557 65 8609
rect 1633 8557 1639 8609
rect 1691 8557 1697 8609
rect 3265 8557 3271 8609
rect 3323 8557 3329 8609
rect 4897 8557 4903 8609
rect 4955 8557 4961 8609
rect 6529 8557 6535 8609
rect 6587 8557 6593 8609
rect 8161 8557 8167 8609
rect 8219 8557 8225 8609
rect 9793 8557 9799 8609
rect 9851 8557 9857 8609
rect 8 8550 59 8557
rect 1640 8550 1691 8557
rect 3272 8550 3323 8557
rect 4904 8550 4955 8557
rect 6536 8550 6587 8557
rect 8168 8550 8219 8557
rect 9800 8550 9851 8557
rect 8 8405 59 8412
rect 1640 8405 1691 8412
rect 3272 8405 3323 8412
rect 4904 8405 4955 8412
rect 6536 8405 6587 8412
rect 8168 8405 8219 8412
rect 9800 8405 9851 8412
rect 1 8353 7 8405
rect 59 8353 65 8405
rect 1633 8353 1639 8405
rect 1691 8353 1697 8405
rect 3265 8353 3271 8405
rect 3323 8353 3329 8405
rect 4897 8353 4903 8405
rect 4955 8353 4961 8405
rect 6529 8353 6535 8405
rect 6587 8353 6593 8405
rect 8161 8353 8167 8405
rect 8219 8353 8225 8405
rect 9793 8353 9799 8405
rect 9851 8353 9857 8405
rect 8 8346 59 8353
rect 1640 8346 1691 8353
rect 3272 8346 3323 8353
rect 4904 8346 4955 8353
rect 6536 8346 6587 8353
rect 8168 8346 8219 8353
rect 9800 8346 9851 8353
rect 8 8201 59 8208
rect 1640 8201 1691 8208
rect 3272 8201 3323 8208
rect 4904 8201 4955 8208
rect 6536 8201 6587 8208
rect 8168 8201 8219 8208
rect 9800 8201 9851 8208
rect 1 8149 7 8201
rect 59 8149 65 8201
rect 1633 8149 1639 8201
rect 1691 8149 1697 8201
rect 3265 8149 3271 8201
rect 3323 8149 3329 8201
rect 4897 8149 4903 8201
rect 4955 8149 4961 8201
rect 6529 8149 6535 8201
rect 6587 8149 6593 8201
rect 8161 8149 8167 8201
rect 8219 8149 8225 8201
rect 9793 8149 9799 8201
rect 9851 8149 9857 8201
rect 8 8142 59 8149
rect 1640 8142 1691 8149
rect 3272 8142 3323 8149
rect 4904 8142 4955 8149
rect 6536 8142 6587 8149
rect 8168 8142 8219 8149
rect 9800 8142 9851 8149
rect 8 7997 59 8004
rect 1640 7997 1691 8004
rect 3272 7997 3323 8004
rect 4904 7997 4955 8004
rect 6536 7997 6587 8004
rect 8168 7997 8219 8004
rect 9800 7997 9851 8004
rect 1 7945 7 7997
rect 59 7945 65 7997
rect 1633 7945 1639 7997
rect 1691 7945 1697 7997
rect 3265 7945 3271 7997
rect 3323 7945 3329 7997
rect 4897 7945 4903 7997
rect 4955 7945 4961 7997
rect 6529 7945 6535 7997
rect 6587 7945 6593 7997
rect 8161 7945 8167 7997
rect 8219 7945 8225 7997
rect 9793 7945 9799 7997
rect 9851 7945 9857 7997
rect 8 7938 59 7945
rect 1640 7938 1691 7945
rect 3272 7938 3323 7945
rect 4904 7938 4955 7945
rect 6536 7938 6587 7945
rect 8168 7938 8219 7945
rect 9800 7938 9851 7945
rect 128 7713 156 7921
rect 218 7843 270 7849
rect 218 7785 270 7791
rect 332 7713 360 7921
rect 422 7843 474 7849
rect 422 7785 474 7791
rect 536 7713 564 7921
rect 626 7843 678 7849
rect 626 7785 678 7791
rect 740 7713 768 7921
rect 830 7843 882 7849
rect 830 7785 882 7791
rect 944 7713 972 7921
rect 1034 7843 1086 7849
rect 1034 7785 1086 7791
rect 1148 7713 1176 7921
rect 1238 7843 1290 7849
rect 1238 7785 1290 7791
rect 1352 7713 1380 7921
rect 1442 7843 1494 7849
rect 1442 7785 1494 7791
rect 1556 7713 1584 7921
rect 1646 7843 1698 7849
rect 1646 7785 1698 7791
rect 1760 7713 1788 7921
rect 1850 7843 1902 7849
rect 1850 7785 1902 7791
rect 1964 7713 1992 7921
rect 2054 7843 2106 7849
rect 2054 7785 2106 7791
rect 2168 7713 2196 7921
rect 2258 7843 2310 7849
rect 2258 7785 2310 7791
rect 2372 7713 2400 7921
rect 2462 7843 2514 7849
rect 2462 7785 2514 7791
rect 2576 7713 2604 7921
rect 2666 7843 2718 7849
rect 2666 7785 2718 7791
rect 2780 7713 2808 7921
rect 2870 7843 2922 7849
rect 2870 7785 2922 7791
rect 2984 7713 3012 7921
rect 3074 7843 3126 7849
rect 3074 7785 3126 7791
rect 3188 7713 3216 7921
rect 3278 7843 3330 7849
rect 3278 7785 3330 7791
rect 3392 7713 3420 7921
rect 3482 7843 3534 7849
rect 3482 7785 3534 7791
rect 3596 7713 3624 7921
rect 3686 7843 3738 7849
rect 3686 7785 3738 7791
rect 3800 7713 3828 7921
rect 3890 7843 3942 7849
rect 3890 7785 3942 7791
rect 4004 7713 4032 7921
rect 4094 7843 4146 7849
rect 4094 7785 4146 7791
rect 4208 7713 4236 7921
rect 4298 7843 4350 7849
rect 4298 7785 4350 7791
rect 4412 7713 4440 7921
rect 4502 7843 4554 7849
rect 4502 7785 4554 7791
rect 4616 7713 4644 7921
rect 4706 7843 4758 7849
rect 4706 7785 4758 7791
rect 4820 7713 4848 7921
rect 4910 7843 4962 7849
rect 4910 7785 4962 7791
rect 5024 7713 5052 7921
rect 5114 7843 5166 7849
rect 5114 7785 5166 7791
rect 5228 7713 5256 7921
rect 5318 7843 5370 7849
rect 5318 7785 5370 7791
rect 5432 7713 5460 7921
rect 5522 7843 5574 7849
rect 5522 7785 5574 7791
rect 5636 7713 5664 7921
rect 5726 7843 5778 7849
rect 5726 7785 5778 7791
rect 5840 7713 5868 7921
rect 5930 7843 5982 7849
rect 5930 7785 5982 7791
rect 6044 7713 6072 7921
rect 6134 7843 6186 7849
rect 6134 7785 6186 7791
rect 6248 7713 6276 7921
rect 6338 7843 6390 7849
rect 6338 7785 6390 7791
rect 6452 7713 6480 7921
rect 6542 7843 6594 7849
rect 6542 7785 6594 7791
rect 6656 7713 6684 7921
rect 6746 7843 6798 7849
rect 6746 7785 6798 7791
rect 6860 7713 6888 7921
rect 6950 7843 7002 7849
rect 6950 7785 7002 7791
rect 7064 7713 7092 7921
rect 7154 7843 7206 7849
rect 7154 7785 7206 7791
rect 7268 7713 7296 7921
rect 7358 7843 7410 7849
rect 7358 7785 7410 7791
rect 7472 7713 7500 7921
rect 7562 7843 7614 7849
rect 7562 7785 7614 7791
rect 7676 7713 7704 7921
rect 7766 7843 7818 7849
rect 7766 7785 7818 7791
rect 7880 7713 7908 7921
rect 7970 7843 8022 7849
rect 7970 7785 8022 7791
rect 8084 7713 8112 7921
rect 8174 7843 8226 7849
rect 8174 7785 8226 7791
rect 8288 7713 8316 7921
rect 8378 7843 8430 7849
rect 8378 7785 8430 7791
rect 8492 7713 8520 7921
rect 8582 7843 8634 7849
rect 8582 7785 8634 7791
rect 8696 7713 8724 7921
rect 8786 7843 8838 7849
rect 8786 7785 8838 7791
rect 8900 7713 8928 7921
rect 8990 7843 9042 7849
rect 8990 7785 9042 7791
rect 9104 7713 9132 7921
rect 9194 7843 9246 7849
rect 9194 7785 9246 7791
rect 9308 7713 9336 7921
rect 9398 7843 9450 7849
rect 9398 7785 9450 7791
rect 9512 7713 9540 7921
rect 9602 7843 9654 7849
rect 9602 7785 9654 7791
rect 9716 7713 9744 7921
rect 9820 7843 9872 7849
rect 9820 7785 9872 7791
rect 8 7689 59 7696
rect 1640 7689 1691 7696
rect 3272 7689 3323 7696
rect 4904 7689 4955 7696
rect 6536 7689 6587 7696
rect 8168 7689 8219 7696
rect 9800 7689 9851 7696
rect 1 7637 7 7689
rect 59 7637 65 7689
rect 1633 7637 1639 7689
rect 1691 7637 1697 7689
rect 3265 7637 3271 7689
rect 3323 7637 3329 7689
rect 4897 7637 4903 7689
rect 4955 7637 4961 7689
rect 6529 7637 6535 7689
rect 6587 7637 6593 7689
rect 8161 7637 8167 7689
rect 8219 7637 8225 7689
rect 9793 7637 9799 7689
rect 9851 7637 9857 7689
rect 8 7630 59 7637
rect 1640 7630 1691 7637
rect 3272 7630 3323 7637
rect 4904 7630 4955 7637
rect 6536 7630 6587 7637
rect 8168 7630 8219 7637
rect 9800 7630 9851 7637
rect 8 7485 59 7492
rect 1640 7485 1691 7492
rect 3272 7485 3323 7492
rect 4904 7485 4955 7492
rect 6536 7485 6587 7492
rect 8168 7485 8219 7492
rect 9800 7485 9851 7492
rect 1 7433 7 7485
rect 59 7433 65 7485
rect 1633 7433 1639 7485
rect 1691 7433 1697 7485
rect 3265 7433 3271 7485
rect 3323 7433 3329 7485
rect 4897 7433 4903 7485
rect 4955 7433 4961 7485
rect 6529 7433 6535 7485
rect 6587 7433 6593 7485
rect 8161 7433 8167 7485
rect 8219 7433 8225 7485
rect 9793 7433 9799 7485
rect 9851 7433 9857 7485
rect 8 7426 59 7433
rect 1640 7426 1691 7433
rect 3272 7426 3323 7433
rect 4904 7426 4955 7433
rect 6536 7426 6587 7433
rect 8168 7426 8219 7433
rect 9800 7426 9851 7433
rect 8 7281 59 7288
rect 1640 7281 1691 7288
rect 3272 7281 3323 7288
rect 4904 7281 4955 7288
rect 6536 7281 6587 7288
rect 8168 7281 8219 7288
rect 9800 7281 9851 7288
rect 1 7229 7 7281
rect 59 7229 65 7281
rect 1633 7229 1639 7281
rect 1691 7229 1697 7281
rect 3265 7229 3271 7281
rect 3323 7229 3329 7281
rect 4897 7229 4903 7281
rect 4955 7229 4961 7281
rect 6529 7229 6535 7281
rect 6587 7229 6593 7281
rect 8161 7229 8167 7281
rect 8219 7229 8225 7281
rect 9793 7229 9799 7281
rect 9851 7229 9857 7281
rect 8 7222 59 7229
rect 1640 7222 1691 7229
rect 3272 7222 3323 7229
rect 4904 7222 4955 7229
rect 6536 7222 6587 7229
rect 8168 7222 8219 7229
rect 9800 7222 9851 7229
rect 8 7077 59 7084
rect 1640 7077 1691 7084
rect 3272 7077 3323 7084
rect 4904 7077 4955 7084
rect 6536 7077 6587 7084
rect 8168 7077 8219 7084
rect 9800 7077 9851 7084
rect 1 7025 7 7077
rect 59 7025 65 7077
rect 1633 7025 1639 7077
rect 1691 7025 1697 7077
rect 3265 7025 3271 7077
rect 3323 7025 3329 7077
rect 4897 7025 4903 7077
rect 4955 7025 4961 7077
rect 6529 7025 6535 7077
rect 6587 7025 6593 7077
rect 8161 7025 8167 7077
rect 8219 7025 8225 7077
rect 9793 7025 9799 7077
rect 9851 7025 9857 7077
rect 8 7018 59 7025
rect 1640 7018 1691 7025
rect 3272 7018 3323 7025
rect 4904 7018 4955 7025
rect 6536 7018 6587 7025
rect 8168 7018 8219 7025
rect 9800 7018 9851 7025
rect 8 6873 59 6880
rect 1640 6873 1691 6880
rect 3272 6873 3323 6880
rect 4904 6873 4955 6880
rect 6536 6873 6587 6880
rect 8168 6873 8219 6880
rect 9800 6873 9851 6880
rect 1 6821 7 6873
rect 59 6821 65 6873
rect 1633 6821 1639 6873
rect 1691 6821 1697 6873
rect 3265 6821 3271 6873
rect 3323 6821 3329 6873
rect 4897 6821 4903 6873
rect 4955 6821 4961 6873
rect 6529 6821 6535 6873
rect 6587 6821 6593 6873
rect 8161 6821 8167 6873
rect 8219 6821 8225 6873
rect 9793 6821 9799 6873
rect 9851 6821 9857 6873
rect 8 6814 59 6821
rect 1640 6814 1691 6821
rect 3272 6814 3323 6821
rect 4904 6814 4955 6821
rect 6536 6814 6587 6821
rect 8168 6814 8219 6821
rect 9800 6814 9851 6821
rect 8 6669 59 6676
rect 1640 6669 1691 6676
rect 3272 6669 3323 6676
rect 4904 6669 4955 6676
rect 6536 6669 6587 6676
rect 8168 6669 8219 6676
rect 9800 6669 9851 6676
rect 1 6617 7 6669
rect 59 6617 65 6669
rect 1633 6617 1639 6669
rect 1691 6617 1697 6669
rect 3265 6617 3271 6669
rect 3323 6617 3329 6669
rect 4897 6617 4903 6669
rect 4955 6617 4961 6669
rect 6529 6617 6535 6669
rect 6587 6617 6593 6669
rect 8161 6617 8167 6669
rect 8219 6617 8225 6669
rect 9793 6617 9799 6669
rect 9851 6617 9857 6669
rect 8 6610 59 6617
rect 1640 6610 1691 6617
rect 3272 6610 3323 6617
rect 4904 6610 4955 6617
rect 6536 6610 6587 6617
rect 8168 6610 8219 6617
rect 9800 6610 9851 6617
rect 8 6465 59 6472
rect 1640 6465 1691 6472
rect 3272 6465 3323 6472
rect 4904 6465 4955 6472
rect 6536 6465 6587 6472
rect 8168 6465 8219 6472
rect 9800 6465 9851 6472
rect 1 6413 7 6465
rect 59 6413 65 6465
rect 1633 6413 1639 6465
rect 1691 6413 1697 6465
rect 3265 6413 3271 6465
rect 3323 6413 3329 6465
rect 4897 6413 4903 6465
rect 4955 6413 4961 6465
rect 6529 6413 6535 6465
rect 6587 6413 6593 6465
rect 8161 6413 8167 6465
rect 8219 6413 8225 6465
rect 9793 6413 9799 6465
rect 9851 6413 9857 6465
rect 8 6406 59 6413
rect 1640 6406 1691 6413
rect 3272 6406 3323 6413
rect 4904 6406 4955 6413
rect 6536 6406 6587 6413
rect 8168 6406 8219 6413
rect 9800 6406 9851 6413
rect 8 6261 59 6268
rect 1640 6261 1691 6268
rect 3272 6261 3323 6268
rect 4904 6261 4955 6268
rect 6536 6261 6587 6268
rect 8168 6261 8219 6268
rect 9800 6261 9851 6268
rect 1 6209 7 6261
rect 59 6209 65 6261
rect 1633 6209 1639 6261
rect 1691 6209 1697 6261
rect 3265 6209 3271 6261
rect 3323 6209 3329 6261
rect 4897 6209 4903 6261
rect 4955 6209 4961 6261
rect 6529 6209 6535 6261
rect 6587 6209 6593 6261
rect 8161 6209 8167 6261
rect 8219 6209 8225 6261
rect 9793 6209 9799 6261
rect 9851 6209 9857 6261
rect 8 6202 59 6209
rect 1640 6202 1691 6209
rect 3272 6202 3323 6209
rect 4904 6202 4955 6209
rect 6536 6202 6587 6209
rect 8168 6202 8219 6209
rect 9800 6202 9851 6209
rect 128 5977 156 6185
rect 218 6107 270 6113
rect 218 6049 270 6055
rect 332 5977 360 6185
rect 422 6107 474 6113
rect 422 6049 474 6055
rect 536 5977 564 6185
rect 626 6107 678 6113
rect 626 6049 678 6055
rect 740 5977 768 6185
rect 830 6107 882 6113
rect 830 6049 882 6055
rect 944 5977 972 6185
rect 1034 6107 1086 6113
rect 1034 6049 1086 6055
rect 1148 5977 1176 6185
rect 1238 6107 1290 6113
rect 1238 6049 1290 6055
rect 1352 5977 1380 6185
rect 1442 6107 1494 6113
rect 1442 6049 1494 6055
rect 1556 5977 1584 6185
rect 1646 6107 1698 6113
rect 1646 6049 1698 6055
rect 1760 5977 1788 6185
rect 1850 6107 1902 6113
rect 1850 6049 1902 6055
rect 1964 5977 1992 6185
rect 2054 6107 2106 6113
rect 2054 6049 2106 6055
rect 2168 5977 2196 6185
rect 2258 6107 2310 6113
rect 2258 6049 2310 6055
rect 2372 5977 2400 6185
rect 2462 6107 2514 6113
rect 2462 6049 2514 6055
rect 2576 5977 2604 6185
rect 2666 6107 2718 6113
rect 2666 6049 2718 6055
rect 2780 5977 2808 6185
rect 2870 6107 2922 6113
rect 2870 6049 2922 6055
rect 2984 5977 3012 6185
rect 3074 6107 3126 6113
rect 3074 6049 3126 6055
rect 3188 5977 3216 6185
rect 3278 6107 3330 6113
rect 3278 6049 3330 6055
rect 3392 5977 3420 6185
rect 3482 6107 3534 6113
rect 3482 6049 3534 6055
rect 3596 5977 3624 6185
rect 3686 6107 3738 6113
rect 3686 6049 3738 6055
rect 3800 5977 3828 6185
rect 3890 6107 3942 6113
rect 3890 6049 3942 6055
rect 4004 5977 4032 6185
rect 4094 6107 4146 6113
rect 4094 6049 4146 6055
rect 4208 5977 4236 6185
rect 4298 6107 4350 6113
rect 4298 6049 4350 6055
rect 4412 5977 4440 6185
rect 4502 6107 4554 6113
rect 4502 6049 4554 6055
rect 4616 5977 4644 6185
rect 4706 6107 4758 6113
rect 4706 6049 4758 6055
rect 4820 5977 4848 6185
rect 4910 6107 4962 6113
rect 4910 6049 4962 6055
rect 5024 5977 5052 6185
rect 5114 6107 5166 6113
rect 5114 6049 5166 6055
rect 5228 5977 5256 6185
rect 5318 6107 5370 6113
rect 5318 6049 5370 6055
rect 5432 5977 5460 6185
rect 5522 6107 5574 6113
rect 5522 6049 5574 6055
rect 5636 5977 5664 6185
rect 5726 6107 5778 6113
rect 5726 6049 5778 6055
rect 5840 5977 5868 6185
rect 5930 6107 5982 6113
rect 5930 6049 5982 6055
rect 6044 5977 6072 6185
rect 6134 6107 6186 6113
rect 6134 6049 6186 6055
rect 6248 5977 6276 6185
rect 6338 6107 6390 6113
rect 6338 6049 6390 6055
rect 6452 5977 6480 6185
rect 6542 6107 6594 6113
rect 6542 6049 6594 6055
rect 6656 5977 6684 6185
rect 6746 6107 6798 6113
rect 6746 6049 6798 6055
rect 6860 5977 6888 6185
rect 6950 6107 7002 6113
rect 6950 6049 7002 6055
rect 7064 5977 7092 6185
rect 7154 6107 7206 6113
rect 7154 6049 7206 6055
rect 7268 5977 7296 6185
rect 7358 6107 7410 6113
rect 7358 6049 7410 6055
rect 7472 5977 7500 6185
rect 7562 6107 7614 6113
rect 7562 6049 7614 6055
rect 7676 5977 7704 6185
rect 7766 6107 7818 6113
rect 7766 6049 7818 6055
rect 7880 5977 7908 6185
rect 7970 6107 8022 6113
rect 7970 6049 8022 6055
rect 8084 5977 8112 6185
rect 8174 6107 8226 6113
rect 8174 6049 8226 6055
rect 8288 5977 8316 6185
rect 8378 6107 8430 6113
rect 8378 6049 8430 6055
rect 8492 5977 8520 6185
rect 8582 6107 8634 6113
rect 8582 6049 8634 6055
rect 8696 5977 8724 6185
rect 8786 6107 8838 6113
rect 8786 6049 8838 6055
rect 8900 5977 8928 6185
rect 8990 6107 9042 6113
rect 8990 6049 9042 6055
rect 9104 5977 9132 6185
rect 9194 6107 9246 6113
rect 9194 6049 9246 6055
rect 9308 5977 9336 6185
rect 9398 6107 9450 6113
rect 9398 6049 9450 6055
rect 9512 5977 9540 6185
rect 9602 6107 9654 6113
rect 9602 6049 9654 6055
rect 9716 5977 9744 6185
rect 9820 6107 9872 6113
rect 9820 6049 9872 6055
rect 8 5953 59 5960
rect 1640 5953 1691 5960
rect 3272 5953 3323 5960
rect 4904 5953 4955 5960
rect 6536 5953 6587 5960
rect 8168 5953 8219 5960
rect 9800 5953 9851 5960
rect 1 5901 7 5953
rect 59 5901 65 5953
rect 1633 5901 1639 5953
rect 1691 5901 1697 5953
rect 3265 5901 3271 5953
rect 3323 5901 3329 5953
rect 4897 5901 4903 5953
rect 4955 5901 4961 5953
rect 6529 5901 6535 5953
rect 6587 5901 6593 5953
rect 8161 5901 8167 5953
rect 8219 5901 8225 5953
rect 9793 5901 9799 5953
rect 9851 5901 9857 5953
rect 8 5894 59 5901
rect 1640 5894 1691 5901
rect 3272 5894 3323 5901
rect 4904 5894 4955 5901
rect 6536 5894 6587 5901
rect 8168 5894 8219 5901
rect 9800 5894 9851 5901
rect 8 5749 59 5756
rect 1640 5749 1691 5756
rect 3272 5749 3323 5756
rect 4904 5749 4955 5756
rect 6536 5749 6587 5756
rect 8168 5749 8219 5756
rect 9800 5749 9851 5756
rect 1 5697 7 5749
rect 59 5697 65 5749
rect 1633 5697 1639 5749
rect 1691 5697 1697 5749
rect 3265 5697 3271 5749
rect 3323 5697 3329 5749
rect 4897 5697 4903 5749
rect 4955 5697 4961 5749
rect 6529 5697 6535 5749
rect 6587 5697 6593 5749
rect 8161 5697 8167 5749
rect 8219 5697 8225 5749
rect 9793 5697 9799 5749
rect 9851 5697 9857 5749
rect 8 5690 59 5697
rect 1640 5690 1691 5697
rect 3272 5690 3323 5697
rect 4904 5690 4955 5697
rect 6536 5690 6587 5697
rect 8168 5690 8219 5697
rect 9800 5690 9851 5697
rect 8 5545 59 5552
rect 1640 5545 1691 5552
rect 3272 5545 3323 5552
rect 4904 5545 4955 5552
rect 6536 5545 6587 5552
rect 8168 5545 8219 5552
rect 9800 5545 9851 5552
rect 1 5493 7 5545
rect 59 5493 65 5545
rect 1633 5493 1639 5545
rect 1691 5493 1697 5545
rect 3265 5493 3271 5545
rect 3323 5493 3329 5545
rect 4897 5493 4903 5545
rect 4955 5493 4961 5545
rect 6529 5493 6535 5545
rect 6587 5493 6593 5545
rect 8161 5493 8167 5545
rect 8219 5493 8225 5545
rect 9793 5493 9799 5545
rect 9851 5493 9857 5545
rect 8 5486 59 5493
rect 1640 5486 1691 5493
rect 3272 5486 3323 5493
rect 4904 5486 4955 5493
rect 6536 5486 6587 5493
rect 8168 5486 8219 5493
rect 9800 5486 9851 5493
rect 8 5341 59 5348
rect 1640 5341 1691 5348
rect 3272 5341 3323 5348
rect 4904 5341 4955 5348
rect 6536 5341 6587 5348
rect 8168 5341 8219 5348
rect 9800 5341 9851 5348
rect 1 5289 7 5341
rect 59 5289 65 5341
rect 1633 5289 1639 5341
rect 1691 5289 1697 5341
rect 3265 5289 3271 5341
rect 3323 5289 3329 5341
rect 4897 5289 4903 5341
rect 4955 5289 4961 5341
rect 6529 5289 6535 5341
rect 6587 5289 6593 5341
rect 8161 5289 8167 5341
rect 8219 5289 8225 5341
rect 9793 5289 9799 5341
rect 9851 5289 9857 5341
rect 8 5282 59 5289
rect 1640 5282 1691 5289
rect 3272 5282 3323 5289
rect 4904 5282 4955 5289
rect 6536 5282 6587 5289
rect 8168 5282 8219 5289
rect 9800 5282 9851 5289
rect 8 5137 59 5144
rect 1640 5137 1691 5144
rect 3272 5137 3323 5144
rect 4904 5137 4955 5144
rect 6536 5137 6587 5144
rect 8168 5137 8219 5144
rect 9800 5137 9851 5144
rect 1 5085 7 5137
rect 59 5085 65 5137
rect 1633 5085 1639 5137
rect 1691 5085 1697 5137
rect 3265 5085 3271 5137
rect 3323 5085 3329 5137
rect 4897 5085 4903 5137
rect 4955 5085 4961 5137
rect 6529 5085 6535 5137
rect 6587 5085 6593 5137
rect 8161 5085 8167 5137
rect 8219 5085 8225 5137
rect 9793 5085 9799 5137
rect 9851 5085 9857 5137
rect 8 5078 59 5085
rect 1640 5078 1691 5085
rect 3272 5078 3323 5085
rect 4904 5078 4955 5085
rect 6536 5078 6587 5085
rect 8168 5078 8219 5085
rect 9800 5078 9851 5085
rect 8 4933 59 4940
rect 1640 4933 1691 4940
rect 3272 4933 3323 4940
rect 4904 4933 4955 4940
rect 6536 4933 6587 4940
rect 8168 4933 8219 4940
rect 9800 4933 9851 4940
rect 1 4881 7 4933
rect 59 4881 65 4933
rect 1633 4881 1639 4933
rect 1691 4881 1697 4933
rect 3265 4881 3271 4933
rect 3323 4881 3329 4933
rect 4897 4881 4903 4933
rect 4955 4881 4961 4933
rect 6529 4881 6535 4933
rect 6587 4881 6593 4933
rect 8161 4881 8167 4933
rect 8219 4881 8225 4933
rect 9793 4881 9799 4933
rect 9851 4881 9857 4933
rect 8 4874 59 4881
rect 1640 4874 1691 4881
rect 3272 4874 3323 4881
rect 4904 4874 4955 4881
rect 6536 4874 6587 4881
rect 8168 4874 8219 4881
rect 9800 4874 9851 4881
rect 8 4729 59 4736
rect 1640 4729 1691 4736
rect 3272 4729 3323 4736
rect 4904 4729 4955 4736
rect 6536 4729 6587 4736
rect 8168 4729 8219 4736
rect 9800 4729 9851 4736
rect 1 4677 7 4729
rect 59 4677 65 4729
rect 1633 4677 1639 4729
rect 1691 4677 1697 4729
rect 3265 4677 3271 4729
rect 3323 4677 3329 4729
rect 4897 4677 4903 4729
rect 4955 4677 4961 4729
rect 6529 4677 6535 4729
rect 6587 4677 6593 4729
rect 8161 4677 8167 4729
rect 8219 4677 8225 4729
rect 9793 4677 9799 4729
rect 9851 4677 9857 4729
rect 8 4670 59 4677
rect 1640 4670 1691 4677
rect 3272 4670 3323 4677
rect 4904 4670 4955 4677
rect 6536 4670 6587 4677
rect 8168 4670 8219 4677
rect 9800 4670 9851 4677
rect 8 4525 59 4532
rect 1640 4525 1691 4532
rect 3272 4525 3323 4532
rect 4904 4525 4955 4532
rect 6536 4525 6587 4532
rect 8168 4525 8219 4532
rect 9800 4525 9851 4532
rect 1 4473 7 4525
rect 59 4473 65 4525
rect 1633 4473 1639 4525
rect 1691 4473 1697 4525
rect 3265 4473 3271 4525
rect 3323 4473 3329 4525
rect 4897 4473 4903 4525
rect 4955 4473 4961 4525
rect 6529 4473 6535 4525
rect 6587 4473 6593 4525
rect 8161 4473 8167 4525
rect 8219 4473 8225 4525
rect 9793 4473 9799 4525
rect 9851 4473 9857 4525
rect 8 4466 59 4473
rect 1640 4466 1691 4473
rect 3272 4466 3323 4473
rect 4904 4466 4955 4473
rect 6536 4466 6587 4473
rect 8168 4466 8219 4473
rect 9800 4466 9851 4473
rect 128 4241 156 4449
rect 218 4371 270 4377
rect 218 4313 270 4319
rect 332 4241 360 4449
rect 422 4371 474 4377
rect 422 4313 474 4319
rect 536 4241 564 4449
rect 626 4371 678 4377
rect 626 4313 678 4319
rect 740 4241 768 4449
rect 830 4371 882 4377
rect 830 4313 882 4319
rect 944 4241 972 4449
rect 1034 4371 1086 4377
rect 1034 4313 1086 4319
rect 1148 4241 1176 4449
rect 1238 4371 1290 4377
rect 1238 4313 1290 4319
rect 1352 4241 1380 4449
rect 1442 4371 1494 4377
rect 1442 4313 1494 4319
rect 1556 4241 1584 4449
rect 1646 4371 1698 4377
rect 1646 4313 1698 4319
rect 1760 4241 1788 4449
rect 1850 4371 1902 4377
rect 1850 4313 1902 4319
rect 1964 4241 1992 4449
rect 2054 4371 2106 4377
rect 2054 4313 2106 4319
rect 2168 4241 2196 4449
rect 2258 4371 2310 4377
rect 2258 4313 2310 4319
rect 2372 4241 2400 4449
rect 2462 4371 2514 4377
rect 2462 4313 2514 4319
rect 2576 4241 2604 4449
rect 2666 4371 2718 4377
rect 2666 4313 2718 4319
rect 2780 4241 2808 4449
rect 2870 4371 2922 4377
rect 2870 4313 2922 4319
rect 2984 4241 3012 4449
rect 3074 4371 3126 4377
rect 3074 4313 3126 4319
rect 3188 4241 3216 4449
rect 3278 4371 3330 4377
rect 3278 4313 3330 4319
rect 3392 4241 3420 4449
rect 3482 4371 3534 4377
rect 3482 4313 3534 4319
rect 3596 4241 3624 4449
rect 3686 4371 3738 4377
rect 3686 4313 3738 4319
rect 3800 4241 3828 4449
rect 3890 4371 3942 4377
rect 3890 4313 3942 4319
rect 4004 4241 4032 4449
rect 4094 4371 4146 4377
rect 4094 4313 4146 4319
rect 4208 4241 4236 4449
rect 4298 4371 4350 4377
rect 4298 4313 4350 4319
rect 4412 4241 4440 4449
rect 4502 4371 4554 4377
rect 4502 4313 4554 4319
rect 4616 4241 4644 4449
rect 4706 4371 4758 4377
rect 4706 4313 4758 4319
rect 4820 4241 4848 4449
rect 4910 4371 4962 4377
rect 4910 4313 4962 4319
rect 5024 4241 5052 4449
rect 5114 4371 5166 4377
rect 5114 4313 5166 4319
rect 5228 4241 5256 4449
rect 5318 4371 5370 4377
rect 5318 4313 5370 4319
rect 5432 4241 5460 4449
rect 5522 4371 5574 4377
rect 5522 4313 5574 4319
rect 5636 4241 5664 4449
rect 5726 4371 5778 4377
rect 5726 4313 5778 4319
rect 5840 4241 5868 4449
rect 5930 4371 5982 4377
rect 5930 4313 5982 4319
rect 6044 4241 6072 4449
rect 6134 4371 6186 4377
rect 6134 4313 6186 4319
rect 6248 4241 6276 4449
rect 6338 4371 6390 4377
rect 6338 4313 6390 4319
rect 6452 4241 6480 4449
rect 6542 4371 6594 4377
rect 6542 4313 6594 4319
rect 6656 4241 6684 4449
rect 6746 4371 6798 4377
rect 6746 4313 6798 4319
rect 6860 4241 6888 4449
rect 6950 4371 7002 4377
rect 6950 4313 7002 4319
rect 7064 4241 7092 4449
rect 7154 4371 7206 4377
rect 7154 4313 7206 4319
rect 7268 4241 7296 4449
rect 7358 4371 7410 4377
rect 7358 4313 7410 4319
rect 7472 4241 7500 4449
rect 7562 4371 7614 4377
rect 7562 4313 7614 4319
rect 7676 4241 7704 4449
rect 7766 4371 7818 4377
rect 7766 4313 7818 4319
rect 7880 4241 7908 4449
rect 7970 4371 8022 4377
rect 7970 4313 8022 4319
rect 8084 4241 8112 4449
rect 8174 4371 8226 4377
rect 8174 4313 8226 4319
rect 8288 4241 8316 4449
rect 8378 4371 8430 4377
rect 8378 4313 8430 4319
rect 8492 4241 8520 4449
rect 8582 4371 8634 4377
rect 8582 4313 8634 4319
rect 8696 4241 8724 4449
rect 8786 4371 8838 4377
rect 8786 4313 8838 4319
rect 8900 4241 8928 4449
rect 8990 4371 9042 4377
rect 8990 4313 9042 4319
rect 9104 4241 9132 4449
rect 9194 4371 9246 4377
rect 9194 4313 9246 4319
rect 9308 4241 9336 4449
rect 9398 4371 9450 4377
rect 9398 4313 9450 4319
rect 9512 4241 9540 4449
rect 9602 4371 9654 4377
rect 9602 4313 9654 4319
rect 9716 4241 9744 4449
rect 9820 4371 9872 4377
rect 9820 4313 9872 4319
rect 8 4217 59 4224
rect 1640 4217 1691 4224
rect 3272 4217 3323 4224
rect 4904 4217 4955 4224
rect 6536 4217 6587 4224
rect 8168 4217 8219 4224
rect 9800 4217 9851 4224
rect 1 4165 7 4217
rect 59 4165 65 4217
rect 1633 4165 1639 4217
rect 1691 4165 1697 4217
rect 3265 4165 3271 4217
rect 3323 4165 3329 4217
rect 4897 4165 4903 4217
rect 4955 4165 4961 4217
rect 6529 4165 6535 4217
rect 6587 4165 6593 4217
rect 8161 4165 8167 4217
rect 8219 4165 8225 4217
rect 9793 4165 9799 4217
rect 9851 4165 9857 4217
rect 8 4158 59 4165
rect 1640 4158 1691 4165
rect 3272 4158 3323 4165
rect 4904 4158 4955 4165
rect 6536 4158 6587 4165
rect 8168 4158 8219 4165
rect 9800 4158 9851 4165
rect 8 4013 59 4020
rect 1640 4013 1691 4020
rect 3272 4013 3323 4020
rect 4904 4013 4955 4020
rect 6536 4013 6587 4020
rect 8168 4013 8219 4020
rect 9800 4013 9851 4020
rect 1 3961 7 4013
rect 59 3961 65 4013
rect 1633 3961 1639 4013
rect 1691 3961 1697 4013
rect 3265 3961 3271 4013
rect 3323 3961 3329 4013
rect 4897 3961 4903 4013
rect 4955 3961 4961 4013
rect 6529 3961 6535 4013
rect 6587 3961 6593 4013
rect 8161 3961 8167 4013
rect 8219 3961 8225 4013
rect 9793 3961 9799 4013
rect 9851 3961 9857 4013
rect 8 3954 59 3961
rect 1640 3954 1691 3961
rect 3272 3954 3323 3961
rect 4904 3954 4955 3961
rect 6536 3954 6587 3961
rect 8168 3954 8219 3961
rect 9800 3954 9851 3961
rect 8 3809 59 3816
rect 1640 3809 1691 3816
rect 3272 3809 3323 3816
rect 4904 3809 4955 3816
rect 6536 3809 6587 3816
rect 8168 3809 8219 3816
rect 9800 3809 9851 3816
rect 1 3757 7 3809
rect 59 3757 65 3809
rect 1633 3757 1639 3809
rect 1691 3757 1697 3809
rect 3265 3757 3271 3809
rect 3323 3757 3329 3809
rect 4897 3757 4903 3809
rect 4955 3757 4961 3809
rect 6529 3757 6535 3809
rect 6587 3757 6593 3809
rect 8161 3757 8167 3809
rect 8219 3757 8225 3809
rect 9793 3757 9799 3809
rect 9851 3757 9857 3809
rect 8 3750 59 3757
rect 1640 3750 1691 3757
rect 3272 3750 3323 3757
rect 4904 3750 4955 3757
rect 6536 3750 6587 3757
rect 8168 3750 8219 3757
rect 9800 3750 9851 3757
rect 8 3605 59 3612
rect 1640 3605 1691 3612
rect 3272 3605 3323 3612
rect 4904 3605 4955 3612
rect 6536 3605 6587 3612
rect 8168 3605 8219 3612
rect 9800 3605 9851 3612
rect 1 3553 7 3605
rect 59 3553 65 3605
rect 1633 3553 1639 3605
rect 1691 3553 1697 3605
rect 3265 3553 3271 3605
rect 3323 3553 3329 3605
rect 4897 3553 4903 3605
rect 4955 3553 4961 3605
rect 6529 3553 6535 3605
rect 6587 3553 6593 3605
rect 8161 3553 8167 3605
rect 8219 3553 8225 3605
rect 9793 3553 9799 3605
rect 9851 3553 9857 3605
rect 8 3546 59 3553
rect 1640 3546 1691 3553
rect 3272 3546 3323 3553
rect 4904 3546 4955 3553
rect 6536 3546 6587 3553
rect 8168 3546 8219 3553
rect 9800 3546 9851 3553
rect 8 3401 59 3408
rect 1640 3401 1691 3408
rect 3272 3401 3323 3408
rect 4904 3401 4955 3408
rect 6536 3401 6587 3408
rect 8168 3401 8219 3408
rect 9800 3401 9851 3408
rect 1 3349 7 3401
rect 59 3349 65 3401
rect 1633 3349 1639 3401
rect 1691 3349 1697 3401
rect 3265 3349 3271 3401
rect 3323 3349 3329 3401
rect 4897 3349 4903 3401
rect 4955 3349 4961 3401
rect 6529 3349 6535 3401
rect 6587 3349 6593 3401
rect 8161 3349 8167 3401
rect 8219 3349 8225 3401
rect 9793 3349 9799 3401
rect 9851 3349 9857 3401
rect 8 3342 59 3349
rect 1640 3342 1691 3349
rect 3272 3342 3323 3349
rect 4904 3342 4955 3349
rect 6536 3342 6587 3349
rect 8168 3342 8219 3349
rect 9800 3342 9851 3349
rect 8 3197 59 3204
rect 1640 3197 1691 3204
rect 3272 3197 3323 3204
rect 4904 3197 4955 3204
rect 6536 3197 6587 3204
rect 8168 3197 8219 3204
rect 9800 3197 9851 3204
rect 1 3145 7 3197
rect 59 3145 65 3197
rect 1633 3145 1639 3197
rect 1691 3145 1697 3197
rect 3265 3145 3271 3197
rect 3323 3145 3329 3197
rect 4897 3145 4903 3197
rect 4955 3145 4961 3197
rect 6529 3145 6535 3197
rect 6587 3145 6593 3197
rect 8161 3145 8167 3197
rect 8219 3145 8225 3197
rect 9793 3145 9799 3197
rect 9851 3145 9857 3197
rect 8 3138 59 3145
rect 1640 3138 1691 3145
rect 3272 3138 3323 3145
rect 4904 3138 4955 3145
rect 6536 3138 6587 3145
rect 8168 3138 8219 3145
rect 9800 3138 9851 3145
rect 8 2993 59 3000
rect 1640 2993 1691 3000
rect 3272 2993 3323 3000
rect 4904 2993 4955 3000
rect 6536 2993 6587 3000
rect 8168 2993 8219 3000
rect 9800 2993 9851 3000
rect 1 2941 7 2993
rect 59 2941 65 2993
rect 1633 2941 1639 2993
rect 1691 2941 1697 2993
rect 3265 2941 3271 2993
rect 3323 2941 3329 2993
rect 4897 2941 4903 2993
rect 4955 2941 4961 2993
rect 6529 2941 6535 2993
rect 6587 2941 6593 2993
rect 8161 2941 8167 2993
rect 8219 2941 8225 2993
rect 9793 2941 9799 2993
rect 9851 2941 9857 2993
rect 8 2934 59 2941
rect 1640 2934 1691 2941
rect 3272 2934 3323 2941
rect 4904 2934 4955 2941
rect 6536 2934 6587 2941
rect 8168 2934 8219 2941
rect 9800 2934 9851 2941
rect 8 2789 59 2796
rect 1640 2789 1691 2796
rect 3272 2789 3323 2796
rect 4904 2789 4955 2796
rect 6536 2789 6587 2796
rect 8168 2789 8219 2796
rect 9800 2789 9851 2796
rect 1 2737 7 2789
rect 59 2737 65 2789
rect 1633 2737 1639 2789
rect 1691 2737 1697 2789
rect 3265 2737 3271 2789
rect 3323 2737 3329 2789
rect 4897 2737 4903 2789
rect 4955 2737 4961 2789
rect 6529 2737 6535 2789
rect 6587 2737 6593 2789
rect 8161 2737 8167 2789
rect 8219 2737 8225 2789
rect 9793 2737 9799 2789
rect 9851 2737 9857 2789
rect 8 2730 59 2737
rect 1640 2730 1691 2737
rect 3272 2730 3323 2737
rect 4904 2730 4955 2737
rect 6536 2730 6587 2737
rect 8168 2730 8219 2737
rect 9800 2730 9851 2737
rect 128 2505 156 2713
rect 218 2635 270 2641
rect 218 2577 270 2583
rect 332 2505 360 2713
rect 422 2635 474 2641
rect 422 2577 474 2583
rect 536 2505 564 2713
rect 626 2635 678 2641
rect 626 2577 678 2583
rect 740 2505 768 2713
rect 830 2635 882 2641
rect 830 2577 882 2583
rect 944 2505 972 2713
rect 1034 2635 1086 2641
rect 1034 2577 1086 2583
rect 1148 2505 1176 2713
rect 1238 2635 1290 2641
rect 1238 2577 1290 2583
rect 1352 2505 1380 2713
rect 1442 2635 1494 2641
rect 1442 2577 1494 2583
rect 1556 2505 1584 2713
rect 1646 2635 1698 2641
rect 1646 2577 1698 2583
rect 1760 2505 1788 2713
rect 1850 2635 1902 2641
rect 1850 2577 1902 2583
rect 1964 2505 1992 2713
rect 2054 2635 2106 2641
rect 2054 2577 2106 2583
rect 2168 2505 2196 2713
rect 2258 2635 2310 2641
rect 2258 2577 2310 2583
rect 2372 2505 2400 2713
rect 2462 2635 2514 2641
rect 2462 2577 2514 2583
rect 2576 2505 2604 2713
rect 2666 2635 2718 2641
rect 2666 2577 2718 2583
rect 2780 2505 2808 2713
rect 2870 2635 2922 2641
rect 2870 2577 2922 2583
rect 2984 2505 3012 2713
rect 3074 2635 3126 2641
rect 3074 2577 3126 2583
rect 3188 2505 3216 2713
rect 3278 2635 3330 2641
rect 3278 2577 3330 2583
rect 3392 2505 3420 2713
rect 3482 2635 3534 2641
rect 3482 2577 3534 2583
rect 3596 2505 3624 2713
rect 3686 2635 3738 2641
rect 3686 2577 3738 2583
rect 3800 2505 3828 2713
rect 3890 2635 3942 2641
rect 3890 2577 3942 2583
rect 4004 2505 4032 2713
rect 4094 2635 4146 2641
rect 4094 2577 4146 2583
rect 4208 2505 4236 2713
rect 4298 2635 4350 2641
rect 4298 2577 4350 2583
rect 4412 2505 4440 2713
rect 4502 2635 4554 2641
rect 4502 2577 4554 2583
rect 4616 2505 4644 2713
rect 4706 2635 4758 2641
rect 4706 2577 4758 2583
rect 4820 2505 4848 2713
rect 4910 2635 4962 2641
rect 4910 2577 4962 2583
rect 5024 2505 5052 2713
rect 5114 2635 5166 2641
rect 5114 2577 5166 2583
rect 5228 2505 5256 2713
rect 5318 2635 5370 2641
rect 5318 2577 5370 2583
rect 5432 2505 5460 2713
rect 5522 2635 5574 2641
rect 5522 2577 5574 2583
rect 5636 2505 5664 2713
rect 5726 2635 5778 2641
rect 5726 2577 5778 2583
rect 5840 2505 5868 2713
rect 5930 2635 5982 2641
rect 5930 2577 5982 2583
rect 6044 2505 6072 2713
rect 6134 2635 6186 2641
rect 6134 2577 6186 2583
rect 6248 2505 6276 2713
rect 6338 2635 6390 2641
rect 6338 2577 6390 2583
rect 6452 2505 6480 2713
rect 6542 2635 6594 2641
rect 6542 2577 6594 2583
rect 6656 2505 6684 2713
rect 6746 2635 6798 2641
rect 6746 2577 6798 2583
rect 6860 2505 6888 2713
rect 6950 2635 7002 2641
rect 6950 2577 7002 2583
rect 7064 2505 7092 2713
rect 7154 2635 7206 2641
rect 7154 2577 7206 2583
rect 7268 2505 7296 2713
rect 7358 2635 7410 2641
rect 7358 2577 7410 2583
rect 7472 2505 7500 2713
rect 7562 2635 7614 2641
rect 7562 2577 7614 2583
rect 7676 2505 7704 2713
rect 7766 2635 7818 2641
rect 7766 2577 7818 2583
rect 7880 2505 7908 2713
rect 7970 2635 8022 2641
rect 7970 2577 8022 2583
rect 8084 2505 8112 2713
rect 8174 2635 8226 2641
rect 8174 2577 8226 2583
rect 8288 2505 8316 2713
rect 8378 2635 8430 2641
rect 8378 2577 8430 2583
rect 8492 2505 8520 2713
rect 8582 2635 8634 2641
rect 8582 2577 8634 2583
rect 8696 2505 8724 2713
rect 8786 2635 8838 2641
rect 8786 2577 8838 2583
rect 8900 2505 8928 2713
rect 8990 2635 9042 2641
rect 8990 2577 9042 2583
rect 9104 2505 9132 2713
rect 9194 2635 9246 2641
rect 9194 2577 9246 2583
rect 9308 2505 9336 2713
rect 9398 2635 9450 2641
rect 9398 2577 9450 2583
rect 9512 2505 9540 2713
rect 9602 2635 9654 2641
rect 9602 2577 9654 2583
rect 9716 2505 9744 2713
rect 9820 2635 9872 2641
rect 9820 2577 9872 2583
rect 8 2481 59 2488
rect 1640 2481 1691 2488
rect 3272 2481 3323 2488
rect 4904 2481 4955 2488
rect 6536 2481 6587 2488
rect 8168 2481 8219 2488
rect 9800 2481 9851 2488
rect 1 2429 7 2481
rect 59 2429 65 2481
rect 1633 2429 1639 2481
rect 1691 2429 1697 2481
rect 3265 2429 3271 2481
rect 3323 2429 3329 2481
rect 4897 2429 4903 2481
rect 4955 2429 4961 2481
rect 6529 2429 6535 2481
rect 6587 2429 6593 2481
rect 8161 2429 8167 2481
rect 8219 2429 8225 2481
rect 9793 2429 9799 2481
rect 9851 2429 9857 2481
rect 8 2422 59 2429
rect 1640 2422 1691 2429
rect 3272 2422 3323 2429
rect 4904 2422 4955 2429
rect 6536 2422 6587 2429
rect 8168 2422 8219 2429
rect 9800 2422 9851 2429
rect 8 2277 59 2284
rect 1640 2277 1691 2284
rect 3272 2277 3323 2284
rect 4904 2277 4955 2284
rect 6536 2277 6587 2284
rect 8168 2277 8219 2284
rect 9800 2277 9851 2284
rect 1 2225 7 2277
rect 59 2225 65 2277
rect 1633 2225 1639 2277
rect 1691 2225 1697 2277
rect 3265 2225 3271 2277
rect 3323 2225 3329 2277
rect 4897 2225 4903 2277
rect 4955 2225 4961 2277
rect 6529 2225 6535 2277
rect 6587 2225 6593 2277
rect 8161 2225 8167 2277
rect 8219 2225 8225 2277
rect 9793 2225 9799 2277
rect 9851 2225 9857 2277
rect 8 2218 59 2225
rect 1640 2218 1691 2225
rect 3272 2218 3323 2225
rect 4904 2218 4955 2225
rect 6536 2218 6587 2225
rect 8168 2218 8219 2225
rect 9800 2218 9851 2225
rect 8 2073 59 2080
rect 1640 2073 1691 2080
rect 3272 2073 3323 2080
rect 4904 2073 4955 2080
rect 6536 2073 6587 2080
rect 8168 2073 8219 2080
rect 9800 2073 9851 2080
rect 1 2021 7 2073
rect 59 2021 65 2073
rect 1633 2021 1639 2073
rect 1691 2021 1697 2073
rect 3265 2021 3271 2073
rect 3323 2021 3329 2073
rect 4897 2021 4903 2073
rect 4955 2021 4961 2073
rect 6529 2021 6535 2073
rect 6587 2021 6593 2073
rect 8161 2021 8167 2073
rect 8219 2021 8225 2073
rect 9793 2021 9799 2073
rect 9851 2021 9857 2073
rect 8 2014 59 2021
rect 1640 2014 1691 2021
rect 3272 2014 3323 2021
rect 4904 2014 4955 2021
rect 6536 2014 6587 2021
rect 8168 2014 8219 2021
rect 9800 2014 9851 2021
rect 8 1869 59 1876
rect 1640 1869 1691 1876
rect 3272 1869 3323 1876
rect 4904 1869 4955 1876
rect 6536 1869 6587 1876
rect 8168 1869 8219 1876
rect 9800 1869 9851 1876
rect 1 1817 7 1869
rect 59 1817 65 1869
rect 1633 1817 1639 1869
rect 1691 1817 1697 1869
rect 3265 1817 3271 1869
rect 3323 1817 3329 1869
rect 4897 1817 4903 1869
rect 4955 1817 4961 1869
rect 6529 1817 6535 1869
rect 6587 1817 6593 1869
rect 8161 1817 8167 1869
rect 8219 1817 8225 1869
rect 9793 1817 9799 1869
rect 9851 1817 9857 1869
rect 8 1810 59 1817
rect 1640 1810 1691 1817
rect 3272 1810 3323 1817
rect 4904 1810 4955 1817
rect 6536 1810 6587 1817
rect 8168 1810 8219 1817
rect 9800 1810 9851 1817
rect 8 1665 59 1672
rect 1640 1665 1691 1672
rect 3272 1665 3323 1672
rect 4904 1665 4955 1672
rect 6536 1665 6587 1672
rect 8168 1665 8219 1672
rect 9800 1665 9851 1672
rect 1 1613 7 1665
rect 59 1613 65 1665
rect 1633 1613 1639 1665
rect 1691 1613 1697 1665
rect 3265 1613 3271 1665
rect 3323 1613 3329 1665
rect 4897 1613 4903 1665
rect 4955 1613 4961 1665
rect 6529 1613 6535 1665
rect 6587 1613 6593 1665
rect 8161 1613 8167 1665
rect 8219 1613 8225 1665
rect 9793 1613 9799 1665
rect 9851 1613 9857 1665
rect 8 1606 59 1613
rect 1640 1606 1691 1613
rect 3272 1606 3323 1613
rect 4904 1606 4955 1613
rect 6536 1606 6587 1613
rect 8168 1606 8219 1613
rect 9800 1606 9851 1613
rect 8 1461 59 1468
rect 1640 1461 1691 1468
rect 3272 1461 3323 1468
rect 4904 1461 4955 1468
rect 6536 1461 6587 1468
rect 8168 1461 8219 1468
rect 9800 1461 9851 1468
rect 1 1409 7 1461
rect 59 1409 65 1461
rect 1633 1409 1639 1461
rect 1691 1409 1697 1461
rect 3265 1409 3271 1461
rect 3323 1409 3329 1461
rect 4897 1409 4903 1461
rect 4955 1409 4961 1461
rect 6529 1409 6535 1461
rect 6587 1409 6593 1461
rect 8161 1409 8167 1461
rect 8219 1409 8225 1461
rect 9793 1409 9799 1461
rect 9851 1409 9857 1461
rect 8 1402 59 1409
rect 1640 1402 1691 1409
rect 3272 1402 3323 1409
rect 4904 1402 4955 1409
rect 6536 1402 6587 1409
rect 8168 1402 8219 1409
rect 9800 1402 9851 1409
rect 8 1257 59 1264
rect 1640 1257 1691 1264
rect 3272 1257 3323 1264
rect 4904 1257 4955 1264
rect 6536 1257 6587 1264
rect 8168 1257 8219 1264
rect 9800 1257 9851 1264
rect 1 1205 7 1257
rect 59 1205 65 1257
rect 1633 1205 1639 1257
rect 1691 1205 1697 1257
rect 3265 1205 3271 1257
rect 3323 1205 3329 1257
rect 4897 1205 4903 1257
rect 4955 1205 4961 1257
rect 6529 1205 6535 1257
rect 6587 1205 6593 1257
rect 8161 1205 8167 1257
rect 8219 1205 8225 1257
rect 9793 1205 9799 1257
rect 9851 1205 9857 1257
rect 8 1198 59 1205
rect 1640 1198 1691 1205
rect 3272 1198 3323 1205
rect 4904 1198 4955 1205
rect 6536 1198 6587 1205
rect 8168 1198 8219 1205
rect 9800 1198 9851 1205
rect 8 1053 59 1060
rect 1640 1053 1691 1060
rect 3272 1053 3323 1060
rect 4904 1053 4955 1060
rect 6536 1053 6587 1060
rect 8168 1053 8219 1060
rect 9800 1053 9851 1060
rect 1 1001 7 1053
rect 59 1001 65 1053
rect 1633 1001 1639 1053
rect 1691 1001 1697 1053
rect 3265 1001 3271 1053
rect 3323 1001 3329 1053
rect 4897 1001 4903 1053
rect 4955 1001 4961 1053
rect 6529 1001 6535 1053
rect 6587 1001 6593 1053
rect 8161 1001 8167 1053
rect 8219 1001 8225 1053
rect 9793 1001 9799 1053
rect 9851 1001 9857 1053
rect 8 994 59 1001
rect 1640 994 1691 1001
rect 3272 994 3323 1001
rect 4904 994 4955 1001
rect 6536 994 6587 1001
rect 8168 994 8219 1001
rect 9800 994 9851 1001
rect 128 -14 156 977
rect 218 899 270 905
rect 218 841 270 847
rect 332 -14 360 977
rect 422 899 474 905
rect 422 841 474 847
rect 536 -14 564 977
rect 626 899 678 905
rect 626 841 678 847
rect 740 -14 768 977
rect 830 899 882 905
rect 830 841 882 847
rect 944 -14 972 977
rect 1034 899 1086 905
rect 1034 841 1086 847
rect 1148 -14 1176 977
rect 1238 899 1290 905
rect 1238 841 1290 847
rect 1352 -14 1380 977
rect 1442 899 1494 905
rect 1442 841 1494 847
rect 1556 -14 1584 977
rect 1646 899 1698 905
rect 1646 841 1698 847
rect 1760 -14 1788 977
rect 1850 899 1902 905
rect 1850 841 1902 847
rect 1964 -14 1992 977
rect 2054 899 2106 905
rect 2054 841 2106 847
rect 2168 -14 2196 977
rect 2258 899 2310 905
rect 2258 841 2310 847
rect 2372 -14 2400 977
rect 2462 899 2514 905
rect 2462 841 2514 847
rect 2576 -14 2604 977
rect 2666 899 2718 905
rect 2666 841 2718 847
rect 2780 -14 2808 977
rect 2870 899 2922 905
rect 2870 841 2922 847
rect 2984 -14 3012 977
rect 3074 899 3126 905
rect 3074 841 3126 847
rect 3188 -14 3216 977
rect 3278 899 3330 905
rect 3278 841 3330 847
rect 3392 -14 3420 977
rect 3482 899 3534 905
rect 3482 841 3534 847
rect 3596 -14 3624 977
rect 3686 899 3738 905
rect 3686 841 3738 847
rect 3800 -14 3828 977
rect 3890 899 3942 905
rect 3890 841 3942 847
rect 4004 -14 4032 977
rect 4094 899 4146 905
rect 4094 841 4146 847
rect 4208 -14 4236 977
rect 4298 899 4350 905
rect 4298 841 4350 847
rect 4412 -14 4440 977
rect 4502 899 4554 905
rect 4502 841 4554 847
rect 4616 -14 4644 977
rect 4706 899 4758 905
rect 4706 841 4758 847
rect 4820 -14 4848 977
rect 4910 899 4962 905
rect 4910 841 4962 847
rect 5024 -14 5052 977
rect 5114 899 5166 905
rect 5114 841 5166 847
rect 5228 -14 5256 977
rect 5318 899 5370 905
rect 5318 841 5370 847
rect 5432 -14 5460 977
rect 5522 899 5574 905
rect 5522 841 5574 847
rect 5636 -14 5664 977
rect 5726 899 5778 905
rect 5726 841 5778 847
rect 5840 -14 5868 977
rect 5930 899 5982 905
rect 5930 841 5982 847
rect 6044 -14 6072 977
rect 6134 899 6186 905
rect 6134 841 6186 847
rect 6248 -14 6276 977
rect 6338 899 6390 905
rect 6338 841 6390 847
rect 6452 -14 6480 977
rect 6542 899 6594 905
rect 6542 841 6594 847
rect 6656 -14 6684 977
rect 6746 899 6798 905
rect 6746 841 6798 847
rect 6860 -14 6888 977
rect 6950 899 7002 905
rect 6950 841 7002 847
rect 7064 -14 7092 977
rect 7154 899 7206 905
rect 7154 841 7206 847
rect 7268 -14 7296 977
rect 7358 899 7410 905
rect 7358 841 7410 847
rect 7472 -14 7500 977
rect 7562 899 7614 905
rect 7562 841 7614 847
rect 7676 -14 7704 977
rect 7766 899 7818 905
rect 7766 841 7818 847
rect 7880 -14 7908 977
rect 7970 899 8022 905
rect 7970 841 8022 847
rect 8084 -14 8112 977
rect 8174 899 8226 905
rect 8174 841 8226 847
rect 8288 -14 8316 977
rect 8378 899 8430 905
rect 8378 841 8430 847
rect 8492 -14 8520 977
rect 8582 899 8634 905
rect 8582 841 8634 847
rect 8696 -14 8724 977
rect 8786 899 8838 905
rect 8786 841 8838 847
rect 8900 -14 8928 977
rect 8990 899 9042 905
rect 8990 841 9042 847
rect 9104 -14 9132 977
rect 9194 899 9246 905
rect 9194 841 9246 847
rect 9308 -14 9336 977
rect 9398 899 9450 905
rect 9398 841 9450 847
rect 9512 -14 9540 977
rect 9602 899 9654 905
rect 9602 841 9654 847
rect 9716 -14 9744 977
rect 9820 899 9872 905
rect 9820 841 9872 847
rect 10013 396 10041 10101
rect 9867 368 10041 396
<< via1 >>
rect 7 10132 59 10141
rect 7 10098 16 10132
rect 16 10098 50 10132
rect 50 10098 59 10132
rect 7 10089 59 10098
rect 1639 10132 1691 10141
rect 1639 10098 1648 10132
rect 1648 10098 1682 10132
rect 1682 10098 1691 10132
rect 1639 10089 1691 10098
rect 3271 10132 3323 10141
rect 3271 10098 3280 10132
rect 3280 10098 3314 10132
rect 3314 10098 3323 10132
rect 3271 10089 3323 10098
rect 4903 10132 4955 10141
rect 4903 10098 4912 10132
rect 4912 10098 4946 10132
rect 4946 10098 4955 10132
rect 4903 10089 4955 10098
rect 6535 10132 6587 10141
rect 6535 10098 6544 10132
rect 6544 10098 6578 10132
rect 6578 10098 6587 10132
rect 6535 10089 6587 10098
rect 8167 10132 8219 10141
rect 8167 10098 8176 10132
rect 8176 10098 8210 10132
rect 8210 10098 8219 10132
rect 8167 10089 8219 10098
rect 9799 10132 9851 10141
rect 9799 10098 9808 10132
rect 9808 10098 9842 10132
rect 9842 10098 9851 10132
rect 9799 10089 9851 10098
rect 7 9928 59 9937
rect 7 9894 16 9928
rect 16 9894 50 9928
rect 50 9894 59 9928
rect 7 9885 59 9894
rect 1639 9928 1691 9937
rect 1639 9894 1648 9928
rect 1648 9894 1682 9928
rect 1682 9894 1691 9928
rect 1639 9885 1691 9894
rect 3271 9928 3323 9937
rect 3271 9894 3280 9928
rect 3280 9894 3314 9928
rect 3314 9894 3323 9928
rect 3271 9885 3323 9894
rect 4903 9928 4955 9937
rect 4903 9894 4912 9928
rect 4912 9894 4946 9928
rect 4946 9894 4955 9928
rect 4903 9885 4955 9894
rect 6535 9928 6587 9937
rect 6535 9894 6544 9928
rect 6544 9894 6578 9928
rect 6578 9894 6587 9928
rect 6535 9885 6587 9894
rect 8167 9928 8219 9937
rect 8167 9894 8176 9928
rect 8176 9894 8210 9928
rect 8210 9894 8219 9928
rect 8167 9885 8219 9894
rect 9799 9928 9851 9937
rect 9799 9894 9808 9928
rect 9808 9894 9842 9928
rect 9842 9894 9851 9928
rect 9799 9885 9851 9894
rect 7 9724 59 9733
rect 7 9690 16 9724
rect 16 9690 50 9724
rect 50 9690 59 9724
rect 7 9681 59 9690
rect 1639 9724 1691 9733
rect 1639 9690 1648 9724
rect 1648 9690 1682 9724
rect 1682 9690 1691 9724
rect 1639 9681 1691 9690
rect 3271 9724 3323 9733
rect 3271 9690 3280 9724
rect 3280 9690 3314 9724
rect 3314 9690 3323 9724
rect 3271 9681 3323 9690
rect 4903 9724 4955 9733
rect 4903 9690 4912 9724
rect 4912 9690 4946 9724
rect 4946 9690 4955 9724
rect 4903 9681 4955 9690
rect 6535 9724 6587 9733
rect 6535 9690 6544 9724
rect 6544 9690 6578 9724
rect 6578 9690 6587 9724
rect 6535 9681 6587 9690
rect 8167 9724 8219 9733
rect 8167 9690 8176 9724
rect 8176 9690 8210 9724
rect 8210 9690 8219 9724
rect 8167 9681 8219 9690
rect 9799 9724 9851 9733
rect 9799 9690 9808 9724
rect 9808 9690 9842 9724
rect 9842 9690 9851 9724
rect 9799 9681 9851 9690
rect 218 9570 270 9579
rect 218 9536 227 9570
rect 227 9536 261 9570
rect 261 9536 270 9570
rect 218 9527 270 9536
rect 422 9570 474 9579
rect 422 9536 431 9570
rect 431 9536 465 9570
rect 465 9536 474 9570
rect 422 9527 474 9536
rect 626 9570 678 9579
rect 626 9536 635 9570
rect 635 9536 669 9570
rect 669 9536 678 9570
rect 626 9527 678 9536
rect 830 9570 882 9579
rect 830 9536 839 9570
rect 839 9536 873 9570
rect 873 9536 882 9570
rect 830 9527 882 9536
rect 1034 9570 1086 9579
rect 1034 9536 1043 9570
rect 1043 9536 1077 9570
rect 1077 9536 1086 9570
rect 1034 9527 1086 9536
rect 1238 9570 1290 9579
rect 1238 9536 1247 9570
rect 1247 9536 1281 9570
rect 1281 9536 1290 9570
rect 1238 9527 1290 9536
rect 1442 9570 1494 9579
rect 1442 9536 1451 9570
rect 1451 9536 1485 9570
rect 1485 9536 1494 9570
rect 1442 9527 1494 9536
rect 1646 9570 1698 9579
rect 1646 9536 1655 9570
rect 1655 9536 1689 9570
rect 1689 9536 1698 9570
rect 1646 9527 1698 9536
rect 1850 9570 1902 9579
rect 1850 9536 1859 9570
rect 1859 9536 1893 9570
rect 1893 9536 1902 9570
rect 1850 9527 1902 9536
rect 2054 9570 2106 9579
rect 2054 9536 2063 9570
rect 2063 9536 2097 9570
rect 2097 9536 2106 9570
rect 2054 9527 2106 9536
rect 2258 9570 2310 9579
rect 2258 9536 2267 9570
rect 2267 9536 2301 9570
rect 2301 9536 2310 9570
rect 2258 9527 2310 9536
rect 2462 9570 2514 9579
rect 2462 9536 2471 9570
rect 2471 9536 2505 9570
rect 2505 9536 2514 9570
rect 2462 9527 2514 9536
rect 2666 9570 2718 9579
rect 2666 9536 2675 9570
rect 2675 9536 2709 9570
rect 2709 9536 2718 9570
rect 2666 9527 2718 9536
rect 2870 9570 2922 9579
rect 2870 9536 2879 9570
rect 2879 9536 2913 9570
rect 2913 9536 2922 9570
rect 2870 9527 2922 9536
rect 3074 9570 3126 9579
rect 3074 9536 3083 9570
rect 3083 9536 3117 9570
rect 3117 9536 3126 9570
rect 3074 9527 3126 9536
rect 3278 9570 3330 9579
rect 3278 9536 3287 9570
rect 3287 9536 3321 9570
rect 3321 9536 3330 9570
rect 3278 9527 3330 9536
rect 3482 9570 3534 9579
rect 3482 9536 3491 9570
rect 3491 9536 3525 9570
rect 3525 9536 3534 9570
rect 3482 9527 3534 9536
rect 3686 9570 3738 9579
rect 3686 9536 3695 9570
rect 3695 9536 3729 9570
rect 3729 9536 3738 9570
rect 3686 9527 3738 9536
rect 3890 9570 3942 9579
rect 3890 9536 3899 9570
rect 3899 9536 3933 9570
rect 3933 9536 3942 9570
rect 3890 9527 3942 9536
rect 4094 9570 4146 9579
rect 4094 9536 4103 9570
rect 4103 9536 4137 9570
rect 4137 9536 4146 9570
rect 4094 9527 4146 9536
rect 4298 9570 4350 9579
rect 4298 9536 4307 9570
rect 4307 9536 4341 9570
rect 4341 9536 4350 9570
rect 4298 9527 4350 9536
rect 4502 9570 4554 9579
rect 4502 9536 4511 9570
rect 4511 9536 4545 9570
rect 4545 9536 4554 9570
rect 4502 9527 4554 9536
rect 4706 9570 4758 9579
rect 4706 9536 4715 9570
rect 4715 9536 4749 9570
rect 4749 9536 4758 9570
rect 4706 9527 4758 9536
rect 4910 9570 4962 9579
rect 4910 9536 4919 9570
rect 4919 9536 4953 9570
rect 4953 9536 4962 9570
rect 4910 9527 4962 9536
rect 5114 9570 5166 9579
rect 5114 9536 5123 9570
rect 5123 9536 5157 9570
rect 5157 9536 5166 9570
rect 5114 9527 5166 9536
rect 5318 9570 5370 9579
rect 5318 9536 5327 9570
rect 5327 9536 5361 9570
rect 5361 9536 5370 9570
rect 5318 9527 5370 9536
rect 5522 9570 5574 9579
rect 5522 9536 5531 9570
rect 5531 9536 5565 9570
rect 5565 9536 5574 9570
rect 5522 9527 5574 9536
rect 5726 9570 5778 9579
rect 5726 9536 5735 9570
rect 5735 9536 5769 9570
rect 5769 9536 5778 9570
rect 5726 9527 5778 9536
rect 5930 9570 5982 9579
rect 5930 9536 5939 9570
rect 5939 9536 5973 9570
rect 5973 9536 5982 9570
rect 5930 9527 5982 9536
rect 6134 9570 6186 9579
rect 6134 9536 6143 9570
rect 6143 9536 6177 9570
rect 6177 9536 6186 9570
rect 6134 9527 6186 9536
rect 6338 9570 6390 9579
rect 6338 9536 6347 9570
rect 6347 9536 6381 9570
rect 6381 9536 6390 9570
rect 6338 9527 6390 9536
rect 6542 9570 6594 9579
rect 6542 9536 6551 9570
rect 6551 9536 6585 9570
rect 6585 9536 6594 9570
rect 6542 9527 6594 9536
rect 6746 9570 6798 9579
rect 6746 9536 6755 9570
rect 6755 9536 6789 9570
rect 6789 9536 6798 9570
rect 6746 9527 6798 9536
rect 6950 9570 7002 9579
rect 6950 9536 6959 9570
rect 6959 9536 6993 9570
rect 6993 9536 7002 9570
rect 6950 9527 7002 9536
rect 7154 9570 7206 9579
rect 7154 9536 7163 9570
rect 7163 9536 7197 9570
rect 7197 9536 7206 9570
rect 7154 9527 7206 9536
rect 7358 9570 7410 9579
rect 7358 9536 7367 9570
rect 7367 9536 7401 9570
rect 7401 9536 7410 9570
rect 7358 9527 7410 9536
rect 7562 9570 7614 9579
rect 7562 9536 7571 9570
rect 7571 9536 7605 9570
rect 7605 9536 7614 9570
rect 7562 9527 7614 9536
rect 7766 9570 7818 9579
rect 7766 9536 7775 9570
rect 7775 9536 7809 9570
rect 7809 9536 7818 9570
rect 7766 9527 7818 9536
rect 7970 9570 8022 9579
rect 7970 9536 7979 9570
rect 7979 9536 8013 9570
rect 8013 9536 8022 9570
rect 7970 9527 8022 9536
rect 8174 9570 8226 9579
rect 8174 9536 8183 9570
rect 8183 9536 8217 9570
rect 8217 9536 8226 9570
rect 8174 9527 8226 9536
rect 8378 9570 8430 9579
rect 8378 9536 8387 9570
rect 8387 9536 8421 9570
rect 8421 9536 8430 9570
rect 8378 9527 8430 9536
rect 8582 9570 8634 9579
rect 8582 9536 8591 9570
rect 8591 9536 8625 9570
rect 8625 9536 8634 9570
rect 8582 9527 8634 9536
rect 8786 9570 8838 9579
rect 8786 9536 8795 9570
rect 8795 9536 8829 9570
rect 8829 9536 8838 9570
rect 8786 9527 8838 9536
rect 8990 9570 9042 9579
rect 8990 9536 8999 9570
rect 8999 9536 9033 9570
rect 9033 9536 9042 9570
rect 8990 9527 9042 9536
rect 9194 9570 9246 9579
rect 9194 9536 9203 9570
rect 9203 9536 9237 9570
rect 9237 9536 9246 9570
rect 9194 9527 9246 9536
rect 9398 9570 9450 9579
rect 9398 9536 9407 9570
rect 9407 9536 9441 9570
rect 9441 9536 9450 9570
rect 9398 9527 9450 9536
rect 9602 9570 9654 9579
rect 9602 9536 9611 9570
rect 9611 9536 9645 9570
rect 9645 9536 9654 9570
rect 9602 9527 9654 9536
rect 9820 9570 9872 9579
rect 9820 9536 9829 9570
rect 9829 9536 9863 9570
rect 9863 9536 9872 9570
rect 9820 9527 9872 9536
rect 7 9416 59 9425
rect 7 9382 16 9416
rect 16 9382 50 9416
rect 50 9382 59 9416
rect 7 9373 59 9382
rect 1639 9416 1691 9425
rect 1639 9382 1648 9416
rect 1648 9382 1682 9416
rect 1682 9382 1691 9416
rect 1639 9373 1691 9382
rect 3271 9416 3323 9425
rect 3271 9382 3280 9416
rect 3280 9382 3314 9416
rect 3314 9382 3323 9416
rect 3271 9373 3323 9382
rect 4903 9416 4955 9425
rect 4903 9382 4912 9416
rect 4912 9382 4946 9416
rect 4946 9382 4955 9416
rect 4903 9373 4955 9382
rect 6535 9416 6587 9425
rect 6535 9382 6544 9416
rect 6544 9382 6578 9416
rect 6578 9382 6587 9416
rect 6535 9373 6587 9382
rect 8167 9416 8219 9425
rect 8167 9382 8176 9416
rect 8176 9382 8210 9416
rect 8210 9382 8219 9416
rect 8167 9373 8219 9382
rect 9799 9416 9851 9425
rect 9799 9382 9808 9416
rect 9808 9382 9842 9416
rect 9842 9382 9851 9416
rect 9799 9373 9851 9382
rect 7 9212 59 9221
rect 7 9178 16 9212
rect 16 9178 50 9212
rect 50 9178 59 9212
rect 7 9169 59 9178
rect 1639 9212 1691 9221
rect 1639 9178 1648 9212
rect 1648 9178 1682 9212
rect 1682 9178 1691 9212
rect 1639 9169 1691 9178
rect 3271 9212 3323 9221
rect 3271 9178 3280 9212
rect 3280 9178 3314 9212
rect 3314 9178 3323 9212
rect 3271 9169 3323 9178
rect 4903 9212 4955 9221
rect 4903 9178 4912 9212
rect 4912 9178 4946 9212
rect 4946 9178 4955 9212
rect 4903 9169 4955 9178
rect 6535 9212 6587 9221
rect 6535 9178 6544 9212
rect 6544 9178 6578 9212
rect 6578 9178 6587 9212
rect 6535 9169 6587 9178
rect 8167 9212 8219 9221
rect 8167 9178 8176 9212
rect 8176 9178 8210 9212
rect 8210 9178 8219 9212
rect 8167 9169 8219 9178
rect 9799 9212 9851 9221
rect 9799 9178 9808 9212
rect 9808 9178 9842 9212
rect 9842 9178 9851 9212
rect 9799 9169 9851 9178
rect 7 9008 59 9017
rect 7 8974 16 9008
rect 16 8974 50 9008
rect 50 8974 59 9008
rect 7 8965 59 8974
rect 1639 9008 1691 9017
rect 1639 8974 1648 9008
rect 1648 8974 1682 9008
rect 1682 8974 1691 9008
rect 1639 8965 1691 8974
rect 3271 9008 3323 9017
rect 3271 8974 3280 9008
rect 3280 8974 3314 9008
rect 3314 8974 3323 9008
rect 3271 8965 3323 8974
rect 4903 9008 4955 9017
rect 4903 8974 4912 9008
rect 4912 8974 4946 9008
rect 4946 8974 4955 9008
rect 4903 8965 4955 8974
rect 6535 9008 6587 9017
rect 6535 8974 6544 9008
rect 6544 8974 6578 9008
rect 6578 8974 6587 9008
rect 6535 8965 6587 8974
rect 8167 9008 8219 9017
rect 8167 8974 8176 9008
rect 8176 8974 8210 9008
rect 8210 8974 8219 9008
rect 8167 8965 8219 8974
rect 9799 9008 9851 9017
rect 9799 8974 9808 9008
rect 9808 8974 9842 9008
rect 9842 8974 9851 9008
rect 9799 8965 9851 8974
rect 7 8804 59 8813
rect 7 8770 16 8804
rect 16 8770 50 8804
rect 50 8770 59 8804
rect 7 8761 59 8770
rect 1639 8804 1691 8813
rect 1639 8770 1648 8804
rect 1648 8770 1682 8804
rect 1682 8770 1691 8804
rect 1639 8761 1691 8770
rect 3271 8804 3323 8813
rect 3271 8770 3280 8804
rect 3280 8770 3314 8804
rect 3314 8770 3323 8804
rect 3271 8761 3323 8770
rect 4903 8804 4955 8813
rect 4903 8770 4912 8804
rect 4912 8770 4946 8804
rect 4946 8770 4955 8804
rect 4903 8761 4955 8770
rect 6535 8804 6587 8813
rect 6535 8770 6544 8804
rect 6544 8770 6578 8804
rect 6578 8770 6587 8804
rect 6535 8761 6587 8770
rect 8167 8804 8219 8813
rect 8167 8770 8176 8804
rect 8176 8770 8210 8804
rect 8210 8770 8219 8804
rect 8167 8761 8219 8770
rect 9799 8804 9851 8813
rect 9799 8770 9808 8804
rect 9808 8770 9842 8804
rect 9842 8770 9851 8804
rect 9799 8761 9851 8770
rect 7 8600 59 8609
rect 7 8566 16 8600
rect 16 8566 50 8600
rect 50 8566 59 8600
rect 7 8557 59 8566
rect 1639 8600 1691 8609
rect 1639 8566 1648 8600
rect 1648 8566 1682 8600
rect 1682 8566 1691 8600
rect 1639 8557 1691 8566
rect 3271 8600 3323 8609
rect 3271 8566 3280 8600
rect 3280 8566 3314 8600
rect 3314 8566 3323 8600
rect 3271 8557 3323 8566
rect 4903 8600 4955 8609
rect 4903 8566 4912 8600
rect 4912 8566 4946 8600
rect 4946 8566 4955 8600
rect 4903 8557 4955 8566
rect 6535 8600 6587 8609
rect 6535 8566 6544 8600
rect 6544 8566 6578 8600
rect 6578 8566 6587 8600
rect 6535 8557 6587 8566
rect 8167 8600 8219 8609
rect 8167 8566 8176 8600
rect 8176 8566 8210 8600
rect 8210 8566 8219 8600
rect 8167 8557 8219 8566
rect 9799 8600 9851 8609
rect 9799 8566 9808 8600
rect 9808 8566 9842 8600
rect 9842 8566 9851 8600
rect 9799 8557 9851 8566
rect 7 8396 59 8405
rect 7 8362 16 8396
rect 16 8362 50 8396
rect 50 8362 59 8396
rect 7 8353 59 8362
rect 1639 8396 1691 8405
rect 1639 8362 1648 8396
rect 1648 8362 1682 8396
rect 1682 8362 1691 8396
rect 1639 8353 1691 8362
rect 3271 8396 3323 8405
rect 3271 8362 3280 8396
rect 3280 8362 3314 8396
rect 3314 8362 3323 8396
rect 3271 8353 3323 8362
rect 4903 8396 4955 8405
rect 4903 8362 4912 8396
rect 4912 8362 4946 8396
rect 4946 8362 4955 8396
rect 4903 8353 4955 8362
rect 6535 8396 6587 8405
rect 6535 8362 6544 8396
rect 6544 8362 6578 8396
rect 6578 8362 6587 8396
rect 6535 8353 6587 8362
rect 8167 8396 8219 8405
rect 8167 8362 8176 8396
rect 8176 8362 8210 8396
rect 8210 8362 8219 8396
rect 8167 8353 8219 8362
rect 9799 8396 9851 8405
rect 9799 8362 9808 8396
rect 9808 8362 9842 8396
rect 9842 8362 9851 8396
rect 9799 8353 9851 8362
rect 7 8192 59 8201
rect 7 8158 16 8192
rect 16 8158 50 8192
rect 50 8158 59 8192
rect 7 8149 59 8158
rect 1639 8192 1691 8201
rect 1639 8158 1648 8192
rect 1648 8158 1682 8192
rect 1682 8158 1691 8192
rect 1639 8149 1691 8158
rect 3271 8192 3323 8201
rect 3271 8158 3280 8192
rect 3280 8158 3314 8192
rect 3314 8158 3323 8192
rect 3271 8149 3323 8158
rect 4903 8192 4955 8201
rect 4903 8158 4912 8192
rect 4912 8158 4946 8192
rect 4946 8158 4955 8192
rect 4903 8149 4955 8158
rect 6535 8192 6587 8201
rect 6535 8158 6544 8192
rect 6544 8158 6578 8192
rect 6578 8158 6587 8192
rect 6535 8149 6587 8158
rect 8167 8192 8219 8201
rect 8167 8158 8176 8192
rect 8176 8158 8210 8192
rect 8210 8158 8219 8192
rect 8167 8149 8219 8158
rect 9799 8192 9851 8201
rect 9799 8158 9808 8192
rect 9808 8158 9842 8192
rect 9842 8158 9851 8192
rect 9799 8149 9851 8158
rect 7 7988 59 7997
rect 7 7954 16 7988
rect 16 7954 50 7988
rect 50 7954 59 7988
rect 7 7945 59 7954
rect 1639 7988 1691 7997
rect 1639 7954 1648 7988
rect 1648 7954 1682 7988
rect 1682 7954 1691 7988
rect 1639 7945 1691 7954
rect 3271 7988 3323 7997
rect 3271 7954 3280 7988
rect 3280 7954 3314 7988
rect 3314 7954 3323 7988
rect 3271 7945 3323 7954
rect 4903 7988 4955 7997
rect 4903 7954 4912 7988
rect 4912 7954 4946 7988
rect 4946 7954 4955 7988
rect 4903 7945 4955 7954
rect 6535 7988 6587 7997
rect 6535 7954 6544 7988
rect 6544 7954 6578 7988
rect 6578 7954 6587 7988
rect 6535 7945 6587 7954
rect 8167 7988 8219 7997
rect 8167 7954 8176 7988
rect 8176 7954 8210 7988
rect 8210 7954 8219 7988
rect 8167 7945 8219 7954
rect 9799 7988 9851 7997
rect 9799 7954 9808 7988
rect 9808 7954 9842 7988
rect 9842 7954 9851 7988
rect 9799 7945 9851 7954
rect 218 7834 270 7843
rect 218 7800 227 7834
rect 227 7800 261 7834
rect 261 7800 270 7834
rect 218 7791 270 7800
rect 422 7834 474 7843
rect 422 7800 431 7834
rect 431 7800 465 7834
rect 465 7800 474 7834
rect 422 7791 474 7800
rect 626 7834 678 7843
rect 626 7800 635 7834
rect 635 7800 669 7834
rect 669 7800 678 7834
rect 626 7791 678 7800
rect 830 7834 882 7843
rect 830 7800 839 7834
rect 839 7800 873 7834
rect 873 7800 882 7834
rect 830 7791 882 7800
rect 1034 7834 1086 7843
rect 1034 7800 1043 7834
rect 1043 7800 1077 7834
rect 1077 7800 1086 7834
rect 1034 7791 1086 7800
rect 1238 7834 1290 7843
rect 1238 7800 1247 7834
rect 1247 7800 1281 7834
rect 1281 7800 1290 7834
rect 1238 7791 1290 7800
rect 1442 7834 1494 7843
rect 1442 7800 1451 7834
rect 1451 7800 1485 7834
rect 1485 7800 1494 7834
rect 1442 7791 1494 7800
rect 1646 7834 1698 7843
rect 1646 7800 1655 7834
rect 1655 7800 1689 7834
rect 1689 7800 1698 7834
rect 1646 7791 1698 7800
rect 1850 7834 1902 7843
rect 1850 7800 1859 7834
rect 1859 7800 1893 7834
rect 1893 7800 1902 7834
rect 1850 7791 1902 7800
rect 2054 7834 2106 7843
rect 2054 7800 2063 7834
rect 2063 7800 2097 7834
rect 2097 7800 2106 7834
rect 2054 7791 2106 7800
rect 2258 7834 2310 7843
rect 2258 7800 2267 7834
rect 2267 7800 2301 7834
rect 2301 7800 2310 7834
rect 2258 7791 2310 7800
rect 2462 7834 2514 7843
rect 2462 7800 2471 7834
rect 2471 7800 2505 7834
rect 2505 7800 2514 7834
rect 2462 7791 2514 7800
rect 2666 7834 2718 7843
rect 2666 7800 2675 7834
rect 2675 7800 2709 7834
rect 2709 7800 2718 7834
rect 2666 7791 2718 7800
rect 2870 7834 2922 7843
rect 2870 7800 2879 7834
rect 2879 7800 2913 7834
rect 2913 7800 2922 7834
rect 2870 7791 2922 7800
rect 3074 7834 3126 7843
rect 3074 7800 3083 7834
rect 3083 7800 3117 7834
rect 3117 7800 3126 7834
rect 3074 7791 3126 7800
rect 3278 7834 3330 7843
rect 3278 7800 3287 7834
rect 3287 7800 3321 7834
rect 3321 7800 3330 7834
rect 3278 7791 3330 7800
rect 3482 7834 3534 7843
rect 3482 7800 3491 7834
rect 3491 7800 3525 7834
rect 3525 7800 3534 7834
rect 3482 7791 3534 7800
rect 3686 7834 3738 7843
rect 3686 7800 3695 7834
rect 3695 7800 3729 7834
rect 3729 7800 3738 7834
rect 3686 7791 3738 7800
rect 3890 7834 3942 7843
rect 3890 7800 3899 7834
rect 3899 7800 3933 7834
rect 3933 7800 3942 7834
rect 3890 7791 3942 7800
rect 4094 7834 4146 7843
rect 4094 7800 4103 7834
rect 4103 7800 4137 7834
rect 4137 7800 4146 7834
rect 4094 7791 4146 7800
rect 4298 7834 4350 7843
rect 4298 7800 4307 7834
rect 4307 7800 4341 7834
rect 4341 7800 4350 7834
rect 4298 7791 4350 7800
rect 4502 7834 4554 7843
rect 4502 7800 4511 7834
rect 4511 7800 4545 7834
rect 4545 7800 4554 7834
rect 4502 7791 4554 7800
rect 4706 7834 4758 7843
rect 4706 7800 4715 7834
rect 4715 7800 4749 7834
rect 4749 7800 4758 7834
rect 4706 7791 4758 7800
rect 4910 7834 4962 7843
rect 4910 7800 4919 7834
rect 4919 7800 4953 7834
rect 4953 7800 4962 7834
rect 4910 7791 4962 7800
rect 5114 7834 5166 7843
rect 5114 7800 5123 7834
rect 5123 7800 5157 7834
rect 5157 7800 5166 7834
rect 5114 7791 5166 7800
rect 5318 7834 5370 7843
rect 5318 7800 5327 7834
rect 5327 7800 5361 7834
rect 5361 7800 5370 7834
rect 5318 7791 5370 7800
rect 5522 7834 5574 7843
rect 5522 7800 5531 7834
rect 5531 7800 5565 7834
rect 5565 7800 5574 7834
rect 5522 7791 5574 7800
rect 5726 7834 5778 7843
rect 5726 7800 5735 7834
rect 5735 7800 5769 7834
rect 5769 7800 5778 7834
rect 5726 7791 5778 7800
rect 5930 7834 5982 7843
rect 5930 7800 5939 7834
rect 5939 7800 5973 7834
rect 5973 7800 5982 7834
rect 5930 7791 5982 7800
rect 6134 7834 6186 7843
rect 6134 7800 6143 7834
rect 6143 7800 6177 7834
rect 6177 7800 6186 7834
rect 6134 7791 6186 7800
rect 6338 7834 6390 7843
rect 6338 7800 6347 7834
rect 6347 7800 6381 7834
rect 6381 7800 6390 7834
rect 6338 7791 6390 7800
rect 6542 7834 6594 7843
rect 6542 7800 6551 7834
rect 6551 7800 6585 7834
rect 6585 7800 6594 7834
rect 6542 7791 6594 7800
rect 6746 7834 6798 7843
rect 6746 7800 6755 7834
rect 6755 7800 6789 7834
rect 6789 7800 6798 7834
rect 6746 7791 6798 7800
rect 6950 7834 7002 7843
rect 6950 7800 6959 7834
rect 6959 7800 6993 7834
rect 6993 7800 7002 7834
rect 6950 7791 7002 7800
rect 7154 7834 7206 7843
rect 7154 7800 7163 7834
rect 7163 7800 7197 7834
rect 7197 7800 7206 7834
rect 7154 7791 7206 7800
rect 7358 7834 7410 7843
rect 7358 7800 7367 7834
rect 7367 7800 7401 7834
rect 7401 7800 7410 7834
rect 7358 7791 7410 7800
rect 7562 7834 7614 7843
rect 7562 7800 7571 7834
rect 7571 7800 7605 7834
rect 7605 7800 7614 7834
rect 7562 7791 7614 7800
rect 7766 7834 7818 7843
rect 7766 7800 7775 7834
rect 7775 7800 7809 7834
rect 7809 7800 7818 7834
rect 7766 7791 7818 7800
rect 7970 7834 8022 7843
rect 7970 7800 7979 7834
rect 7979 7800 8013 7834
rect 8013 7800 8022 7834
rect 7970 7791 8022 7800
rect 8174 7834 8226 7843
rect 8174 7800 8183 7834
rect 8183 7800 8217 7834
rect 8217 7800 8226 7834
rect 8174 7791 8226 7800
rect 8378 7834 8430 7843
rect 8378 7800 8387 7834
rect 8387 7800 8421 7834
rect 8421 7800 8430 7834
rect 8378 7791 8430 7800
rect 8582 7834 8634 7843
rect 8582 7800 8591 7834
rect 8591 7800 8625 7834
rect 8625 7800 8634 7834
rect 8582 7791 8634 7800
rect 8786 7834 8838 7843
rect 8786 7800 8795 7834
rect 8795 7800 8829 7834
rect 8829 7800 8838 7834
rect 8786 7791 8838 7800
rect 8990 7834 9042 7843
rect 8990 7800 8999 7834
rect 8999 7800 9033 7834
rect 9033 7800 9042 7834
rect 8990 7791 9042 7800
rect 9194 7834 9246 7843
rect 9194 7800 9203 7834
rect 9203 7800 9237 7834
rect 9237 7800 9246 7834
rect 9194 7791 9246 7800
rect 9398 7834 9450 7843
rect 9398 7800 9407 7834
rect 9407 7800 9441 7834
rect 9441 7800 9450 7834
rect 9398 7791 9450 7800
rect 9602 7834 9654 7843
rect 9602 7800 9611 7834
rect 9611 7800 9645 7834
rect 9645 7800 9654 7834
rect 9602 7791 9654 7800
rect 9820 7834 9872 7843
rect 9820 7800 9829 7834
rect 9829 7800 9863 7834
rect 9863 7800 9872 7834
rect 9820 7791 9872 7800
rect 7 7680 59 7689
rect 7 7646 16 7680
rect 16 7646 50 7680
rect 50 7646 59 7680
rect 7 7637 59 7646
rect 1639 7680 1691 7689
rect 1639 7646 1648 7680
rect 1648 7646 1682 7680
rect 1682 7646 1691 7680
rect 1639 7637 1691 7646
rect 3271 7680 3323 7689
rect 3271 7646 3280 7680
rect 3280 7646 3314 7680
rect 3314 7646 3323 7680
rect 3271 7637 3323 7646
rect 4903 7680 4955 7689
rect 4903 7646 4912 7680
rect 4912 7646 4946 7680
rect 4946 7646 4955 7680
rect 4903 7637 4955 7646
rect 6535 7680 6587 7689
rect 6535 7646 6544 7680
rect 6544 7646 6578 7680
rect 6578 7646 6587 7680
rect 6535 7637 6587 7646
rect 8167 7680 8219 7689
rect 8167 7646 8176 7680
rect 8176 7646 8210 7680
rect 8210 7646 8219 7680
rect 8167 7637 8219 7646
rect 9799 7680 9851 7689
rect 9799 7646 9808 7680
rect 9808 7646 9842 7680
rect 9842 7646 9851 7680
rect 9799 7637 9851 7646
rect 7 7476 59 7485
rect 7 7442 16 7476
rect 16 7442 50 7476
rect 50 7442 59 7476
rect 7 7433 59 7442
rect 1639 7476 1691 7485
rect 1639 7442 1648 7476
rect 1648 7442 1682 7476
rect 1682 7442 1691 7476
rect 1639 7433 1691 7442
rect 3271 7476 3323 7485
rect 3271 7442 3280 7476
rect 3280 7442 3314 7476
rect 3314 7442 3323 7476
rect 3271 7433 3323 7442
rect 4903 7476 4955 7485
rect 4903 7442 4912 7476
rect 4912 7442 4946 7476
rect 4946 7442 4955 7476
rect 4903 7433 4955 7442
rect 6535 7476 6587 7485
rect 6535 7442 6544 7476
rect 6544 7442 6578 7476
rect 6578 7442 6587 7476
rect 6535 7433 6587 7442
rect 8167 7476 8219 7485
rect 8167 7442 8176 7476
rect 8176 7442 8210 7476
rect 8210 7442 8219 7476
rect 8167 7433 8219 7442
rect 9799 7476 9851 7485
rect 9799 7442 9808 7476
rect 9808 7442 9842 7476
rect 9842 7442 9851 7476
rect 9799 7433 9851 7442
rect 7 7272 59 7281
rect 7 7238 16 7272
rect 16 7238 50 7272
rect 50 7238 59 7272
rect 7 7229 59 7238
rect 1639 7272 1691 7281
rect 1639 7238 1648 7272
rect 1648 7238 1682 7272
rect 1682 7238 1691 7272
rect 1639 7229 1691 7238
rect 3271 7272 3323 7281
rect 3271 7238 3280 7272
rect 3280 7238 3314 7272
rect 3314 7238 3323 7272
rect 3271 7229 3323 7238
rect 4903 7272 4955 7281
rect 4903 7238 4912 7272
rect 4912 7238 4946 7272
rect 4946 7238 4955 7272
rect 4903 7229 4955 7238
rect 6535 7272 6587 7281
rect 6535 7238 6544 7272
rect 6544 7238 6578 7272
rect 6578 7238 6587 7272
rect 6535 7229 6587 7238
rect 8167 7272 8219 7281
rect 8167 7238 8176 7272
rect 8176 7238 8210 7272
rect 8210 7238 8219 7272
rect 8167 7229 8219 7238
rect 9799 7272 9851 7281
rect 9799 7238 9808 7272
rect 9808 7238 9842 7272
rect 9842 7238 9851 7272
rect 9799 7229 9851 7238
rect 7 7068 59 7077
rect 7 7034 16 7068
rect 16 7034 50 7068
rect 50 7034 59 7068
rect 7 7025 59 7034
rect 1639 7068 1691 7077
rect 1639 7034 1648 7068
rect 1648 7034 1682 7068
rect 1682 7034 1691 7068
rect 1639 7025 1691 7034
rect 3271 7068 3323 7077
rect 3271 7034 3280 7068
rect 3280 7034 3314 7068
rect 3314 7034 3323 7068
rect 3271 7025 3323 7034
rect 4903 7068 4955 7077
rect 4903 7034 4912 7068
rect 4912 7034 4946 7068
rect 4946 7034 4955 7068
rect 4903 7025 4955 7034
rect 6535 7068 6587 7077
rect 6535 7034 6544 7068
rect 6544 7034 6578 7068
rect 6578 7034 6587 7068
rect 6535 7025 6587 7034
rect 8167 7068 8219 7077
rect 8167 7034 8176 7068
rect 8176 7034 8210 7068
rect 8210 7034 8219 7068
rect 8167 7025 8219 7034
rect 9799 7068 9851 7077
rect 9799 7034 9808 7068
rect 9808 7034 9842 7068
rect 9842 7034 9851 7068
rect 9799 7025 9851 7034
rect 7 6864 59 6873
rect 7 6830 16 6864
rect 16 6830 50 6864
rect 50 6830 59 6864
rect 7 6821 59 6830
rect 1639 6864 1691 6873
rect 1639 6830 1648 6864
rect 1648 6830 1682 6864
rect 1682 6830 1691 6864
rect 1639 6821 1691 6830
rect 3271 6864 3323 6873
rect 3271 6830 3280 6864
rect 3280 6830 3314 6864
rect 3314 6830 3323 6864
rect 3271 6821 3323 6830
rect 4903 6864 4955 6873
rect 4903 6830 4912 6864
rect 4912 6830 4946 6864
rect 4946 6830 4955 6864
rect 4903 6821 4955 6830
rect 6535 6864 6587 6873
rect 6535 6830 6544 6864
rect 6544 6830 6578 6864
rect 6578 6830 6587 6864
rect 6535 6821 6587 6830
rect 8167 6864 8219 6873
rect 8167 6830 8176 6864
rect 8176 6830 8210 6864
rect 8210 6830 8219 6864
rect 8167 6821 8219 6830
rect 9799 6864 9851 6873
rect 9799 6830 9808 6864
rect 9808 6830 9842 6864
rect 9842 6830 9851 6864
rect 9799 6821 9851 6830
rect 7 6660 59 6669
rect 7 6626 16 6660
rect 16 6626 50 6660
rect 50 6626 59 6660
rect 7 6617 59 6626
rect 1639 6660 1691 6669
rect 1639 6626 1648 6660
rect 1648 6626 1682 6660
rect 1682 6626 1691 6660
rect 1639 6617 1691 6626
rect 3271 6660 3323 6669
rect 3271 6626 3280 6660
rect 3280 6626 3314 6660
rect 3314 6626 3323 6660
rect 3271 6617 3323 6626
rect 4903 6660 4955 6669
rect 4903 6626 4912 6660
rect 4912 6626 4946 6660
rect 4946 6626 4955 6660
rect 4903 6617 4955 6626
rect 6535 6660 6587 6669
rect 6535 6626 6544 6660
rect 6544 6626 6578 6660
rect 6578 6626 6587 6660
rect 6535 6617 6587 6626
rect 8167 6660 8219 6669
rect 8167 6626 8176 6660
rect 8176 6626 8210 6660
rect 8210 6626 8219 6660
rect 8167 6617 8219 6626
rect 9799 6660 9851 6669
rect 9799 6626 9808 6660
rect 9808 6626 9842 6660
rect 9842 6626 9851 6660
rect 9799 6617 9851 6626
rect 7 6456 59 6465
rect 7 6422 16 6456
rect 16 6422 50 6456
rect 50 6422 59 6456
rect 7 6413 59 6422
rect 1639 6456 1691 6465
rect 1639 6422 1648 6456
rect 1648 6422 1682 6456
rect 1682 6422 1691 6456
rect 1639 6413 1691 6422
rect 3271 6456 3323 6465
rect 3271 6422 3280 6456
rect 3280 6422 3314 6456
rect 3314 6422 3323 6456
rect 3271 6413 3323 6422
rect 4903 6456 4955 6465
rect 4903 6422 4912 6456
rect 4912 6422 4946 6456
rect 4946 6422 4955 6456
rect 4903 6413 4955 6422
rect 6535 6456 6587 6465
rect 6535 6422 6544 6456
rect 6544 6422 6578 6456
rect 6578 6422 6587 6456
rect 6535 6413 6587 6422
rect 8167 6456 8219 6465
rect 8167 6422 8176 6456
rect 8176 6422 8210 6456
rect 8210 6422 8219 6456
rect 8167 6413 8219 6422
rect 9799 6456 9851 6465
rect 9799 6422 9808 6456
rect 9808 6422 9842 6456
rect 9842 6422 9851 6456
rect 9799 6413 9851 6422
rect 7 6252 59 6261
rect 7 6218 16 6252
rect 16 6218 50 6252
rect 50 6218 59 6252
rect 7 6209 59 6218
rect 1639 6252 1691 6261
rect 1639 6218 1648 6252
rect 1648 6218 1682 6252
rect 1682 6218 1691 6252
rect 1639 6209 1691 6218
rect 3271 6252 3323 6261
rect 3271 6218 3280 6252
rect 3280 6218 3314 6252
rect 3314 6218 3323 6252
rect 3271 6209 3323 6218
rect 4903 6252 4955 6261
rect 4903 6218 4912 6252
rect 4912 6218 4946 6252
rect 4946 6218 4955 6252
rect 4903 6209 4955 6218
rect 6535 6252 6587 6261
rect 6535 6218 6544 6252
rect 6544 6218 6578 6252
rect 6578 6218 6587 6252
rect 6535 6209 6587 6218
rect 8167 6252 8219 6261
rect 8167 6218 8176 6252
rect 8176 6218 8210 6252
rect 8210 6218 8219 6252
rect 8167 6209 8219 6218
rect 9799 6252 9851 6261
rect 9799 6218 9808 6252
rect 9808 6218 9842 6252
rect 9842 6218 9851 6252
rect 9799 6209 9851 6218
rect 218 6098 270 6107
rect 218 6064 227 6098
rect 227 6064 261 6098
rect 261 6064 270 6098
rect 218 6055 270 6064
rect 422 6098 474 6107
rect 422 6064 431 6098
rect 431 6064 465 6098
rect 465 6064 474 6098
rect 422 6055 474 6064
rect 626 6098 678 6107
rect 626 6064 635 6098
rect 635 6064 669 6098
rect 669 6064 678 6098
rect 626 6055 678 6064
rect 830 6098 882 6107
rect 830 6064 839 6098
rect 839 6064 873 6098
rect 873 6064 882 6098
rect 830 6055 882 6064
rect 1034 6098 1086 6107
rect 1034 6064 1043 6098
rect 1043 6064 1077 6098
rect 1077 6064 1086 6098
rect 1034 6055 1086 6064
rect 1238 6098 1290 6107
rect 1238 6064 1247 6098
rect 1247 6064 1281 6098
rect 1281 6064 1290 6098
rect 1238 6055 1290 6064
rect 1442 6098 1494 6107
rect 1442 6064 1451 6098
rect 1451 6064 1485 6098
rect 1485 6064 1494 6098
rect 1442 6055 1494 6064
rect 1646 6098 1698 6107
rect 1646 6064 1655 6098
rect 1655 6064 1689 6098
rect 1689 6064 1698 6098
rect 1646 6055 1698 6064
rect 1850 6098 1902 6107
rect 1850 6064 1859 6098
rect 1859 6064 1893 6098
rect 1893 6064 1902 6098
rect 1850 6055 1902 6064
rect 2054 6098 2106 6107
rect 2054 6064 2063 6098
rect 2063 6064 2097 6098
rect 2097 6064 2106 6098
rect 2054 6055 2106 6064
rect 2258 6098 2310 6107
rect 2258 6064 2267 6098
rect 2267 6064 2301 6098
rect 2301 6064 2310 6098
rect 2258 6055 2310 6064
rect 2462 6098 2514 6107
rect 2462 6064 2471 6098
rect 2471 6064 2505 6098
rect 2505 6064 2514 6098
rect 2462 6055 2514 6064
rect 2666 6098 2718 6107
rect 2666 6064 2675 6098
rect 2675 6064 2709 6098
rect 2709 6064 2718 6098
rect 2666 6055 2718 6064
rect 2870 6098 2922 6107
rect 2870 6064 2879 6098
rect 2879 6064 2913 6098
rect 2913 6064 2922 6098
rect 2870 6055 2922 6064
rect 3074 6098 3126 6107
rect 3074 6064 3083 6098
rect 3083 6064 3117 6098
rect 3117 6064 3126 6098
rect 3074 6055 3126 6064
rect 3278 6098 3330 6107
rect 3278 6064 3287 6098
rect 3287 6064 3321 6098
rect 3321 6064 3330 6098
rect 3278 6055 3330 6064
rect 3482 6098 3534 6107
rect 3482 6064 3491 6098
rect 3491 6064 3525 6098
rect 3525 6064 3534 6098
rect 3482 6055 3534 6064
rect 3686 6098 3738 6107
rect 3686 6064 3695 6098
rect 3695 6064 3729 6098
rect 3729 6064 3738 6098
rect 3686 6055 3738 6064
rect 3890 6098 3942 6107
rect 3890 6064 3899 6098
rect 3899 6064 3933 6098
rect 3933 6064 3942 6098
rect 3890 6055 3942 6064
rect 4094 6098 4146 6107
rect 4094 6064 4103 6098
rect 4103 6064 4137 6098
rect 4137 6064 4146 6098
rect 4094 6055 4146 6064
rect 4298 6098 4350 6107
rect 4298 6064 4307 6098
rect 4307 6064 4341 6098
rect 4341 6064 4350 6098
rect 4298 6055 4350 6064
rect 4502 6098 4554 6107
rect 4502 6064 4511 6098
rect 4511 6064 4545 6098
rect 4545 6064 4554 6098
rect 4502 6055 4554 6064
rect 4706 6098 4758 6107
rect 4706 6064 4715 6098
rect 4715 6064 4749 6098
rect 4749 6064 4758 6098
rect 4706 6055 4758 6064
rect 4910 6098 4962 6107
rect 4910 6064 4919 6098
rect 4919 6064 4953 6098
rect 4953 6064 4962 6098
rect 4910 6055 4962 6064
rect 5114 6098 5166 6107
rect 5114 6064 5123 6098
rect 5123 6064 5157 6098
rect 5157 6064 5166 6098
rect 5114 6055 5166 6064
rect 5318 6098 5370 6107
rect 5318 6064 5327 6098
rect 5327 6064 5361 6098
rect 5361 6064 5370 6098
rect 5318 6055 5370 6064
rect 5522 6098 5574 6107
rect 5522 6064 5531 6098
rect 5531 6064 5565 6098
rect 5565 6064 5574 6098
rect 5522 6055 5574 6064
rect 5726 6098 5778 6107
rect 5726 6064 5735 6098
rect 5735 6064 5769 6098
rect 5769 6064 5778 6098
rect 5726 6055 5778 6064
rect 5930 6098 5982 6107
rect 5930 6064 5939 6098
rect 5939 6064 5973 6098
rect 5973 6064 5982 6098
rect 5930 6055 5982 6064
rect 6134 6098 6186 6107
rect 6134 6064 6143 6098
rect 6143 6064 6177 6098
rect 6177 6064 6186 6098
rect 6134 6055 6186 6064
rect 6338 6098 6390 6107
rect 6338 6064 6347 6098
rect 6347 6064 6381 6098
rect 6381 6064 6390 6098
rect 6338 6055 6390 6064
rect 6542 6098 6594 6107
rect 6542 6064 6551 6098
rect 6551 6064 6585 6098
rect 6585 6064 6594 6098
rect 6542 6055 6594 6064
rect 6746 6098 6798 6107
rect 6746 6064 6755 6098
rect 6755 6064 6789 6098
rect 6789 6064 6798 6098
rect 6746 6055 6798 6064
rect 6950 6098 7002 6107
rect 6950 6064 6959 6098
rect 6959 6064 6993 6098
rect 6993 6064 7002 6098
rect 6950 6055 7002 6064
rect 7154 6098 7206 6107
rect 7154 6064 7163 6098
rect 7163 6064 7197 6098
rect 7197 6064 7206 6098
rect 7154 6055 7206 6064
rect 7358 6098 7410 6107
rect 7358 6064 7367 6098
rect 7367 6064 7401 6098
rect 7401 6064 7410 6098
rect 7358 6055 7410 6064
rect 7562 6098 7614 6107
rect 7562 6064 7571 6098
rect 7571 6064 7605 6098
rect 7605 6064 7614 6098
rect 7562 6055 7614 6064
rect 7766 6098 7818 6107
rect 7766 6064 7775 6098
rect 7775 6064 7809 6098
rect 7809 6064 7818 6098
rect 7766 6055 7818 6064
rect 7970 6098 8022 6107
rect 7970 6064 7979 6098
rect 7979 6064 8013 6098
rect 8013 6064 8022 6098
rect 7970 6055 8022 6064
rect 8174 6098 8226 6107
rect 8174 6064 8183 6098
rect 8183 6064 8217 6098
rect 8217 6064 8226 6098
rect 8174 6055 8226 6064
rect 8378 6098 8430 6107
rect 8378 6064 8387 6098
rect 8387 6064 8421 6098
rect 8421 6064 8430 6098
rect 8378 6055 8430 6064
rect 8582 6098 8634 6107
rect 8582 6064 8591 6098
rect 8591 6064 8625 6098
rect 8625 6064 8634 6098
rect 8582 6055 8634 6064
rect 8786 6098 8838 6107
rect 8786 6064 8795 6098
rect 8795 6064 8829 6098
rect 8829 6064 8838 6098
rect 8786 6055 8838 6064
rect 8990 6098 9042 6107
rect 8990 6064 8999 6098
rect 8999 6064 9033 6098
rect 9033 6064 9042 6098
rect 8990 6055 9042 6064
rect 9194 6098 9246 6107
rect 9194 6064 9203 6098
rect 9203 6064 9237 6098
rect 9237 6064 9246 6098
rect 9194 6055 9246 6064
rect 9398 6098 9450 6107
rect 9398 6064 9407 6098
rect 9407 6064 9441 6098
rect 9441 6064 9450 6098
rect 9398 6055 9450 6064
rect 9602 6098 9654 6107
rect 9602 6064 9611 6098
rect 9611 6064 9645 6098
rect 9645 6064 9654 6098
rect 9602 6055 9654 6064
rect 9820 6098 9872 6107
rect 9820 6064 9829 6098
rect 9829 6064 9863 6098
rect 9863 6064 9872 6098
rect 9820 6055 9872 6064
rect 7 5944 59 5953
rect 7 5910 16 5944
rect 16 5910 50 5944
rect 50 5910 59 5944
rect 7 5901 59 5910
rect 1639 5944 1691 5953
rect 1639 5910 1648 5944
rect 1648 5910 1682 5944
rect 1682 5910 1691 5944
rect 1639 5901 1691 5910
rect 3271 5944 3323 5953
rect 3271 5910 3280 5944
rect 3280 5910 3314 5944
rect 3314 5910 3323 5944
rect 3271 5901 3323 5910
rect 4903 5944 4955 5953
rect 4903 5910 4912 5944
rect 4912 5910 4946 5944
rect 4946 5910 4955 5944
rect 4903 5901 4955 5910
rect 6535 5944 6587 5953
rect 6535 5910 6544 5944
rect 6544 5910 6578 5944
rect 6578 5910 6587 5944
rect 6535 5901 6587 5910
rect 8167 5944 8219 5953
rect 8167 5910 8176 5944
rect 8176 5910 8210 5944
rect 8210 5910 8219 5944
rect 8167 5901 8219 5910
rect 9799 5944 9851 5953
rect 9799 5910 9808 5944
rect 9808 5910 9842 5944
rect 9842 5910 9851 5944
rect 9799 5901 9851 5910
rect 7 5740 59 5749
rect 7 5706 16 5740
rect 16 5706 50 5740
rect 50 5706 59 5740
rect 7 5697 59 5706
rect 1639 5740 1691 5749
rect 1639 5706 1648 5740
rect 1648 5706 1682 5740
rect 1682 5706 1691 5740
rect 1639 5697 1691 5706
rect 3271 5740 3323 5749
rect 3271 5706 3280 5740
rect 3280 5706 3314 5740
rect 3314 5706 3323 5740
rect 3271 5697 3323 5706
rect 4903 5740 4955 5749
rect 4903 5706 4912 5740
rect 4912 5706 4946 5740
rect 4946 5706 4955 5740
rect 4903 5697 4955 5706
rect 6535 5740 6587 5749
rect 6535 5706 6544 5740
rect 6544 5706 6578 5740
rect 6578 5706 6587 5740
rect 6535 5697 6587 5706
rect 8167 5740 8219 5749
rect 8167 5706 8176 5740
rect 8176 5706 8210 5740
rect 8210 5706 8219 5740
rect 8167 5697 8219 5706
rect 9799 5740 9851 5749
rect 9799 5706 9808 5740
rect 9808 5706 9842 5740
rect 9842 5706 9851 5740
rect 9799 5697 9851 5706
rect 7 5536 59 5545
rect 7 5502 16 5536
rect 16 5502 50 5536
rect 50 5502 59 5536
rect 7 5493 59 5502
rect 1639 5536 1691 5545
rect 1639 5502 1648 5536
rect 1648 5502 1682 5536
rect 1682 5502 1691 5536
rect 1639 5493 1691 5502
rect 3271 5536 3323 5545
rect 3271 5502 3280 5536
rect 3280 5502 3314 5536
rect 3314 5502 3323 5536
rect 3271 5493 3323 5502
rect 4903 5536 4955 5545
rect 4903 5502 4912 5536
rect 4912 5502 4946 5536
rect 4946 5502 4955 5536
rect 4903 5493 4955 5502
rect 6535 5536 6587 5545
rect 6535 5502 6544 5536
rect 6544 5502 6578 5536
rect 6578 5502 6587 5536
rect 6535 5493 6587 5502
rect 8167 5536 8219 5545
rect 8167 5502 8176 5536
rect 8176 5502 8210 5536
rect 8210 5502 8219 5536
rect 8167 5493 8219 5502
rect 9799 5536 9851 5545
rect 9799 5502 9808 5536
rect 9808 5502 9842 5536
rect 9842 5502 9851 5536
rect 9799 5493 9851 5502
rect 7 5332 59 5341
rect 7 5298 16 5332
rect 16 5298 50 5332
rect 50 5298 59 5332
rect 7 5289 59 5298
rect 1639 5332 1691 5341
rect 1639 5298 1648 5332
rect 1648 5298 1682 5332
rect 1682 5298 1691 5332
rect 1639 5289 1691 5298
rect 3271 5332 3323 5341
rect 3271 5298 3280 5332
rect 3280 5298 3314 5332
rect 3314 5298 3323 5332
rect 3271 5289 3323 5298
rect 4903 5332 4955 5341
rect 4903 5298 4912 5332
rect 4912 5298 4946 5332
rect 4946 5298 4955 5332
rect 4903 5289 4955 5298
rect 6535 5332 6587 5341
rect 6535 5298 6544 5332
rect 6544 5298 6578 5332
rect 6578 5298 6587 5332
rect 6535 5289 6587 5298
rect 8167 5332 8219 5341
rect 8167 5298 8176 5332
rect 8176 5298 8210 5332
rect 8210 5298 8219 5332
rect 8167 5289 8219 5298
rect 9799 5332 9851 5341
rect 9799 5298 9808 5332
rect 9808 5298 9842 5332
rect 9842 5298 9851 5332
rect 9799 5289 9851 5298
rect 7 5128 59 5137
rect 7 5094 16 5128
rect 16 5094 50 5128
rect 50 5094 59 5128
rect 7 5085 59 5094
rect 1639 5128 1691 5137
rect 1639 5094 1648 5128
rect 1648 5094 1682 5128
rect 1682 5094 1691 5128
rect 1639 5085 1691 5094
rect 3271 5128 3323 5137
rect 3271 5094 3280 5128
rect 3280 5094 3314 5128
rect 3314 5094 3323 5128
rect 3271 5085 3323 5094
rect 4903 5128 4955 5137
rect 4903 5094 4912 5128
rect 4912 5094 4946 5128
rect 4946 5094 4955 5128
rect 4903 5085 4955 5094
rect 6535 5128 6587 5137
rect 6535 5094 6544 5128
rect 6544 5094 6578 5128
rect 6578 5094 6587 5128
rect 6535 5085 6587 5094
rect 8167 5128 8219 5137
rect 8167 5094 8176 5128
rect 8176 5094 8210 5128
rect 8210 5094 8219 5128
rect 8167 5085 8219 5094
rect 9799 5128 9851 5137
rect 9799 5094 9808 5128
rect 9808 5094 9842 5128
rect 9842 5094 9851 5128
rect 9799 5085 9851 5094
rect 7 4924 59 4933
rect 7 4890 16 4924
rect 16 4890 50 4924
rect 50 4890 59 4924
rect 7 4881 59 4890
rect 1639 4924 1691 4933
rect 1639 4890 1648 4924
rect 1648 4890 1682 4924
rect 1682 4890 1691 4924
rect 1639 4881 1691 4890
rect 3271 4924 3323 4933
rect 3271 4890 3280 4924
rect 3280 4890 3314 4924
rect 3314 4890 3323 4924
rect 3271 4881 3323 4890
rect 4903 4924 4955 4933
rect 4903 4890 4912 4924
rect 4912 4890 4946 4924
rect 4946 4890 4955 4924
rect 4903 4881 4955 4890
rect 6535 4924 6587 4933
rect 6535 4890 6544 4924
rect 6544 4890 6578 4924
rect 6578 4890 6587 4924
rect 6535 4881 6587 4890
rect 8167 4924 8219 4933
rect 8167 4890 8176 4924
rect 8176 4890 8210 4924
rect 8210 4890 8219 4924
rect 8167 4881 8219 4890
rect 9799 4924 9851 4933
rect 9799 4890 9808 4924
rect 9808 4890 9842 4924
rect 9842 4890 9851 4924
rect 9799 4881 9851 4890
rect 7 4720 59 4729
rect 7 4686 16 4720
rect 16 4686 50 4720
rect 50 4686 59 4720
rect 7 4677 59 4686
rect 1639 4720 1691 4729
rect 1639 4686 1648 4720
rect 1648 4686 1682 4720
rect 1682 4686 1691 4720
rect 1639 4677 1691 4686
rect 3271 4720 3323 4729
rect 3271 4686 3280 4720
rect 3280 4686 3314 4720
rect 3314 4686 3323 4720
rect 3271 4677 3323 4686
rect 4903 4720 4955 4729
rect 4903 4686 4912 4720
rect 4912 4686 4946 4720
rect 4946 4686 4955 4720
rect 4903 4677 4955 4686
rect 6535 4720 6587 4729
rect 6535 4686 6544 4720
rect 6544 4686 6578 4720
rect 6578 4686 6587 4720
rect 6535 4677 6587 4686
rect 8167 4720 8219 4729
rect 8167 4686 8176 4720
rect 8176 4686 8210 4720
rect 8210 4686 8219 4720
rect 8167 4677 8219 4686
rect 9799 4720 9851 4729
rect 9799 4686 9808 4720
rect 9808 4686 9842 4720
rect 9842 4686 9851 4720
rect 9799 4677 9851 4686
rect 7 4516 59 4525
rect 7 4482 16 4516
rect 16 4482 50 4516
rect 50 4482 59 4516
rect 7 4473 59 4482
rect 1639 4516 1691 4525
rect 1639 4482 1648 4516
rect 1648 4482 1682 4516
rect 1682 4482 1691 4516
rect 1639 4473 1691 4482
rect 3271 4516 3323 4525
rect 3271 4482 3280 4516
rect 3280 4482 3314 4516
rect 3314 4482 3323 4516
rect 3271 4473 3323 4482
rect 4903 4516 4955 4525
rect 4903 4482 4912 4516
rect 4912 4482 4946 4516
rect 4946 4482 4955 4516
rect 4903 4473 4955 4482
rect 6535 4516 6587 4525
rect 6535 4482 6544 4516
rect 6544 4482 6578 4516
rect 6578 4482 6587 4516
rect 6535 4473 6587 4482
rect 8167 4516 8219 4525
rect 8167 4482 8176 4516
rect 8176 4482 8210 4516
rect 8210 4482 8219 4516
rect 8167 4473 8219 4482
rect 9799 4516 9851 4525
rect 9799 4482 9808 4516
rect 9808 4482 9842 4516
rect 9842 4482 9851 4516
rect 9799 4473 9851 4482
rect 218 4362 270 4371
rect 218 4328 227 4362
rect 227 4328 261 4362
rect 261 4328 270 4362
rect 218 4319 270 4328
rect 422 4362 474 4371
rect 422 4328 431 4362
rect 431 4328 465 4362
rect 465 4328 474 4362
rect 422 4319 474 4328
rect 626 4362 678 4371
rect 626 4328 635 4362
rect 635 4328 669 4362
rect 669 4328 678 4362
rect 626 4319 678 4328
rect 830 4362 882 4371
rect 830 4328 839 4362
rect 839 4328 873 4362
rect 873 4328 882 4362
rect 830 4319 882 4328
rect 1034 4362 1086 4371
rect 1034 4328 1043 4362
rect 1043 4328 1077 4362
rect 1077 4328 1086 4362
rect 1034 4319 1086 4328
rect 1238 4362 1290 4371
rect 1238 4328 1247 4362
rect 1247 4328 1281 4362
rect 1281 4328 1290 4362
rect 1238 4319 1290 4328
rect 1442 4362 1494 4371
rect 1442 4328 1451 4362
rect 1451 4328 1485 4362
rect 1485 4328 1494 4362
rect 1442 4319 1494 4328
rect 1646 4362 1698 4371
rect 1646 4328 1655 4362
rect 1655 4328 1689 4362
rect 1689 4328 1698 4362
rect 1646 4319 1698 4328
rect 1850 4362 1902 4371
rect 1850 4328 1859 4362
rect 1859 4328 1893 4362
rect 1893 4328 1902 4362
rect 1850 4319 1902 4328
rect 2054 4362 2106 4371
rect 2054 4328 2063 4362
rect 2063 4328 2097 4362
rect 2097 4328 2106 4362
rect 2054 4319 2106 4328
rect 2258 4362 2310 4371
rect 2258 4328 2267 4362
rect 2267 4328 2301 4362
rect 2301 4328 2310 4362
rect 2258 4319 2310 4328
rect 2462 4362 2514 4371
rect 2462 4328 2471 4362
rect 2471 4328 2505 4362
rect 2505 4328 2514 4362
rect 2462 4319 2514 4328
rect 2666 4362 2718 4371
rect 2666 4328 2675 4362
rect 2675 4328 2709 4362
rect 2709 4328 2718 4362
rect 2666 4319 2718 4328
rect 2870 4362 2922 4371
rect 2870 4328 2879 4362
rect 2879 4328 2913 4362
rect 2913 4328 2922 4362
rect 2870 4319 2922 4328
rect 3074 4362 3126 4371
rect 3074 4328 3083 4362
rect 3083 4328 3117 4362
rect 3117 4328 3126 4362
rect 3074 4319 3126 4328
rect 3278 4362 3330 4371
rect 3278 4328 3287 4362
rect 3287 4328 3321 4362
rect 3321 4328 3330 4362
rect 3278 4319 3330 4328
rect 3482 4362 3534 4371
rect 3482 4328 3491 4362
rect 3491 4328 3525 4362
rect 3525 4328 3534 4362
rect 3482 4319 3534 4328
rect 3686 4362 3738 4371
rect 3686 4328 3695 4362
rect 3695 4328 3729 4362
rect 3729 4328 3738 4362
rect 3686 4319 3738 4328
rect 3890 4362 3942 4371
rect 3890 4328 3899 4362
rect 3899 4328 3933 4362
rect 3933 4328 3942 4362
rect 3890 4319 3942 4328
rect 4094 4362 4146 4371
rect 4094 4328 4103 4362
rect 4103 4328 4137 4362
rect 4137 4328 4146 4362
rect 4094 4319 4146 4328
rect 4298 4362 4350 4371
rect 4298 4328 4307 4362
rect 4307 4328 4341 4362
rect 4341 4328 4350 4362
rect 4298 4319 4350 4328
rect 4502 4362 4554 4371
rect 4502 4328 4511 4362
rect 4511 4328 4545 4362
rect 4545 4328 4554 4362
rect 4502 4319 4554 4328
rect 4706 4362 4758 4371
rect 4706 4328 4715 4362
rect 4715 4328 4749 4362
rect 4749 4328 4758 4362
rect 4706 4319 4758 4328
rect 4910 4362 4962 4371
rect 4910 4328 4919 4362
rect 4919 4328 4953 4362
rect 4953 4328 4962 4362
rect 4910 4319 4962 4328
rect 5114 4362 5166 4371
rect 5114 4328 5123 4362
rect 5123 4328 5157 4362
rect 5157 4328 5166 4362
rect 5114 4319 5166 4328
rect 5318 4362 5370 4371
rect 5318 4328 5327 4362
rect 5327 4328 5361 4362
rect 5361 4328 5370 4362
rect 5318 4319 5370 4328
rect 5522 4362 5574 4371
rect 5522 4328 5531 4362
rect 5531 4328 5565 4362
rect 5565 4328 5574 4362
rect 5522 4319 5574 4328
rect 5726 4362 5778 4371
rect 5726 4328 5735 4362
rect 5735 4328 5769 4362
rect 5769 4328 5778 4362
rect 5726 4319 5778 4328
rect 5930 4362 5982 4371
rect 5930 4328 5939 4362
rect 5939 4328 5973 4362
rect 5973 4328 5982 4362
rect 5930 4319 5982 4328
rect 6134 4362 6186 4371
rect 6134 4328 6143 4362
rect 6143 4328 6177 4362
rect 6177 4328 6186 4362
rect 6134 4319 6186 4328
rect 6338 4362 6390 4371
rect 6338 4328 6347 4362
rect 6347 4328 6381 4362
rect 6381 4328 6390 4362
rect 6338 4319 6390 4328
rect 6542 4362 6594 4371
rect 6542 4328 6551 4362
rect 6551 4328 6585 4362
rect 6585 4328 6594 4362
rect 6542 4319 6594 4328
rect 6746 4362 6798 4371
rect 6746 4328 6755 4362
rect 6755 4328 6789 4362
rect 6789 4328 6798 4362
rect 6746 4319 6798 4328
rect 6950 4362 7002 4371
rect 6950 4328 6959 4362
rect 6959 4328 6993 4362
rect 6993 4328 7002 4362
rect 6950 4319 7002 4328
rect 7154 4362 7206 4371
rect 7154 4328 7163 4362
rect 7163 4328 7197 4362
rect 7197 4328 7206 4362
rect 7154 4319 7206 4328
rect 7358 4362 7410 4371
rect 7358 4328 7367 4362
rect 7367 4328 7401 4362
rect 7401 4328 7410 4362
rect 7358 4319 7410 4328
rect 7562 4362 7614 4371
rect 7562 4328 7571 4362
rect 7571 4328 7605 4362
rect 7605 4328 7614 4362
rect 7562 4319 7614 4328
rect 7766 4362 7818 4371
rect 7766 4328 7775 4362
rect 7775 4328 7809 4362
rect 7809 4328 7818 4362
rect 7766 4319 7818 4328
rect 7970 4362 8022 4371
rect 7970 4328 7979 4362
rect 7979 4328 8013 4362
rect 8013 4328 8022 4362
rect 7970 4319 8022 4328
rect 8174 4362 8226 4371
rect 8174 4328 8183 4362
rect 8183 4328 8217 4362
rect 8217 4328 8226 4362
rect 8174 4319 8226 4328
rect 8378 4362 8430 4371
rect 8378 4328 8387 4362
rect 8387 4328 8421 4362
rect 8421 4328 8430 4362
rect 8378 4319 8430 4328
rect 8582 4362 8634 4371
rect 8582 4328 8591 4362
rect 8591 4328 8625 4362
rect 8625 4328 8634 4362
rect 8582 4319 8634 4328
rect 8786 4362 8838 4371
rect 8786 4328 8795 4362
rect 8795 4328 8829 4362
rect 8829 4328 8838 4362
rect 8786 4319 8838 4328
rect 8990 4362 9042 4371
rect 8990 4328 8999 4362
rect 8999 4328 9033 4362
rect 9033 4328 9042 4362
rect 8990 4319 9042 4328
rect 9194 4362 9246 4371
rect 9194 4328 9203 4362
rect 9203 4328 9237 4362
rect 9237 4328 9246 4362
rect 9194 4319 9246 4328
rect 9398 4362 9450 4371
rect 9398 4328 9407 4362
rect 9407 4328 9441 4362
rect 9441 4328 9450 4362
rect 9398 4319 9450 4328
rect 9602 4362 9654 4371
rect 9602 4328 9611 4362
rect 9611 4328 9645 4362
rect 9645 4328 9654 4362
rect 9602 4319 9654 4328
rect 9820 4362 9872 4371
rect 9820 4328 9829 4362
rect 9829 4328 9863 4362
rect 9863 4328 9872 4362
rect 9820 4319 9872 4328
rect 7 4208 59 4217
rect 7 4174 16 4208
rect 16 4174 50 4208
rect 50 4174 59 4208
rect 7 4165 59 4174
rect 1639 4208 1691 4217
rect 1639 4174 1648 4208
rect 1648 4174 1682 4208
rect 1682 4174 1691 4208
rect 1639 4165 1691 4174
rect 3271 4208 3323 4217
rect 3271 4174 3280 4208
rect 3280 4174 3314 4208
rect 3314 4174 3323 4208
rect 3271 4165 3323 4174
rect 4903 4208 4955 4217
rect 4903 4174 4912 4208
rect 4912 4174 4946 4208
rect 4946 4174 4955 4208
rect 4903 4165 4955 4174
rect 6535 4208 6587 4217
rect 6535 4174 6544 4208
rect 6544 4174 6578 4208
rect 6578 4174 6587 4208
rect 6535 4165 6587 4174
rect 8167 4208 8219 4217
rect 8167 4174 8176 4208
rect 8176 4174 8210 4208
rect 8210 4174 8219 4208
rect 8167 4165 8219 4174
rect 9799 4208 9851 4217
rect 9799 4174 9808 4208
rect 9808 4174 9842 4208
rect 9842 4174 9851 4208
rect 9799 4165 9851 4174
rect 7 4004 59 4013
rect 7 3970 16 4004
rect 16 3970 50 4004
rect 50 3970 59 4004
rect 7 3961 59 3970
rect 1639 4004 1691 4013
rect 1639 3970 1648 4004
rect 1648 3970 1682 4004
rect 1682 3970 1691 4004
rect 1639 3961 1691 3970
rect 3271 4004 3323 4013
rect 3271 3970 3280 4004
rect 3280 3970 3314 4004
rect 3314 3970 3323 4004
rect 3271 3961 3323 3970
rect 4903 4004 4955 4013
rect 4903 3970 4912 4004
rect 4912 3970 4946 4004
rect 4946 3970 4955 4004
rect 4903 3961 4955 3970
rect 6535 4004 6587 4013
rect 6535 3970 6544 4004
rect 6544 3970 6578 4004
rect 6578 3970 6587 4004
rect 6535 3961 6587 3970
rect 8167 4004 8219 4013
rect 8167 3970 8176 4004
rect 8176 3970 8210 4004
rect 8210 3970 8219 4004
rect 8167 3961 8219 3970
rect 9799 4004 9851 4013
rect 9799 3970 9808 4004
rect 9808 3970 9842 4004
rect 9842 3970 9851 4004
rect 9799 3961 9851 3970
rect 7 3800 59 3809
rect 7 3766 16 3800
rect 16 3766 50 3800
rect 50 3766 59 3800
rect 7 3757 59 3766
rect 1639 3800 1691 3809
rect 1639 3766 1648 3800
rect 1648 3766 1682 3800
rect 1682 3766 1691 3800
rect 1639 3757 1691 3766
rect 3271 3800 3323 3809
rect 3271 3766 3280 3800
rect 3280 3766 3314 3800
rect 3314 3766 3323 3800
rect 3271 3757 3323 3766
rect 4903 3800 4955 3809
rect 4903 3766 4912 3800
rect 4912 3766 4946 3800
rect 4946 3766 4955 3800
rect 4903 3757 4955 3766
rect 6535 3800 6587 3809
rect 6535 3766 6544 3800
rect 6544 3766 6578 3800
rect 6578 3766 6587 3800
rect 6535 3757 6587 3766
rect 8167 3800 8219 3809
rect 8167 3766 8176 3800
rect 8176 3766 8210 3800
rect 8210 3766 8219 3800
rect 8167 3757 8219 3766
rect 9799 3800 9851 3809
rect 9799 3766 9808 3800
rect 9808 3766 9842 3800
rect 9842 3766 9851 3800
rect 9799 3757 9851 3766
rect 7 3596 59 3605
rect 7 3562 16 3596
rect 16 3562 50 3596
rect 50 3562 59 3596
rect 7 3553 59 3562
rect 1639 3596 1691 3605
rect 1639 3562 1648 3596
rect 1648 3562 1682 3596
rect 1682 3562 1691 3596
rect 1639 3553 1691 3562
rect 3271 3596 3323 3605
rect 3271 3562 3280 3596
rect 3280 3562 3314 3596
rect 3314 3562 3323 3596
rect 3271 3553 3323 3562
rect 4903 3596 4955 3605
rect 4903 3562 4912 3596
rect 4912 3562 4946 3596
rect 4946 3562 4955 3596
rect 4903 3553 4955 3562
rect 6535 3596 6587 3605
rect 6535 3562 6544 3596
rect 6544 3562 6578 3596
rect 6578 3562 6587 3596
rect 6535 3553 6587 3562
rect 8167 3596 8219 3605
rect 8167 3562 8176 3596
rect 8176 3562 8210 3596
rect 8210 3562 8219 3596
rect 8167 3553 8219 3562
rect 9799 3596 9851 3605
rect 9799 3562 9808 3596
rect 9808 3562 9842 3596
rect 9842 3562 9851 3596
rect 9799 3553 9851 3562
rect 7 3392 59 3401
rect 7 3358 16 3392
rect 16 3358 50 3392
rect 50 3358 59 3392
rect 7 3349 59 3358
rect 1639 3392 1691 3401
rect 1639 3358 1648 3392
rect 1648 3358 1682 3392
rect 1682 3358 1691 3392
rect 1639 3349 1691 3358
rect 3271 3392 3323 3401
rect 3271 3358 3280 3392
rect 3280 3358 3314 3392
rect 3314 3358 3323 3392
rect 3271 3349 3323 3358
rect 4903 3392 4955 3401
rect 4903 3358 4912 3392
rect 4912 3358 4946 3392
rect 4946 3358 4955 3392
rect 4903 3349 4955 3358
rect 6535 3392 6587 3401
rect 6535 3358 6544 3392
rect 6544 3358 6578 3392
rect 6578 3358 6587 3392
rect 6535 3349 6587 3358
rect 8167 3392 8219 3401
rect 8167 3358 8176 3392
rect 8176 3358 8210 3392
rect 8210 3358 8219 3392
rect 8167 3349 8219 3358
rect 9799 3392 9851 3401
rect 9799 3358 9808 3392
rect 9808 3358 9842 3392
rect 9842 3358 9851 3392
rect 9799 3349 9851 3358
rect 7 3188 59 3197
rect 7 3154 16 3188
rect 16 3154 50 3188
rect 50 3154 59 3188
rect 7 3145 59 3154
rect 1639 3188 1691 3197
rect 1639 3154 1648 3188
rect 1648 3154 1682 3188
rect 1682 3154 1691 3188
rect 1639 3145 1691 3154
rect 3271 3188 3323 3197
rect 3271 3154 3280 3188
rect 3280 3154 3314 3188
rect 3314 3154 3323 3188
rect 3271 3145 3323 3154
rect 4903 3188 4955 3197
rect 4903 3154 4912 3188
rect 4912 3154 4946 3188
rect 4946 3154 4955 3188
rect 4903 3145 4955 3154
rect 6535 3188 6587 3197
rect 6535 3154 6544 3188
rect 6544 3154 6578 3188
rect 6578 3154 6587 3188
rect 6535 3145 6587 3154
rect 8167 3188 8219 3197
rect 8167 3154 8176 3188
rect 8176 3154 8210 3188
rect 8210 3154 8219 3188
rect 8167 3145 8219 3154
rect 9799 3188 9851 3197
rect 9799 3154 9808 3188
rect 9808 3154 9842 3188
rect 9842 3154 9851 3188
rect 9799 3145 9851 3154
rect 7 2984 59 2993
rect 7 2950 16 2984
rect 16 2950 50 2984
rect 50 2950 59 2984
rect 7 2941 59 2950
rect 1639 2984 1691 2993
rect 1639 2950 1648 2984
rect 1648 2950 1682 2984
rect 1682 2950 1691 2984
rect 1639 2941 1691 2950
rect 3271 2984 3323 2993
rect 3271 2950 3280 2984
rect 3280 2950 3314 2984
rect 3314 2950 3323 2984
rect 3271 2941 3323 2950
rect 4903 2984 4955 2993
rect 4903 2950 4912 2984
rect 4912 2950 4946 2984
rect 4946 2950 4955 2984
rect 4903 2941 4955 2950
rect 6535 2984 6587 2993
rect 6535 2950 6544 2984
rect 6544 2950 6578 2984
rect 6578 2950 6587 2984
rect 6535 2941 6587 2950
rect 8167 2984 8219 2993
rect 8167 2950 8176 2984
rect 8176 2950 8210 2984
rect 8210 2950 8219 2984
rect 8167 2941 8219 2950
rect 9799 2984 9851 2993
rect 9799 2950 9808 2984
rect 9808 2950 9842 2984
rect 9842 2950 9851 2984
rect 9799 2941 9851 2950
rect 7 2780 59 2789
rect 7 2746 16 2780
rect 16 2746 50 2780
rect 50 2746 59 2780
rect 7 2737 59 2746
rect 1639 2780 1691 2789
rect 1639 2746 1648 2780
rect 1648 2746 1682 2780
rect 1682 2746 1691 2780
rect 1639 2737 1691 2746
rect 3271 2780 3323 2789
rect 3271 2746 3280 2780
rect 3280 2746 3314 2780
rect 3314 2746 3323 2780
rect 3271 2737 3323 2746
rect 4903 2780 4955 2789
rect 4903 2746 4912 2780
rect 4912 2746 4946 2780
rect 4946 2746 4955 2780
rect 4903 2737 4955 2746
rect 6535 2780 6587 2789
rect 6535 2746 6544 2780
rect 6544 2746 6578 2780
rect 6578 2746 6587 2780
rect 6535 2737 6587 2746
rect 8167 2780 8219 2789
rect 8167 2746 8176 2780
rect 8176 2746 8210 2780
rect 8210 2746 8219 2780
rect 8167 2737 8219 2746
rect 9799 2780 9851 2789
rect 9799 2746 9808 2780
rect 9808 2746 9842 2780
rect 9842 2746 9851 2780
rect 9799 2737 9851 2746
rect 218 2626 270 2635
rect 218 2592 227 2626
rect 227 2592 261 2626
rect 261 2592 270 2626
rect 218 2583 270 2592
rect 422 2626 474 2635
rect 422 2592 431 2626
rect 431 2592 465 2626
rect 465 2592 474 2626
rect 422 2583 474 2592
rect 626 2626 678 2635
rect 626 2592 635 2626
rect 635 2592 669 2626
rect 669 2592 678 2626
rect 626 2583 678 2592
rect 830 2626 882 2635
rect 830 2592 839 2626
rect 839 2592 873 2626
rect 873 2592 882 2626
rect 830 2583 882 2592
rect 1034 2626 1086 2635
rect 1034 2592 1043 2626
rect 1043 2592 1077 2626
rect 1077 2592 1086 2626
rect 1034 2583 1086 2592
rect 1238 2626 1290 2635
rect 1238 2592 1247 2626
rect 1247 2592 1281 2626
rect 1281 2592 1290 2626
rect 1238 2583 1290 2592
rect 1442 2626 1494 2635
rect 1442 2592 1451 2626
rect 1451 2592 1485 2626
rect 1485 2592 1494 2626
rect 1442 2583 1494 2592
rect 1646 2626 1698 2635
rect 1646 2592 1655 2626
rect 1655 2592 1689 2626
rect 1689 2592 1698 2626
rect 1646 2583 1698 2592
rect 1850 2626 1902 2635
rect 1850 2592 1859 2626
rect 1859 2592 1893 2626
rect 1893 2592 1902 2626
rect 1850 2583 1902 2592
rect 2054 2626 2106 2635
rect 2054 2592 2063 2626
rect 2063 2592 2097 2626
rect 2097 2592 2106 2626
rect 2054 2583 2106 2592
rect 2258 2626 2310 2635
rect 2258 2592 2267 2626
rect 2267 2592 2301 2626
rect 2301 2592 2310 2626
rect 2258 2583 2310 2592
rect 2462 2626 2514 2635
rect 2462 2592 2471 2626
rect 2471 2592 2505 2626
rect 2505 2592 2514 2626
rect 2462 2583 2514 2592
rect 2666 2626 2718 2635
rect 2666 2592 2675 2626
rect 2675 2592 2709 2626
rect 2709 2592 2718 2626
rect 2666 2583 2718 2592
rect 2870 2626 2922 2635
rect 2870 2592 2879 2626
rect 2879 2592 2913 2626
rect 2913 2592 2922 2626
rect 2870 2583 2922 2592
rect 3074 2626 3126 2635
rect 3074 2592 3083 2626
rect 3083 2592 3117 2626
rect 3117 2592 3126 2626
rect 3074 2583 3126 2592
rect 3278 2626 3330 2635
rect 3278 2592 3287 2626
rect 3287 2592 3321 2626
rect 3321 2592 3330 2626
rect 3278 2583 3330 2592
rect 3482 2626 3534 2635
rect 3482 2592 3491 2626
rect 3491 2592 3525 2626
rect 3525 2592 3534 2626
rect 3482 2583 3534 2592
rect 3686 2626 3738 2635
rect 3686 2592 3695 2626
rect 3695 2592 3729 2626
rect 3729 2592 3738 2626
rect 3686 2583 3738 2592
rect 3890 2626 3942 2635
rect 3890 2592 3899 2626
rect 3899 2592 3933 2626
rect 3933 2592 3942 2626
rect 3890 2583 3942 2592
rect 4094 2626 4146 2635
rect 4094 2592 4103 2626
rect 4103 2592 4137 2626
rect 4137 2592 4146 2626
rect 4094 2583 4146 2592
rect 4298 2626 4350 2635
rect 4298 2592 4307 2626
rect 4307 2592 4341 2626
rect 4341 2592 4350 2626
rect 4298 2583 4350 2592
rect 4502 2626 4554 2635
rect 4502 2592 4511 2626
rect 4511 2592 4545 2626
rect 4545 2592 4554 2626
rect 4502 2583 4554 2592
rect 4706 2626 4758 2635
rect 4706 2592 4715 2626
rect 4715 2592 4749 2626
rect 4749 2592 4758 2626
rect 4706 2583 4758 2592
rect 4910 2626 4962 2635
rect 4910 2592 4919 2626
rect 4919 2592 4953 2626
rect 4953 2592 4962 2626
rect 4910 2583 4962 2592
rect 5114 2626 5166 2635
rect 5114 2592 5123 2626
rect 5123 2592 5157 2626
rect 5157 2592 5166 2626
rect 5114 2583 5166 2592
rect 5318 2626 5370 2635
rect 5318 2592 5327 2626
rect 5327 2592 5361 2626
rect 5361 2592 5370 2626
rect 5318 2583 5370 2592
rect 5522 2626 5574 2635
rect 5522 2592 5531 2626
rect 5531 2592 5565 2626
rect 5565 2592 5574 2626
rect 5522 2583 5574 2592
rect 5726 2626 5778 2635
rect 5726 2592 5735 2626
rect 5735 2592 5769 2626
rect 5769 2592 5778 2626
rect 5726 2583 5778 2592
rect 5930 2626 5982 2635
rect 5930 2592 5939 2626
rect 5939 2592 5973 2626
rect 5973 2592 5982 2626
rect 5930 2583 5982 2592
rect 6134 2626 6186 2635
rect 6134 2592 6143 2626
rect 6143 2592 6177 2626
rect 6177 2592 6186 2626
rect 6134 2583 6186 2592
rect 6338 2626 6390 2635
rect 6338 2592 6347 2626
rect 6347 2592 6381 2626
rect 6381 2592 6390 2626
rect 6338 2583 6390 2592
rect 6542 2626 6594 2635
rect 6542 2592 6551 2626
rect 6551 2592 6585 2626
rect 6585 2592 6594 2626
rect 6542 2583 6594 2592
rect 6746 2626 6798 2635
rect 6746 2592 6755 2626
rect 6755 2592 6789 2626
rect 6789 2592 6798 2626
rect 6746 2583 6798 2592
rect 6950 2626 7002 2635
rect 6950 2592 6959 2626
rect 6959 2592 6993 2626
rect 6993 2592 7002 2626
rect 6950 2583 7002 2592
rect 7154 2626 7206 2635
rect 7154 2592 7163 2626
rect 7163 2592 7197 2626
rect 7197 2592 7206 2626
rect 7154 2583 7206 2592
rect 7358 2626 7410 2635
rect 7358 2592 7367 2626
rect 7367 2592 7401 2626
rect 7401 2592 7410 2626
rect 7358 2583 7410 2592
rect 7562 2626 7614 2635
rect 7562 2592 7571 2626
rect 7571 2592 7605 2626
rect 7605 2592 7614 2626
rect 7562 2583 7614 2592
rect 7766 2626 7818 2635
rect 7766 2592 7775 2626
rect 7775 2592 7809 2626
rect 7809 2592 7818 2626
rect 7766 2583 7818 2592
rect 7970 2626 8022 2635
rect 7970 2592 7979 2626
rect 7979 2592 8013 2626
rect 8013 2592 8022 2626
rect 7970 2583 8022 2592
rect 8174 2626 8226 2635
rect 8174 2592 8183 2626
rect 8183 2592 8217 2626
rect 8217 2592 8226 2626
rect 8174 2583 8226 2592
rect 8378 2626 8430 2635
rect 8378 2592 8387 2626
rect 8387 2592 8421 2626
rect 8421 2592 8430 2626
rect 8378 2583 8430 2592
rect 8582 2626 8634 2635
rect 8582 2592 8591 2626
rect 8591 2592 8625 2626
rect 8625 2592 8634 2626
rect 8582 2583 8634 2592
rect 8786 2626 8838 2635
rect 8786 2592 8795 2626
rect 8795 2592 8829 2626
rect 8829 2592 8838 2626
rect 8786 2583 8838 2592
rect 8990 2626 9042 2635
rect 8990 2592 8999 2626
rect 8999 2592 9033 2626
rect 9033 2592 9042 2626
rect 8990 2583 9042 2592
rect 9194 2626 9246 2635
rect 9194 2592 9203 2626
rect 9203 2592 9237 2626
rect 9237 2592 9246 2626
rect 9194 2583 9246 2592
rect 9398 2626 9450 2635
rect 9398 2592 9407 2626
rect 9407 2592 9441 2626
rect 9441 2592 9450 2626
rect 9398 2583 9450 2592
rect 9602 2626 9654 2635
rect 9602 2592 9611 2626
rect 9611 2592 9645 2626
rect 9645 2592 9654 2626
rect 9602 2583 9654 2592
rect 9820 2626 9872 2635
rect 9820 2592 9829 2626
rect 9829 2592 9863 2626
rect 9863 2592 9872 2626
rect 9820 2583 9872 2592
rect 7 2472 59 2481
rect 7 2438 16 2472
rect 16 2438 50 2472
rect 50 2438 59 2472
rect 7 2429 59 2438
rect 1639 2472 1691 2481
rect 1639 2438 1648 2472
rect 1648 2438 1682 2472
rect 1682 2438 1691 2472
rect 1639 2429 1691 2438
rect 3271 2472 3323 2481
rect 3271 2438 3280 2472
rect 3280 2438 3314 2472
rect 3314 2438 3323 2472
rect 3271 2429 3323 2438
rect 4903 2472 4955 2481
rect 4903 2438 4912 2472
rect 4912 2438 4946 2472
rect 4946 2438 4955 2472
rect 4903 2429 4955 2438
rect 6535 2472 6587 2481
rect 6535 2438 6544 2472
rect 6544 2438 6578 2472
rect 6578 2438 6587 2472
rect 6535 2429 6587 2438
rect 8167 2472 8219 2481
rect 8167 2438 8176 2472
rect 8176 2438 8210 2472
rect 8210 2438 8219 2472
rect 8167 2429 8219 2438
rect 9799 2472 9851 2481
rect 9799 2438 9808 2472
rect 9808 2438 9842 2472
rect 9842 2438 9851 2472
rect 9799 2429 9851 2438
rect 7 2268 59 2277
rect 7 2234 16 2268
rect 16 2234 50 2268
rect 50 2234 59 2268
rect 7 2225 59 2234
rect 1639 2268 1691 2277
rect 1639 2234 1648 2268
rect 1648 2234 1682 2268
rect 1682 2234 1691 2268
rect 1639 2225 1691 2234
rect 3271 2268 3323 2277
rect 3271 2234 3280 2268
rect 3280 2234 3314 2268
rect 3314 2234 3323 2268
rect 3271 2225 3323 2234
rect 4903 2268 4955 2277
rect 4903 2234 4912 2268
rect 4912 2234 4946 2268
rect 4946 2234 4955 2268
rect 4903 2225 4955 2234
rect 6535 2268 6587 2277
rect 6535 2234 6544 2268
rect 6544 2234 6578 2268
rect 6578 2234 6587 2268
rect 6535 2225 6587 2234
rect 8167 2268 8219 2277
rect 8167 2234 8176 2268
rect 8176 2234 8210 2268
rect 8210 2234 8219 2268
rect 8167 2225 8219 2234
rect 9799 2268 9851 2277
rect 9799 2234 9808 2268
rect 9808 2234 9842 2268
rect 9842 2234 9851 2268
rect 9799 2225 9851 2234
rect 7 2064 59 2073
rect 7 2030 16 2064
rect 16 2030 50 2064
rect 50 2030 59 2064
rect 7 2021 59 2030
rect 1639 2064 1691 2073
rect 1639 2030 1648 2064
rect 1648 2030 1682 2064
rect 1682 2030 1691 2064
rect 1639 2021 1691 2030
rect 3271 2064 3323 2073
rect 3271 2030 3280 2064
rect 3280 2030 3314 2064
rect 3314 2030 3323 2064
rect 3271 2021 3323 2030
rect 4903 2064 4955 2073
rect 4903 2030 4912 2064
rect 4912 2030 4946 2064
rect 4946 2030 4955 2064
rect 4903 2021 4955 2030
rect 6535 2064 6587 2073
rect 6535 2030 6544 2064
rect 6544 2030 6578 2064
rect 6578 2030 6587 2064
rect 6535 2021 6587 2030
rect 8167 2064 8219 2073
rect 8167 2030 8176 2064
rect 8176 2030 8210 2064
rect 8210 2030 8219 2064
rect 8167 2021 8219 2030
rect 9799 2064 9851 2073
rect 9799 2030 9808 2064
rect 9808 2030 9842 2064
rect 9842 2030 9851 2064
rect 9799 2021 9851 2030
rect 7 1860 59 1869
rect 7 1826 16 1860
rect 16 1826 50 1860
rect 50 1826 59 1860
rect 7 1817 59 1826
rect 1639 1860 1691 1869
rect 1639 1826 1648 1860
rect 1648 1826 1682 1860
rect 1682 1826 1691 1860
rect 1639 1817 1691 1826
rect 3271 1860 3323 1869
rect 3271 1826 3280 1860
rect 3280 1826 3314 1860
rect 3314 1826 3323 1860
rect 3271 1817 3323 1826
rect 4903 1860 4955 1869
rect 4903 1826 4912 1860
rect 4912 1826 4946 1860
rect 4946 1826 4955 1860
rect 4903 1817 4955 1826
rect 6535 1860 6587 1869
rect 6535 1826 6544 1860
rect 6544 1826 6578 1860
rect 6578 1826 6587 1860
rect 6535 1817 6587 1826
rect 8167 1860 8219 1869
rect 8167 1826 8176 1860
rect 8176 1826 8210 1860
rect 8210 1826 8219 1860
rect 8167 1817 8219 1826
rect 9799 1860 9851 1869
rect 9799 1826 9808 1860
rect 9808 1826 9842 1860
rect 9842 1826 9851 1860
rect 9799 1817 9851 1826
rect 7 1656 59 1665
rect 7 1622 16 1656
rect 16 1622 50 1656
rect 50 1622 59 1656
rect 7 1613 59 1622
rect 1639 1656 1691 1665
rect 1639 1622 1648 1656
rect 1648 1622 1682 1656
rect 1682 1622 1691 1656
rect 1639 1613 1691 1622
rect 3271 1656 3323 1665
rect 3271 1622 3280 1656
rect 3280 1622 3314 1656
rect 3314 1622 3323 1656
rect 3271 1613 3323 1622
rect 4903 1656 4955 1665
rect 4903 1622 4912 1656
rect 4912 1622 4946 1656
rect 4946 1622 4955 1656
rect 4903 1613 4955 1622
rect 6535 1656 6587 1665
rect 6535 1622 6544 1656
rect 6544 1622 6578 1656
rect 6578 1622 6587 1656
rect 6535 1613 6587 1622
rect 8167 1656 8219 1665
rect 8167 1622 8176 1656
rect 8176 1622 8210 1656
rect 8210 1622 8219 1656
rect 8167 1613 8219 1622
rect 9799 1656 9851 1665
rect 9799 1622 9808 1656
rect 9808 1622 9842 1656
rect 9842 1622 9851 1656
rect 9799 1613 9851 1622
rect 7 1452 59 1461
rect 7 1418 16 1452
rect 16 1418 50 1452
rect 50 1418 59 1452
rect 7 1409 59 1418
rect 1639 1452 1691 1461
rect 1639 1418 1648 1452
rect 1648 1418 1682 1452
rect 1682 1418 1691 1452
rect 1639 1409 1691 1418
rect 3271 1452 3323 1461
rect 3271 1418 3280 1452
rect 3280 1418 3314 1452
rect 3314 1418 3323 1452
rect 3271 1409 3323 1418
rect 4903 1452 4955 1461
rect 4903 1418 4912 1452
rect 4912 1418 4946 1452
rect 4946 1418 4955 1452
rect 4903 1409 4955 1418
rect 6535 1452 6587 1461
rect 6535 1418 6544 1452
rect 6544 1418 6578 1452
rect 6578 1418 6587 1452
rect 6535 1409 6587 1418
rect 8167 1452 8219 1461
rect 8167 1418 8176 1452
rect 8176 1418 8210 1452
rect 8210 1418 8219 1452
rect 8167 1409 8219 1418
rect 9799 1452 9851 1461
rect 9799 1418 9808 1452
rect 9808 1418 9842 1452
rect 9842 1418 9851 1452
rect 9799 1409 9851 1418
rect 7 1248 59 1257
rect 7 1214 16 1248
rect 16 1214 50 1248
rect 50 1214 59 1248
rect 7 1205 59 1214
rect 1639 1248 1691 1257
rect 1639 1214 1648 1248
rect 1648 1214 1682 1248
rect 1682 1214 1691 1248
rect 1639 1205 1691 1214
rect 3271 1248 3323 1257
rect 3271 1214 3280 1248
rect 3280 1214 3314 1248
rect 3314 1214 3323 1248
rect 3271 1205 3323 1214
rect 4903 1248 4955 1257
rect 4903 1214 4912 1248
rect 4912 1214 4946 1248
rect 4946 1214 4955 1248
rect 4903 1205 4955 1214
rect 6535 1248 6587 1257
rect 6535 1214 6544 1248
rect 6544 1214 6578 1248
rect 6578 1214 6587 1248
rect 6535 1205 6587 1214
rect 8167 1248 8219 1257
rect 8167 1214 8176 1248
rect 8176 1214 8210 1248
rect 8210 1214 8219 1248
rect 8167 1205 8219 1214
rect 9799 1248 9851 1257
rect 9799 1214 9808 1248
rect 9808 1214 9842 1248
rect 9842 1214 9851 1248
rect 9799 1205 9851 1214
rect 7 1044 59 1053
rect 7 1010 16 1044
rect 16 1010 50 1044
rect 50 1010 59 1044
rect 7 1001 59 1010
rect 1639 1044 1691 1053
rect 1639 1010 1648 1044
rect 1648 1010 1682 1044
rect 1682 1010 1691 1044
rect 1639 1001 1691 1010
rect 3271 1044 3323 1053
rect 3271 1010 3280 1044
rect 3280 1010 3314 1044
rect 3314 1010 3323 1044
rect 3271 1001 3323 1010
rect 4903 1044 4955 1053
rect 4903 1010 4912 1044
rect 4912 1010 4946 1044
rect 4946 1010 4955 1044
rect 4903 1001 4955 1010
rect 6535 1044 6587 1053
rect 6535 1010 6544 1044
rect 6544 1010 6578 1044
rect 6578 1010 6587 1044
rect 6535 1001 6587 1010
rect 8167 1044 8219 1053
rect 8167 1010 8176 1044
rect 8176 1010 8210 1044
rect 8210 1010 8219 1044
rect 8167 1001 8219 1010
rect 9799 1044 9851 1053
rect 9799 1010 9808 1044
rect 9808 1010 9842 1044
rect 9842 1010 9851 1044
rect 9799 1001 9851 1010
rect 218 890 270 899
rect 218 856 227 890
rect 227 856 261 890
rect 261 856 270 890
rect 218 847 270 856
rect 422 890 474 899
rect 422 856 431 890
rect 431 856 465 890
rect 465 856 474 890
rect 422 847 474 856
rect 626 890 678 899
rect 626 856 635 890
rect 635 856 669 890
rect 669 856 678 890
rect 626 847 678 856
rect 830 890 882 899
rect 830 856 839 890
rect 839 856 873 890
rect 873 856 882 890
rect 830 847 882 856
rect 1034 890 1086 899
rect 1034 856 1043 890
rect 1043 856 1077 890
rect 1077 856 1086 890
rect 1034 847 1086 856
rect 1238 890 1290 899
rect 1238 856 1247 890
rect 1247 856 1281 890
rect 1281 856 1290 890
rect 1238 847 1290 856
rect 1442 890 1494 899
rect 1442 856 1451 890
rect 1451 856 1485 890
rect 1485 856 1494 890
rect 1442 847 1494 856
rect 1646 890 1698 899
rect 1646 856 1655 890
rect 1655 856 1689 890
rect 1689 856 1698 890
rect 1646 847 1698 856
rect 1850 890 1902 899
rect 1850 856 1859 890
rect 1859 856 1893 890
rect 1893 856 1902 890
rect 1850 847 1902 856
rect 2054 890 2106 899
rect 2054 856 2063 890
rect 2063 856 2097 890
rect 2097 856 2106 890
rect 2054 847 2106 856
rect 2258 890 2310 899
rect 2258 856 2267 890
rect 2267 856 2301 890
rect 2301 856 2310 890
rect 2258 847 2310 856
rect 2462 890 2514 899
rect 2462 856 2471 890
rect 2471 856 2505 890
rect 2505 856 2514 890
rect 2462 847 2514 856
rect 2666 890 2718 899
rect 2666 856 2675 890
rect 2675 856 2709 890
rect 2709 856 2718 890
rect 2666 847 2718 856
rect 2870 890 2922 899
rect 2870 856 2879 890
rect 2879 856 2913 890
rect 2913 856 2922 890
rect 2870 847 2922 856
rect 3074 890 3126 899
rect 3074 856 3083 890
rect 3083 856 3117 890
rect 3117 856 3126 890
rect 3074 847 3126 856
rect 3278 890 3330 899
rect 3278 856 3287 890
rect 3287 856 3321 890
rect 3321 856 3330 890
rect 3278 847 3330 856
rect 3482 890 3534 899
rect 3482 856 3491 890
rect 3491 856 3525 890
rect 3525 856 3534 890
rect 3482 847 3534 856
rect 3686 890 3738 899
rect 3686 856 3695 890
rect 3695 856 3729 890
rect 3729 856 3738 890
rect 3686 847 3738 856
rect 3890 890 3942 899
rect 3890 856 3899 890
rect 3899 856 3933 890
rect 3933 856 3942 890
rect 3890 847 3942 856
rect 4094 890 4146 899
rect 4094 856 4103 890
rect 4103 856 4137 890
rect 4137 856 4146 890
rect 4094 847 4146 856
rect 4298 890 4350 899
rect 4298 856 4307 890
rect 4307 856 4341 890
rect 4341 856 4350 890
rect 4298 847 4350 856
rect 4502 890 4554 899
rect 4502 856 4511 890
rect 4511 856 4545 890
rect 4545 856 4554 890
rect 4502 847 4554 856
rect 4706 890 4758 899
rect 4706 856 4715 890
rect 4715 856 4749 890
rect 4749 856 4758 890
rect 4706 847 4758 856
rect 4910 890 4962 899
rect 4910 856 4919 890
rect 4919 856 4953 890
rect 4953 856 4962 890
rect 4910 847 4962 856
rect 5114 890 5166 899
rect 5114 856 5123 890
rect 5123 856 5157 890
rect 5157 856 5166 890
rect 5114 847 5166 856
rect 5318 890 5370 899
rect 5318 856 5327 890
rect 5327 856 5361 890
rect 5361 856 5370 890
rect 5318 847 5370 856
rect 5522 890 5574 899
rect 5522 856 5531 890
rect 5531 856 5565 890
rect 5565 856 5574 890
rect 5522 847 5574 856
rect 5726 890 5778 899
rect 5726 856 5735 890
rect 5735 856 5769 890
rect 5769 856 5778 890
rect 5726 847 5778 856
rect 5930 890 5982 899
rect 5930 856 5939 890
rect 5939 856 5973 890
rect 5973 856 5982 890
rect 5930 847 5982 856
rect 6134 890 6186 899
rect 6134 856 6143 890
rect 6143 856 6177 890
rect 6177 856 6186 890
rect 6134 847 6186 856
rect 6338 890 6390 899
rect 6338 856 6347 890
rect 6347 856 6381 890
rect 6381 856 6390 890
rect 6338 847 6390 856
rect 6542 890 6594 899
rect 6542 856 6551 890
rect 6551 856 6585 890
rect 6585 856 6594 890
rect 6542 847 6594 856
rect 6746 890 6798 899
rect 6746 856 6755 890
rect 6755 856 6789 890
rect 6789 856 6798 890
rect 6746 847 6798 856
rect 6950 890 7002 899
rect 6950 856 6959 890
rect 6959 856 6993 890
rect 6993 856 7002 890
rect 6950 847 7002 856
rect 7154 890 7206 899
rect 7154 856 7163 890
rect 7163 856 7197 890
rect 7197 856 7206 890
rect 7154 847 7206 856
rect 7358 890 7410 899
rect 7358 856 7367 890
rect 7367 856 7401 890
rect 7401 856 7410 890
rect 7358 847 7410 856
rect 7562 890 7614 899
rect 7562 856 7571 890
rect 7571 856 7605 890
rect 7605 856 7614 890
rect 7562 847 7614 856
rect 7766 890 7818 899
rect 7766 856 7775 890
rect 7775 856 7809 890
rect 7809 856 7818 890
rect 7766 847 7818 856
rect 7970 890 8022 899
rect 7970 856 7979 890
rect 7979 856 8013 890
rect 8013 856 8022 890
rect 7970 847 8022 856
rect 8174 890 8226 899
rect 8174 856 8183 890
rect 8183 856 8217 890
rect 8217 856 8226 890
rect 8174 847 8226 856
rect 8378 890 8430 899
rect 8378 856 8387 890
rect 8387 856 8421 890
rect 8421 856 8430 890
rect 8378 847 8430 856
rect 8582 890 8634 899
rect 8582 856 8591 890
rect 8591 856 8625 890
rect 8625 856 8634 890
rect 8582 847 8634 856
rect 8786 890 8838 899
rect 8786 856 8795 890
rect 8795 856 8829 890
rect 8829 856 8838 890
rect 8786 847 8838 856
rect 8990 890 9042 899
rect 8990 856 8999 890
rect 8999 856 9033 890
rect 9033 856 9042 890
rect 8990 847 9042 856
rect 9194 890 9246 899
rect 9194 856 9203 890
rect 9203 856 9237 890
rect 9237 856 9246 890
rect 9194 847 9246 856
rect 9398 890 9450 899
rect 9398 856 9407 890
rect 9407 856 9441 890
rect 9441 856 9450 890
rect 9398 847 9450 856
rect 9602 890 9654 899
rect 9602 856 9611 890
rect 9611 856 9645 890
rect 9645 856 9654 890
rect 9602 847 9654 856
rect 9820 890 9872 899
rect 9820 856 9829 890
rect 9829 856 9863 890
rect 9863 856 9872 890
rect 9820 847 9872 856
<< metal2 >>
rect 7 10141 59 10147
rect 1 10094 7 10137
rect 1639 10141 1691 10147
rect 59 10129 65 10137
rect 1633 10129 1639 10137
rect 59 10101 1639 10129
rect 59 10094 65 10101
rect 1633 10094 1639 10101
rect 7 10083 59 10089
rect 3271 10141 3323 10147
rect 1691 10129 1697 10137
rect 3265 10129 3271 10137
rect 1691 10101 3271 10129
rect 1691 10094 1697 10101
rect 3265 10094 3271 10101
rect 1639 10083 1691 10089
rect 4903 10141 4955 10147
rect 3323 10129 3329 10137
rect 4897 10129 4903 10137
rect 3323 10101 4903 10129
rect 3323 10094 3329 10101
rect 4897 10094 4903 10101
rect 3271 10083 3323 10089
rect 6535 10141 6587 10147
rect 4955 10129 4961 10137
rect 6529 10129 6535 10137
rect 4955 10101 6535 10129
rect 4955 10094 4961 10101
rect 6529 10094 6535 10101
rect 4903 10083 4955 10089
rect 8167 10141 8219 10147
rect 6587 10129 6593 10137
rect 8161 10129 8167 10137
rect 6587 10101 8167 10129
rect 6587 10094 6593 10101
rect 8161 10094 8167 10101
rect 6535 10083 6587 10089
rect 9799 10141 9851 10147
rect 8219 10129 8225 10137
rect 9793 10129 9799 10137
rect 8219 10101 9799 10129
rect 8219 10094 8225 10101
rect 9793 10094 9799 10101
rect 8167 10083 8219 10089
rect 9851 10094 9857 10137
rect 9799 10083 9851 10089
rect 7 9937 59 9943
rect 1 9890 7 9933
rect 1639 9937 1691 9943
rect 59 9925 65 9933
rect 1633 9925 1639 9933
rect 59 9897 1639 9925
rect 59 9890 65 9897
rect 1633 9890 1639 9897
rect 7 9879 59 9885
rect 3271 9937 3323 9943
rect 1691 9925 1697 9933
rect 3265 9925 3271 9933
rect 1691 9897 3271 9925
rect 1691 9890 1697 9897
rect 3265 9890 3271 9897
rect 1639 9879 1691 9885
rect 4903 9937 4955 9943
rect 3323 9925 3329 9933
rect 4897 9925 4903 9933
rect 3323 9897 4903 9925
rect 3323 9890 3329 9897
rect 4897 9890 4903 9897
rect 3271 9879 3323 9885
rect 6535 9937 6587 9943
rect 4955 9925 4961 9933
rect 6529 9925 6535 9933
rect 4955 9897 6535 9925
rect 4955 9890 4961 9897
rect 6529 9890 6535 9897
rect 4903 9879 4955 9885
rect 8167 9937 8219 9943
rect 6587 9925 6593 9933
rect 8161 9925 8167 9933
rect 6587 9897 8167 9925
rect 6587 9890 6593 9897
rect 8161 9890 8167 9897
rect 6535 9879 6587 9885
rect 9799 9937 9851 9943
rect 8219 9925 8225 9933
rect 9793 9925 9799 9933
rect 8219 9897 9799 9925
rect 8219 9890 8225 9897
rect 9793 9890 9799 9897
rect 8167 9879 8219 9885
rect 9851 9890 9857 9933
rect 9799 9879 9851 9885
rect 7 9733 59 9739
rect 1 9686 7 9729
rect 1639 9733 1691 9739
rect 59 9721 65 9729
rect 1633 9721 1639 9729
rect 59 9693 1639 9721
rect 59 9686 65 9693
rect 1633 9686 1639 9693
rect 7 9675 59 9681
rect 3271 9733 3323 9739
rect 1691 9721 1697 9729
rect 3265 9721 3271 9729
rect 1691 9693 3271 9721
rect 1691 9686 1697 9693
rect 3265 9686 3271 9693
rect 1639 9675 1691 9681
rect 4903 9733 4955 9739
rect 3323 9721 3329 9729
rect 4897 9721 4903 9729
rect 3323 9693 4903 9721
rect 3323 9686 3329 9693
rect 4897 9686 4903 9693
rect 3271 9675 3323 9681
rect 6535 9733 6587 9739
rect 4955 9721 4961 9729
rect 6529 9721 6535 9729
rect 4955 9693 6535 9721
rect 4955 9686 4961 9693
rect 6529 9686 6535 9693
rect 4903 9675 4955 9681
rect 8167 9733 8219 9739
rect 6587 9721 6593 9729
rect 8161 9721 8167 9729
rect 6587 9693 8167 9721
rect 6587 9686 6593 9693
rect 8161 9686 8167 9693
rect 6535 9675 6587 9681
rect 9799 9733 9851 9739
rect 8219 9721 8225 9729
rect 9793 9721 9799 9729
rect 8219 9693 9799 9721
rect 8219 9686 8225 9693
rect 9793 9686 9799 9693
rect 8167 9675 8219 9681
rect 9851 9686 9857 9729
rect 9799 9675 9851 9681
rect 212 9527 218 9579
rect 270 9567 276 9579
rect 416 9567 422 9579
rect 270 9539 422 9567
rect 270 9527 276 9539
rect 416 9527 422 9539
rect 474 9567 480 9579
rect 620 9567 626 9579
rect 474 9539 626 9567
rect 474 9527 480 9539
rect 620 9527 626 9539
rect 678 9567 684 9579
rect 824 9567 830 9579
rect 678 9539 830 9567
rect 678 9527 684 9539
rect 824 9527 830 9539
rect 882 9567 888 9579
rect 1028 9567 1034 9579
rect 882 9539 1034 9567
rect 882 9527 888 9539
rect 1028 9527 1034 9539
rect 1086 9567 1092 9579
rect 1232 9567 1238 9579
rect 1086 9539 1238 9567
rect 1086 9527 1092 9539
rect 1232 9527 1238 9539
rect 1290 9567 1296 9579
rect 1436 9567 1442 9579
rect 1290 9539 1442 9567
rect 1290 9527 1296 9539
rect 1436 9527 1442 9539
rect 1494 9567 1500 9579
rect 1640 9567 1646 9579
rect 1494 9539 1646 9567
rect 1494 9527 1500 9539
rect 1640 9527 1646 9539
rect 1698 9567 1704 9579
rect 1844 9567 1850 9579
rect 1698 9539 1850 9567
rect 1698 9527 1704 9539
rect 1844 9527 1850 9539
rect 1902 9567 1908 9579
rect 2048 9567 2054 9579
rect 1902 9539 2054 9567
rect 1902 9527 1908 9539
rect 2048 9527 2054 9539
rect 2106 9567 2112 9579
rect 2252 9567 2258 9579
rect 2106 9539 2258 9567
rect 2106 9527 2112 9539
rect 2252 9527 2258 9539
rect 2310 9567 2316 9579
rect 2456 9567 2462 9579
rect 2310 9539 2462 9567
rect 2310 9527 2316 9539
rect 2456 9527 2462 9539
rect 2514 9567 2520 9579
rect 2660 9567 2666 9579
rect 2514 9539 2666 9567
rect 2514 9527 2520 9539
rect 2660 9527 2666 9539
rect 2718 9567 2724 9579
rect 2864 9567 2870 9579
rect 2718 9539 2870 9567
rect 2718 9527 2724 9539
rect 2864 9527 2870 9539
rect 2922 9567 2928 9579
rect 3068 9567 3074 9579
rect 2922 9539 3074 9567
rect 2922 9527 2928 9539
rect 3068 9527 3074 9539
rect 3126 9567 3132 9579
rect 3272 9567 3278 9579
rect 3126 9539 3278 9567
rect 3126 9527 3132 9539
rect 3272 9527 3278 9539
rect 3330 9567 3336 9579
rect 3476 9567 3482 9579
rect 3330 9539 3482 9567
rect 3330 9527 3336 9539
rect 3476 9527 3482 9539
rect 3534 9567 3540 9579
rect 3680 9567 3686 9579
rect 3534 9539 3686 9567
rect 3534 9527 3540 9539
rect 3680 9527 3686 9539
rect 3738 9567 3744 9579
rect 3884 9567 3890 9579
rect 3738 9539 3890 9567
rect 3738 9527 3744 9539
rect 3884 9527 3890 9539
rect 3942 9567 3948 9579
rect 4088 9567 4094 9579
rect 3942 9539 4094 9567
rect 3942 9527 3948 9539
rect 4088 9527 4094 9539
rect 4146 9567 4152 9579
rect 4292 9567 4298 9579
rect 4146 9539 4298 9567
rect 4146 9527 4152 9539
rect 4292 9527 4298 9539
rect 4350 9567 4356 9579
rect 4496 9567 4502 9579
rect 4350 9539 4502 9567
rect 4350 9527 4356 9539
rect 4496 9527 4502 9539
rect 4554 9567 4560 9579
rect 4700 9567 4706 9579
rect 4554 9539 4706 9567
rect 4554 9527 4560 9539
rect 4700 9527 4706 9539
rect 4758 9567 4764 9579
rect 4904 9567 4910 9579
rect 4758 9539 4910 9567
rect 4758 9527 4764 9539
rect 4904 9527 4910 9539
rect 4962 9567 4968 9579
rect 5108 9567 5114 9579
rect 4962 9539 5114 9567
rect 4962 9527 4968 9539
rect 5108 9527 5114 9539
rect 5166 9567 5172 9579
rect 5312 9567 5318 9579
rect 5166 9539 5318 9567
rect 5166 9527 5172 9539
rect 5312 9527 5318 9539
rect 5370 9567 5376 9579
rect 5516 9567 5522 9579
rect 5370 9539 5522 9567
rect 5370 9527 5376 9539
rect 5516 9527 5522 9539
rect 5574 9567 5580 9579
rect 5720 9567 5726 9579
rect 5574 9539 5726 9567
rect 5574 9527 5580 9539
rect 5720 9527 5726 9539
rect 5778 9567 5784 9579
rect 5924 9567 5930 9579
rect 5778 9539 5930 9567
rect 5778 9527 5784 9539
rect 5924 9527 5930 9539
rect 5982 9567 5988 9579
rect 6128 9567 6134 9579
rect 5982 9539 6134 9567
rect 5982 9527 5988 9539
rect 6128 9527 6134 9539
rect 6186 9567 6192 9579
rect 6332 9567 6338 9579
rect 6186 9539 6338 9567
rect 6186 9527 6192 9539
rect 6332 9527 6338 9539
rect 6390 9567 6396 9579
rect 6536 9567 6542 9579
rect 6390 9539 6542 9567
rect 6390 9527 6396 9539
rect 6536 9527 6542 9539
rect 6594 9567 6600 9579
rect 6740 9567 6746 9579
rect 6594 9539 6746 9567
rect 6594 9527 6600 9539
rect 6740 9527 6746 9539
rect 6798 9567 6804 9579
rect 6944 9567 6950 9579
rect 6798 9539 6950 9567
rect 6798 9527 6804 9539
rect 6944 9527 6950 9539
rect 7002 9567 7008 9579
rect 7148 9567 7154 9579
rect 7002 9539 7154 9567
rect 7002 9527 7008 9539
rect 7148 9527 7154 9539
rect 7206 9567 7212 9579
rect 7352 9567 7358 9579
rect 7206 9539 7358 9567
rect 7206 9527 7212 9539
rect 7352 9527 7358 9539
rect 7410 9567 7416 9579
rect 7556 9567 7562 9579
rect 7410 9539 7562 9567
rect 7410 9527 7416 9539
rect 7556 9527 7562 9539
rect 7614 9567 7620 9579
rect 7760 9567 7766 9579
rect 7614 9539 7766 9567
rect 7614 9527 7620 9539
rect 7760 9527 7766 9539
rect 7818 9567 7824 9579
rect 7964 9567 7970 9579
rect 7818 9539 7970 9567
rect 7818 9527 7824 9539
rect 7964 9527 7970 9539
rect 8022 9567 8028 9579
rect 8168 9567 8174 9579
rect 8022 9539 8174 9567
rect 8022 9527 8028 9539
rect 8168 9527 8174 9539
rect 8226 9567 8232 9579
rect 8372 9567 8378 9579
rect 8226 9539 8378 9567
rect 8226 9527 8232 9539
rect 8372 9527 8378 9539
rect 8430 9567 8436 9579
rect 8576 9567 8582 9579
rect 8430 9539 8582 9567
rect 8430 9527 8436 9539
rect 8576 9527 8582 9539
rect 8634 9567 8640 9579
rect 8780 9567 8786 9579
rect 8634 9539 8786 9567
rect 8634 9527 8640 9539
rect 8780 9527 8786 9539
rect 8838 9567 8844 9579
rect 8984 9567 8990 9579
rect 8838 9539 8990 9567
rect 8838 9527 8844 9539
rect 8984 9527 8990 9539
rect 9042 9567 9048 9579
rect 9188 9567 9194 9579
rect 9042 9539 9194 9567
rect 9042 9527 9048 9539
rect 9188 9527 9194 9539
rect 9246 9567 9252 9579
rect 9392 9567 9398 9579
rect 9246 9539 9398 9567
rect 9246 9527 9252 9539
rect 9392 9527 9398 9539
rect 9450 9567 9456 9579
rect 9596 9567 9602 9579
rect 9450 9539 9602 9567
rect 9450 9527 9456 9539
rect 9596 9527 9602 9539
rect 9654 9567 9660 9579
rect 9814 9567 9820 9579
rect 9654 9539 9820 9567
rect 9654 9527 9660 9539
rect 9814 9527 9820 9539
rect 9872 9527 9878 9579
rect 7 9425 59 9431
rect 1 9378 7 9421
rect 1639 9425 1691 9431
rect 59 9413 65 9421
rect 1633 9413 1639 9421
rect 59 9385 1639 9413
rect 59 9378 65 9385
rect 1633 9378 1639 9385
rect 7 9367 59 9373
rect 3271 9425 3323 9431
rect 1691 9413 1697 9421
rect 3265 9413 3271 9421
rect 1691 9385 3271 9413
rect 1691 9378 1697 9385
rect 3265 9378 3271 9385
rect 1639 9367 1691 9373
rect 4903 9425 4955 9431
rect 3323 9413 3329 9421
rect 4897 9413 4903 9421
rect 3323 9385 4903 9413
rect 3323 9378 3329 9385
rect 4897 9378 4903 9385
rect 3271 9367 3323 9373
rect 6535 9425 6587 9431
rect 4955 9413 4961 9421
rect 6529 9413 6535 9421
rect 4955 9385 6535 9413
rect 4955 9378 4961 9385
rect 6529 9378 6535 9385
rect 4903 9367 4955 9373
rect 8167 9425 8219 9431
rect 6587 9413 6593 9421
rect 8161 9413 8167 9421
rect 6587 9385 8167 9413
rect 6587 9378 6593 9385
rect 8161 9378 8167 9385
rect 6535 9367 6587 9373
rect 9799 9425 9851 9431
rect 8219 9413 8225 9421
rect 9793 9413 9799 9421
rect 8219 9385 9799 9413
rect 8219 9378 8225 9385
rect 9793 9378 9799 9385
rect 8167 9367 8219 9373
rect 9851 9378 9857 9421
rect 9799 9367 9851 9373
rect 7 9221 59 9227
rect 1 9174 7 9217
rect 1639 9221 1691 9227
rect 59 9209 65 9217
rect 1633 9209 1639 9217
rect 59 9181 1639 9209
rect 59 9174 65 9181
rect 1633 9174 1639 9181
rect 7 9163 59 9169
rect 3271 9221 3323 9227
rect 1691 9209 1697 9217
rect 3265 9209 3271 9217
rect 1691 9181 3271 9209
rect 1691 9174 1697 9181
rect 3265 9174 3271 9181
rect 1639 9163 1691 9169
rect 4903 9221 4955 9227
rect 3323 9209 3329 9217
rect 4897 9209 4903 9217
rect 3323 9181 4903 9209
rect 3323 9174 3329 9181
rect 4897 9174 4903 9181
rect 3271 9163 3323 9169
rect 6535 9221 6587 9227
rect 4955 9209 4961 9217
rect 6529 9209 6535 9217
rect 4955 9181 6535 9209
rect 4955 9174 4961 9181
rect 6529 9174 6535 9181
rect 4903 9163 4955 9169
rect 8167 9221 8219 9227
rect 6587 9209 6593 9217
rect 8161 9209 8167 9217
rect 6587 9181 8167 9209
rect 6587 9174 6593 9181
rect 8161 9174 8167 9181
rect 6535 9163 6587 9169
rect 9799 9221 9851 9227
rect 8219 9209 8225 9217
rect 9793 9209 9799 9217
rect 8219 9181 9799 9209
rect 8219 9174 8225 9181
rect 9793 9174 9799 9181
rect 8167 9163 8219 9169
rect 9851 9174 9857 9217
rect 9799 9163 9851 9169
rect 7 9017 59 9023
rect 1 8970 7 9013
rect 1639 9017 1691 9023
rect 59 9005 65 9013
rect 1633 9005 1639 9013
rect 59 8977 1639 9005
rect 59 8970 65 8977
rect 1633 8970 1639 8977
rect 7 8959 59 8965
rect 3271 9017 3323 9023
rect 1691 9005 1697 9013
rect 3265 9005 3271 9013
rect 1691 8977 3271 9005
rect 1691 8970 1697 8977
rect 3265 8970 3271 8977
rect 1639 8959 1691 8965
rect 4903 9017 4955 9023
rect 3323 9005 3329 9013
rect 4897 9005 4903 9013
rect 3323 8977 4903 9005
rect 3323 8970 3329 8977
rect 4897 8970 4903 8977
rect 3271 8959 3323 8965
rect 6535 9017 6587 9023
rect 4955 9005 4961 9013
rect 6529 9005 6535 9013
rect 4955 8977 6535 9005
rect 4955 8970 4961 8977
rect 6529 8970 6535 8977
rect 4903 8959 4955 8965
rect 8167 9017 8219 9023
rect 6587 9005 6593 9013
rect 8161 9005 8167 9013
rect 6587 8977 8167 9005
rect 6587 8970 6593 8977
rect 8161 8970 8167 8977
rect 6535 8959 6587 8965
rect 9799 9017 9851 9023
rect 8219 9005 8225 9013
rect 9793 9005 9799 9013
rect 8219 8977 9799 9005
rect 8219 8970 8225 8977
rect 9793 8970 9799 8977
rect 8167 8959 8219 8965
rect 9851 8970 9857 9013
rect 9799 8959 9851 8965
rect 7 8813 59 8819
rect 1 8766 7 8809
rect 1639 8813 1691 8819
rect 59 8801 65 8809
rect 1633 8801 1639 8809
rect 59 8773 1639 8801
rect 59 8766 65 8773
rect 1633 8766 1639 8773
rect 7 8755 59 8761
rect 3271 8813 3323 8819
rect 1691 8801 1697 8809
rect 3265 8801 3271 8809
rect 1691 8773 3271 8801
rect 1691 8766 1697 8773
rect 3265 8766 3271 8773
rect 1639 8755 1691 8761
rect 4903 8813 4955 8819
rect 3323 8801 3329 8809
rect 4897 8801 4903 8809
rect 3323 8773 4903 8801
rect 3323 8766 3329 8773
rect 4897 8766 4903 8773
rect 3271 8755 3323 8761
rect 6535 8813 6587 8819
rect 4955 8801 4961 8809
rect 6529 8801 6535 8809
rect 4955 8773 6535 8801
rect 4955 8766 4961 8773
rect 6529 8766 6535 8773
rect 4903 8755 4955 8761
rect 8167 8813 8219 8819
rect 6587 8801 6593 8809
rect 8161 8801 8167 8809
rect 6587 8773 8167 8801
rect 6587 8766 6593 8773
rect 8161 8766 8167 8773
rect 6535 8755 6587 8761
rect 9799 8813 9851 8819
rect 8219 8801 8225 8809
rect 9793 8801 9799 8809
rect 8219 8773 9799 8801
rect 8219 8766 8225 8773
rect 9793 8766 9799 8773
rect 8167 8755 8219 8761
rect 9851 8766 9857 8809
rect 9799 8755 9851 8761
rect 7 8609 59 8615
rect 1 8562 7 8605
rect 1639 8609 1691 8615
rect 59 8597 65 8605
rect 1633 8597 1639 8605
rect 59 8569 1639 8597
rect 59 8562 65 8569
rect 1633 8562 1639 8569
rect 7 8551 59 8557
rect 3271 8609 3323 8615
rect 1691 8597 1697 8605
rect 3265 8597 3271 8605
rect 1691 8569 3271 8597
rect 1691 8562 1697 8569
rect 3265 8562 3271 8569
rect 1639 8551 1691 8557
rect 4903 8609 4955 8615
rect 3323 8597 3329 8605
rect 4897 8597 4903 8605
rect 3323 8569 4903 8597
rect 3323 8562 3329 8569
rect 4897 8562 4903 8569
rect 3271 8551 3323 8557
rect 6535 8609 6587 8615
rect 4955 8597 4961 8605
rect 6529 8597 6535 8605
rect 4955 8569 6535 8597
rect 4955 8562 4961 8569
rect 6529 8562 6535 8569
rect 4903 8551 4955 8557
rect 8167 8609 8219 8615
rect 6587 8597 6593 8605
rect 8161 8597 8167 8605
rect 6587 8569 8167 8597
rect 6587 8562 6593 8569
rect 8161 8562 8167 8569
rect 6535 8551 6587 8557
rect 9799 8609 9851 8615
rect 8219 8597 8225 8605
rect 9793 8597 9799 8605
rect 8219 8569 9799 8597
rect 8219 8562 8225 8569
rect 9793 8562 9799 8569
rect 8167 8551 8219 8557
rect 9851 8562 9857 8605
rect 9799 8551 9851 8557
rect 7 8405 59 8411
rect 1 8358 7 8401
rect 1639 8405 1691 8411
rect 59 8393 65 8401
rect 1633 8393 1639 8401
rect 59 8365 1639 8393
rect 59 8358 65 8365
rect 1633 8358 1639 8365
rect 7 8347 59 8353
rect 3271 8405 3323 8411
rect 1691 8393 1697 8401
rect 3265 8393 3271 8401
rect 1691 8365 3271 8393
rect 1691 8358 1697 8365
rect 3265 8358 3271 8365
rect 1639 8347 1691 8353
rect 4903 8405 4955 8411
rect 3323 8393 3329 8401
rect 4897 8393 4903 8401
rect 3323 8365 4903 8393
rect 3323 8358 3329 8365
rect 4897 8358 4903 8365
rect 3271 8347 3323 8353
rect 6535 8405 6587 8411
rect 4955 8393 4961 8401
rect 6529 8393 6535 8401
rect 4955 8365 6535 8393
rect 4955 8358 4961 8365
rect 6529 8358 6535 8365
rect 4903 8347 4955 8353
rect 8167 8405 8219 8411
rect 6587 8393 6593 8401
rect 8161 8393 8167 8401
rect 6587 8365 8167 8393
rect 6587 8358 6593 8365
rect 8161 8358 8167 8365
rect 6535 8347 6587 8353
rect 9799 8405 9851 8411
rect 8219 8393 8225 8401
rect 9793 8393 9799 8401
rect 8219 8365 9799 8393
rect 8219 8358 8225 8365
rect 9793 8358 9799 8365
rect 8167 8347 8219 8353
rect 9851 8358 9857 8401
rect 9799 8347 9851 8353
rect 7 8201 59 8207
rect 1 8154 7 8197
rect 1639 8201 1691 8207
rect 59 8189 65 8197
rect 1633 8189 1639 8197
rect 59 8161 1639 8189
rect 59 8154 65 8161
rect 1633 8154 1639 8161
rect 7 8143 59 8149
rect 3271 8201 3323 8207
rect 1691 8189 1697 8197
rect 3265 8189 3271 8197
rect 1691 8161 3271 8189
rect 1691 8154 1697 8161
rect 3265 8154 3271 8161
rect 1639 8143 1691 8149
rect 4903 8201 4955 8207
rect 3323 8189 3329 8197
rect 4897 8189 4903 8197
rect 3323 8161 4903 8189
rect 3323 8154 3329 8161
rect 4897 8154 4903 8161
rect 3271 8143 3323 8149
rect 6535 8201 6587 8207
rect 4955 8189 4961 8197
rect 6529 8189 6535 8197
rect 4955 8161 6535 8189
rect 4955 8154 4961 8161
rect 6529 8154 6535 8161
rect 4903 8143 4955 8149
rect 8167 8201 8219 8207
rect 6587 8189 6593 8197
rect 8161 8189 8167 8197
rect 6587 8161 8167 8189
rect 6587 8154 6593 8161
rect 8161 8154 8167 8161
rect 6535 8143 6587 8149
rect 9799 8201 9851 8207
rect 8219 8189 8225 8197
rect 9793 8189 9799 8197
rect 8219 8161 9799 8189
rect 8219 8154 8225 8161
rect 9793 8154 9799 8161
rect 8167 8143 8219 8149
rect 9851 8154 9857 8197
rect 9799 8143 9851 8149
rect 7 7997 59 8003
rect 1 7950 7 7993
rect 1639 7997 1691 8003
rect 59 7985 65 7993
rect 1633 7985 1639 7993
rect 59 7957 1639 7985
rect 59 7950 65 7957
rect 1633 7950 1639 7957
rect 7 7939 59 7945
rect 3271 7997 3323 8003
rect 1691 7985 1697 7993
rect 3265 7985 3271 7993
rect 1691 7957 3271 7985
rect 1691 7950 1697 7957
rect 3265 7950 3271 7957
rect 1639 7939 1691 7945
rect 4903 7997 4955 8003
rect 3323 7985 3329 7993
rect 4897 7985 4903 7993
rect 3323 7957 4903 7985
rect 3323 7950 3329 7957
rect 4897 7950 4903 7957
rect 3271 7939 3323 7945
rect 6535 7997 6587 8003
rect 4955 7985 4961 7993
rect 6529 7985 6535 7993
rect 4955 7957 6535 7985
rect 4955 7950 4961 7957
rect 6529 7950 6535 7957
rect 4903 7939 4955 7945
rect 8167 7997 8219 8003
rect 6587 7985 6593 7993
rect 8161 7985 8167 7993
rect 6587 7957 8167 7985
rect 6587 7950 6593 7957
rect 8161 7950 8167 7957
rect 6535 7939 6587 7945
rect 9799 7997 9851 8003
rect 8219 7985 8225 7993
rect 9793 7985 9799 7993
rect 8219 7957 9799 7985
rect 8219 7950 8225 7957
rect 9793 7950 9799 7957
rect 8167 7939 8219 7945
rect 9851 7950 9857 7993
rect 9799 7939 9851 7945
rect 212 7791 218 7843
rect 270 7831 276 7843
rect 416 7831 422 7843
rect 270 7803 422 7831
rect 270 7791 276 7803
rect 416 7791 422 7803
rect 474 7831 480 7843
rect 620 7831 626 7843
rect 474 7803 626 7831
rect 474 7791 480 7803
rect 620 7791 626 7803
rect 678 7831 684 7843
rect 824 7831 830 7843
rect 678 7803 830 7831
rect 678 7791 684 7803
rect 824 7791 830 7803
rect 882 7831 888 7843
rect 1028 7831 1034 7843
rect 882 7803 1034 7831
rect 882 7791 888 7803
rect 1028 7791 1034 7803
rect 1086 7831 1092 7843
rect 1232 7831 1238 7843
rect 1086 7803 1238 7831
rect 1086 7791 1092 7803
rect 1232 7791 1238 7803
rect 1290 7831 1296 7843
rect 1436 7831 1442 7843
rect 1290 7803 1442 7831
rect 1290 7791 1296 7803
rect 1436 7791 1442 7803
rect 1494 7831 1500 7843
rect 1640 7831 1646 7843
rect 1494 7803 1646 7831
rect 1494 7791 1500 7803
rect 1640 7791 1646 7803
rect 1698 7831 1704 7843
rect 1844 7831 1850 7843
rect 1698 7803 1850 7831
rect 1698 7791 1704 7803
rect 1844 7791 1850 7803
rect 1902 7831 1908 7843
rect 2048 7831 2054 7843
rect 1902 7803 2054 7831
rect 1902 7791 1908 7803
rect 2048 7791 2054 7803
rect 2106 7831 2112 7843
rect 2252 7831 2258 7843
rect 2106 7803 2258 7831
rect 2106 7791 2112 7803
rect 2252 7791 2258 7803
rect 2310 7831 2316 7843
rect 2456 7831 2462 7843
rect 2310 7803 2462 7831
rect 2310 7791 2316 7803
rect 2456 7791 2462 7803
rect 2514 7831 2520 7843
rect 2660 7831 2666 7843
rect 2514 7803 2666 7831
rect 2514 7791 2520 7803
rect 2660 7791 2666 7803
rect 2718 7831 2724 7843
rect 2864 7831 2870 7843
rect 2718 7803 2870 7831
rect 2718 7791 2724 7803
rect 2864 7791 2870 7803
rect 2922 7831 2928 7843
rect 3068 7831 3074 7843
rect 2922 7803 3074 7831
rect 2922 7791 2928 7803
rect 3068 7791 3074 7803
rect 3126 7831 3132 7843
rect 3272 7831 3278 7843
rect 3126 7803 3278 7831
rect 3126 7791 3132 7803
rect 3272 7791 3278 7803
rect 3330 7831 3336 7843
rect 3476 7831 3482 7843
rect 3330 7803 3482 7831
rect 3330 7791 3336 7803
rect 3476 7791 3482 7803
rect 3534 7831 3540 7843
rect 3680 7831 3686 7843
rect 3534 7803 3686 7831
rect 3534 7791 3540 7803
rect 3680 7791 3686 7803
rect 3738 7831 3744 7843
rect 3884 7831 3890 7843
rect 3738 7803 3890 7831
rect 3738 7791 3744 7803
rect 3884 7791 3890 7803
rect 3942 7831 3948 7843
rect 4088 7831 4094 7843
rect 3942 7803 4094 7831
rect 3942 7791 3948 7803
rect 4088 7791 4094 7803
rect 4146 7831 4152 7843
rect 4292 7831 4298 7843
rect 4146 7803 4298 7831
rect 4146 7791 4152 7803
rect 4292 7791 4298 7803
rect 4350 7831 4356 7843
rect 4496 7831 4502 7843
rect 4350 7803 4502 7831
rect 4350 7791 4356 7803
rect 4496 7791 4502 7803
rect 4554 7831 4560 7843
rect 4700 7831 4706 7843
rect 4554 7803 4706 7831
rect 4554 7791 4560 7803
rect 4700 7791 4706 7803
rect 4758 7831 4764 7843
rect 4904 7831 4910 7843
rect 4758 7803 4910 7831
rect 4758 7791 4764 7803
rect 4904 7791 4910 7803
rect 4962 7831 4968 7843
rect 5108 7831 5114 7843
rect 4962 7803 5114 7831
rect 4962 7791 4968 7803
rect 5108 7791 5114 7803
rect 5166 7831 5172 7843
rect 5312 7831 5318 7843
rect 5166 7803 5318 7831
rect 5166 7791 5172 7803
rect 5312 7791 5318 7803
rect 5370 7831 5376 7843
rect 5516 7831 5522 7843
rect 5370 7803 5522 7831
rect 5370 7791 5376 7803
rect 5516 7791 5522 7803
rect 5574 7831 5580 7843
rect 5720 7831 5726 7843
rect 5574 7803 5726 7831
rect 5574 7791 5580 7803
rect 5720 7791 5726 7803
rect 5778 7831 5784 7843
rect 5924 7831 5930 7843
rect 5778 7803 5930 7831
rect 5778 7791 5784 7803
rect 5924 7791 5930 7803
rect 5982 7831 5988 7843
rect 6128 7831 6134 7843
rect 5982 7803 6134 7831
rect 5982 7791 5988 7803
rect 6128 7791 6134 7803
rect 6186 7831 6192 7843
rect 6332 7831 6338 7843
rect 6186 7803 6338 7831
rect 6186 7791 6192 7803
rect 6332 7791 6338 7803
rect 6390 7831 6396 7843
rect 6536 7831 6542 7843
rect 6390 7803 6542 7831
rect 6390 7791 6396 7803
rect 6536 7791 6542 7803
rect 6594 7831 6600 7843
rect 6740 7831 6746 7843
rect 6594 7803 6746 7831
rect 6594 7791 6600 7803
rect 6740 7791 6746 7803
rect 6798 7831 6804 7843
rect 6944 7831 6950 7843
rect 6798 7803 6950 7831
rect 6798 7791 6804 7803
rect 6944 7791 6950 7803
rect 7002 7831 7008 7843
rect 7148 7831 7154 7843
rect 7002 7803 7154 7831
rect 7002 7791 7008 7803
rect 7148 7791 7154 7803
rect 7206 7831 7212 7843
rect 7352 7831 7358 7843
rect 7206 7803 7358 7831
rect 7206 7791 7212 7803
rect 7352 7791 7358 7803
rect 7410 7831 7416 7843
rect 7556 7831 7562 7843
rect 7410 7803 7562 7831
rect 7410 7791 7416 7803
rect 7556 7791 7562 7803
rect 7614 7831 7620 7843
rect 7760 7831 7766 7843
rect 7614 7803 7766 7831
rect 7614 7791 7620 7803
rect 7760 7791 7766 7803
rect 7818 7831 7824 7843
rect 7964 7831 7970 7843
rect 7818 7803 7970 7831
rect 7818 7791 7824 7803
rect 7964 7791 7970 7803
rect 8022 7831 8028 7843
rect 8168 7831 8174 7843
rect 8022 7803 8174 7831
rect 8022 7791 8028 7803
rect 8168 7791 8174 7803
rect 8226 7831 8232 7843
rect 8372 7831 8378 7843
rect 8226 7803 8378 7831
rect 8226 7791 8232 7803
rect 8372 7791 8378 7803
rect 8430 7831 8436 7843
rect 8576 7831 8582 7843
rect 8430 7803 8582 7831
rect 8430 7791 8436 7803
rect 8576 7791 8582 7803
rect 8634 7831 8640 7843
rect 8780 7831 8786 7843
rect 8634 7803 8786 7831
rect 8634 7791 8640 7803
rect 8780 7791 8786 7803
rect 8838 7831 8844 7843
rect 8984 7831 8990 7843
rect 8838 7803 8990 7831
rect 8838 7791 8844 7803
rect 8984 7791 8990 7803
rect 9042 7831 9048 7843
rect 9188 7831 9194 7843
rect 9042 7803 9194 7831
rect 9042 7791 9048 7803
rect 9188 7791 9194 7803
rect 9246 7831 9252 7843
rect 9392 7831 9398 7843
rect 9246 7803 9398 7831
rect 9246 7791 9252 7803
rect 9392 7791 9398 7803
rect 9450 7831 9456 7843
rect 9596 7831 9602 7843
rect 9450 7803 9602 7831
rect 9450 7791 9456 7803
rect 9596 7791 9602 7803
rect 9654 7831 9660 7843
rect 9814 7831 9820 7843
rect 9654 7803 9820 7831
rect 9654 7791 9660 7803
rect 9814 7791 9820 7803
rect 9872 7791 9878 7843
rect 7 7689 59 7695
rect 1 7642 7 7685
rect 1639 7689 1691 7695
rect 59 7677 65 7685
rect 1633 7677 1639 7685
rect 59 7649 1639 7677
rect 59 7642 65 7649
rect 1633 7642 1639 7649
rect 7 7631 59 7637
rect 3271 7689 3323 7695
rect 1691 7677 1697 7685
rect 3265 7677 3271 7685
rect 1691 7649 3271 7677
rect 1691 7642 1697 7649
rect 3265 7642 3271 7649
rect 1639 7631 1691 7637
rect 4903 7689 4955 7695
rect 3323 7677 3329 7685
rect 4897 7677 4903 7685
rect 3323 7649 4903 7677
rect 3323 7642 3329 7649
rect 4897 7642 4903 7649
rect 3271 7631 3323 7637
rect 6535 7689 6587 7695
rect 4955 7677 4961 7685
rect 6529 7677 6535 7685
rect 4955 7649 6535 7677
rect 4955 7642 4961 7649
rect 6529 7642 6535 7649
rect 4903 7631 4955 7637
rect 8167 7689 8219 7695
rect 6587 7677 6593 7685
rect 8161 7677 8167 7685
rect 6587 7649 8167 7677
rect 6587 7642 6593 7649
rect 8161 7642 8167 7649
rect 6535 7631 6587 7637
rect 9799 7689 9851 7695
rect 8219 7677 8225 7685
rect 9793 7677 9799 7685
rect 8219 7649 9799 7677
rect 8219 7642 8225 7649
rect 9793 7642 9799 7649
rect 8167 7631 8219 7637
rect 9851 7642 9857 7685
rect 9799 7631 9851 7637
rect 7 7485 59 7491
rect 1 7438 7 7481
rect 1639 7485 1691 7491
rect 59 7473 65 7481
rect 1633 7473 1639 7481
rect 59 7445 1639 7473
rect 59 7438 65 7445
rect 1633 7438 1639 7445
rect 7 7427 59 7433
rect 3271 7485 3323 7491
rect 1691 7473 1697 7481
rect 3265 7473 3271 7481
rect 1691 7445 3271 7473
rect 1691 7438 1697 7445
rect 3265 7438 3271 7445
rect 1639 7427 1691 7433
rect 4903 7485 4955 7491
rect 3323 7473 3329 7481
rect 4897 7473 4903 7481
rect 3323 7445 4903 7473
rect 3323 7438 3329 7445
rect 4897 7438 4903 7445
rect 3271 7427 3323 7433
rect 6535 7485 6587 7491
rect 4955 7473 4961 7481
rect 6529 7473 6535 7481
rect 4955 7445 6535 7473
rect 4955 7438 4961 7445
rect 6529 7438 6535 7445
rect 4903 7427 4955 7433
rect 8167 7485 8219 7491
rect 6587 7473 6593 7481
rect 8161 7473 8167 7481
rect 6587 7445 8167 7473
rect 6587 7438 6593 7445
rect 8161 7438 8167 7445
rect 6535 7427 6587 7433
rect 9799 7485 9851 7491
rect 8219 7473 8225 7481
rect 9793 7473 9799 7481
rect 8219 7445 9799 7473
rect 8219 7438 8225 7445
rect 9793 7438 9799 7445
rect 8167 7427 8219 7433
rect 9851 7438 9857 7481
rect 9799 7427 9851 7433
rect 7 7281 59 7287
rect 1 7234 7 7277
rect 1639 7281 1691 7287
rect 59 7269 65 7277
rect 1633 7269 1639 7277
rect 59 7241 1639 7269
rect 59 7234 65 7241
rect 1633 7234 1639 7241
rect 7 7223 59 7229
rect 3271 7281 3323 7287
rect 1691 7269 1697 7277
rect 3265 7269 3271 7277
rect 1691 7241 3271 7269
rect 1691 7234 1697 7241
rect 3265 7234 3271 7241
rect 1639 7223 1691 7229
rect 4903 7281 4955 7287
rect 3323 7269 3329 7277
rect 4897 7269 4903 7277
rect 3323 7241 4903 7269
rect 3323 7234 3329 7241
rect 4897 7234 4903 7241
rect 3271 7223 3323 7229
rect 6535 7281 6587 7287
rect 4955 7269 4961 7277
rect 6529 7269 6535 7277
rect 4955 7241 6535 7269
rect 4955 7234 4961 7241
rect 6529 7234 6535 7241
rect 4903 7223 4955 7229
rect 8167 7281 8219 7287
rect 6587 7269 6593 7277
rect 8161 7269 8167 7277
rect 6587 7241 8167 7269
rect 6587 7234 6593 7241
rect 8161 7234 8167 7241
rect 6535 7223 6587 7229
rect 9799 7281 9851 7287
rect 8219 7269 8225 7277
rect 9793 7269 9799 7277
rect 8219 7241 9799 7269
rect 8219 7234 8225 7241
rect 9793 7234 9799 7241
rect 8167 7223 8219 7229
rect 9851 7234 9857 7277
rect 9799 7223 9851 7229
rect 7 7077 59 7083
rect 1 7030 7 7073
rect 1639 7077 1691 7083
rect 59 7065 65 7073
rect 1633 7065 1639 7073
rect 59 7037 1639 7065
rect 59 7030 65 7037
rect 1633 7030 1639 7037
rect 7 7019 59 7025
rect 3271 7077 3323 7083
rect 1691 7065 1697 7073
rect 3265 7065 3271 7073
rect 1691 7037 3271 7065
rect 1691 7030 1697 7037
rect 3265 7030 3271 7037
rect 1639 7019 1691 7025
rect 4903 7077 4955 7083
rect 3323 7065 3329 7073
rect 4897 7065 4903 7073
rect 3323 7037 4903 7065
rect 3323 7030 3329 7037
rect 4897 7030 4903 7037
rect 3271 7019 3323 7025
rect 6535 7077 6587 7083
rect 4955 7065 4961 7073
rect 6529 7065 6535 7073
rect 4955 7037 6535 7065
rect 4955 7030 4961 7037
rect 6529 7030 6535 7037
rect 4903 7019 4955 7025
rect 8167 7077 8219 7083
rect 6587 7065 6593 7073
rect 8161 7065 8167 7073
rect 6587 7037 8167 7065
rect 6587 7030 6593 7037
rect 8161 7030 8167 7037
rect 6535 7019 6587 7025
rect 9799 7077 9851 7083
rect 8219 7065 8225 7073
rect 9793 7065 9799 7073
rect 8219 7037 9799 7065
rect 8219 7030 8225 7037
rect 9793 7030 9799 7037
rect 8167 7019 8219 7025
rect 9851 7030 9857 7073
rect 9799 7019 9851 7025
rect 7 6873 59 6879
rect 1 6826 7 6869
rect 1639 6873 1691 6879
rect 59 6861 65 6869
rect 1633 6861 1639 6869
rect 59 6833 1639 6861
rect 59 6826 65 6833
rect 1633 6826 1639 6833
rect 7 6815 59 6821
rect 3271 6873 3323 6879
rect 1691 6861 1697 6869
rect 3265 6861 3271 6869
rect 1691 6833 3271 6861
rect 1691 6826 1697 6833
rect 3265 6826 3271 6833
rect 1639 6815 1691 6821
rect 4903 6873 4955 6879
rect 3323 6861 3329 6869
rect 4897 6861 4903 6869
rect 3323 6833 4903 6861
rect 3323 6826 3329 6833
rect 4897 6826 4903 6833
rect 3271 6815 3323 6821
rect 6535 6873 6587 6879
rect 4955 6861 4961 6869
rect 6529 6861 6535 6869
rect 4955 6833 6535 6861
rect 4955 6826 4961 6833
rect 6529 6826 6535 6833
rect 4903 6815 4955 6821
rect 8167 6873 8219 6879
rect 6587 6861 6593 6869
rect 8161 6861 8167 6869
rect 6587 6833 8167 6861
rect 6587 6826 6593 6833
rect 8161 6826 8167 6833
rect 6535 6815 6587 6821
rect 9799 6873 9851 6879
rect 8219 6861 8225 6869
rect 9793 6861 9799 6869
rect 8219 6833 9799 6861
rect 8219 6826 8225 6833
rect 9793 6826 9799 6833
rect 8167 6815 8219 6821
rect 9851 6826 9857 6869
rect 9799 6815 9851 6821
rect 7 6669 59 6675
rect 1 6622 7 6665
rect 1639 6669 1691 6675
rect 59 6657 65 6665
rect 1633 6657 1639 6665
rect 59 6629 1639 6657
rect 59 6622 65 6629
rect 1633 6622 1639 6629
rect 7 6611 59 6617
rect 3271 6669 3323 6675
rect 1691 6657 1697 6665
rect 3265 6657 3271 6665
rect 1691 6629 3271 6657
rect 1691 6622 1697 6629
rect 3265 6622 3271 6629
rect 1639 6611 1691 6617
rect 4903 6669 4955 6675
rect 3323 6657 3329 6665
rect 4897 6657 4903 6665
rect 3323 6629 4903 6657
rect 3323 6622 3329 6629
rect 4897 6622 4903 6629
rect 3271 6611 3323 6617
rect 6535 6669 6587 6675
rect 4955 6657 4961 6665
rect 6529 6657 6535 6665
rect 4955 6629 6535 6657
rect 4955 6622 4961 6629
rect 6529 6622 6535 6629
rect 4903 6611 4955 6617
rect 8167 6669 8219 6675
rect 6587 6657 6593 6665
rect 8161 6657 8167 6665
rect 6587 6629 8167 6657
rect 6587 6622 6593 6629
rect 8161 6622 8167 6629
rect 6535 6611 6587 6617
rect 9799 6669 9851 6675
rect 8219 6657 8225 6665
rect 9793 6657 9799 6665
rect 8219 6629 9799 6657
rect 8219 6622 8225 6629
rect 9793 6622 9799 6629
rect 8167 6611 8219 6617
rect 9851 6622 9857 6665
rect 9799 6611 9851 6617
rect 7 6465 59 6471
rect 1 6418 7 6461
rect 1639 6465 1691 6471
rect 59 6453 65 6461
rect 1633 6453 1639 6461
rect 59 6425 1639 6453
rect 59 6418 65 6425
rect 1633 6418 1639 6425
rect 7 6407 59 6413
rect 3271 6465 3323 6471
rect 1691 6453 1697 6461
rect 3265 6453 3271 6461
rect 1691 6425 3271 6453
rect 1691 6418 1697 6425
rect 3265 6418 3271 6425
rect 1639 6407 1691 6413
rect 4903 6465 4955 6471
rect 3323 6453 3329 6461
rect 4897 6453 4903 6461
rect 3323 6425 4903 6453
rect 3323 6418 3329 6425
rect 4897 6418 4903 6425
rect 3271 6407 3323 6413
rect 6535 6465 6587 6471
rect 4955 6453 4961 6461
rect 6529 6453 6535 6461
rect 4955 6425 6535 6453
rect 4955 6418 4961 6425
rect 6529 6418 6535 6425
rect 4903 6407 4955 6413
rect 8167 6465 8219 6471
rect 6587 6453 6593 6461
rect 8161 6453 8167 6461
rect 6587 6425 8167 6453
rect 6587 6418 6593 6425
rect 8161 6418 8167 6425
rect 6535 6407 6587 6413
rect 9799 6465 9851 6471
rect 8219 6453 8225 6461
rect 9793 6453 9799 6461
rect 8219 6425 9799 6453
rect 8219 6418 8225 6425
rect 9793 6418 9799 6425
rect 8167 6407 8219 6413
rect 9851 6418 9857 6461
rect 9799 6407 9851 6413
rect 7 6261 59 6267
rect 1 6214 7 6257
rect 1639 6261 1691 6267
rect 59 6249 65 6257
rect 1633 6249 1639 6257
rect 59 6221 1639 6249
rect 59 6214 65 6221
rect 1633 6214 1639 6221
rect 7 6203 59 6209
rect 3271 6261 3323 6267
rect 1691 6249 1697 6257
rect 3265 6249 3271 6257
rect 1691 6221 3271 6249
rect 1691 6214 1697 6221
rect 3265 6214 3271 6221
rect 1639 6203 1691 6209
rect 4903 6261 4955 6267
rect 3323 6249 3329 6257
rect 4897 6249 4903 6257
rect 3323 6221 4903 6249
rect 3323 6214 3329 6221
rect 4897 6214 4903 6221
rect 3271 6203 3323 6209
rect 6535 6261 6587 6267
rect 4955 6249 4961 6257
rect 6529 6249 6535 6257
rect 4955 6221 6535 6249
rect 4955 6214 4961 6221
rect 6529 6214 6535 6221
rect 4903 6203 4955 6209
rect 8167 6261 8219 6267
rect 6587 6249 6593 6257
rect 8161 6249 8167 6257
rect 6587 6221 8167 6249
rect 6587 6214 6593 6221
rect 8161 6214 8167 6221
rect 6535 6203 6587 6209
rect 9799 6261 9851 6267
rect 8219 6249 8225 6257
rect 9793 6249 9799 6257
rect 8219 6221 9799 6249
rect 8219 6214 8225 6221
rect 9793 6214 9799 6221
rect 8167 6203 8219 6209
rect 9851 6214 9857 6257
rect 9799 6203 9851 6209
rect 212 6055 218 6107
rect 270 6095 276 6107
rect 416 6095 422 6107
rect 270 6067 422 6095
rect 270 6055 276 6067
rect 416 6055 422 6067
rect 474 6095 480 6107
rect 620 6095 626 6107
rect 474 6067 626 6095
rect 474 6055 480 6067
rect 620 6055 626 6067
rect 678 6095 684 6107
rect 824 6095 830 6107
rect 678 6067 830 6095
rect 678 6055 684 6067
rect 824 6055 830 6067
rect 882 6095 888 6107
rect 1028 6095 1034 6107
rect 882 6067 1034 6095
rect 882 6055 888 6067
rect 1028 6055 1034 6067
rect 1086 6095 1092 6107
rect 1232 6095 1238 6107
rect 1086 6067 1238 6095
rect 1086 6055 1092 6067
rect 1232 6055 1238 6067
rect 1290 6095 1296 6107
rect 1436 6095 1442 6107
rect 1290 6067 1442 6095
rect 1290 6055 1296 6067
rect 1436 6055 1442 6067
rect 1494 6095 1500 6107
rect 1640 6095 1646 6107
rect 1494 6067 1646 6095
rect 1494 6055 1500 6067
rect 1640 6055 1646 6067
rect 1698 6095 1704 6107
rect 1844 6095 1850 6107
rect 1698 6067 1850 6095
rect 1698 6055 1704 6067
rect 1844 6055 1850 6067
rect 1902 6095 1908 6107
rect 2048 6095 2054 6107
rect 1902 6067 2054 6095
rect 1902 6055 1908 6067
rect 2048 6055 2054 6067
rect 2106 6095 2112 6107
rect 2252 6095 2258 6107
rect 2106 6067 2258 6095
rect 2106 6055 2112 6067
rect 2252 6055 2258 6067
rect 2310 6095 2316 6107
rect 2456 6095 2462 6107
rect 2310 6067 2462 6095
rect 2310 6055 2316 6067
rect 2456 6055 2462 6067
rect 2514 6095 2520 6107
rect 2660 6095 2666 6107
rect 2514 6067 2666 6095
rect 2514 6055 2520 6067
rect 2660 6055 2666 6067
rect 2718 6095 2724 6107
rect 2864 6095 2870 6107
rect 2718 6067 2870 6095
rect 2718 6055 2724 6067
rect 2864 6055 2870 6067
rect 2922 6095 2928 6107
rect 3068 6095 3074 6107
rect 2922 6067 3074 6095
rect 2922 6055 2928 6067
rect 3068 6055 3074 6067
rect 3126 6095 3132 6107
rect 3272 6095 3278 6107
rect 3126 6067 3278 6095
rect 3126 6055 3132 6067
rect 3272 6055 3278 6067
rect 3330 6095 3336 6107
rect 3476 6095 3482 6107
rect 3330 6067 3482 6095
rect 3330 6055 3336 6067
rect 3476 6055 3482 6067
rect 3534 6095 3540 6107
rect 3680 6095 3686 6107
rect 3534 6067 3686 6095
rect 3534 6055 3540 6067
rect 3680 6055 3686 6067
rect 3738 6095 3744 6107
rect 3884 6095 3890 6107
rect 3738 6067 3890 6095
rect 3738 6055 3744 6067
rect 3884 6055 3890 6067
rect 3942 6095 3948 6107
rect 4088 6095 4094 6107
rect 3942 6067 4094 6095
rect 3942 6055 3948 6067
rect 4088 6055 4094 6067
rect 4146 6095 4152 6107
rect 4292 6095 4298 6107
rect 4146 6067 4298 6095
rect 4146 6055 4152 6067
rect 4292 6055 4298 6067
rect 4350 6095 4356 6107
rect 4496 6095 4502 6107
rect 4350 6067 4502 6095
rect 4350 6055 4356 6067
rect 4496 6055 4502 6067
rect 4554 6095 4560 6107
rect 4700 6095 4706 6107
rect 4554 6067 4706 6095
rect 4554 6055 4560 6067
rect 4700 6055 4706 6067
rect 4758 6095 4764 6107
rect 4904 6095 4910 6107
rect 4758 6067 4910 6095
rect 4758 6055 4764 6067
rect 4904 6055 4910 6067
rect 4962 6095 4968 6107
rect 5108 6095 5114 6107
rect 4962 6067 5114 6095
rect 4962 6055 4968 6067
rect 5108 6055 5114 6067
rect 5166 6095 5172 6107
rect 5312 6095 5318 6107
rect 5166 6067 5318 6095
rect 5166 6055 5172 6067
rect 5312 6055 5318 6067
rect 5370 6095 5376 6107
rect 5516 6095 5522 6107
rect 5370 6067 5522 6095
rect 5370 6055 5376 6067
rect 5516 6055 5522 6067
rect 5574 6095 5580 6107
rect 5720 6095 5726 6107
rect 5574 6067 5726 6095
rect 5574 6055 5580 6067
rect 5720 6055 5726 6067
rect 5778 6095 5784 6107
rect 5924 6095 5930 6107
rect 5778 6067 5930 6095
rect 5778 6055 5784 6067
rect 5924 6055 5930 6067
rect 5982 6095 5988 6107
rect 6128 6095 6134 6107
rect 5982 6067 6134 6095
rect 5982 6055 5988 6067
rect 6128 6055 6134 6067
rect 6186 6095 6192 6107
rect 6332 6095 6338 6107
rect 6186 6067 6338 6095
rect 6186 6055 6192 6067
rect 6332 6055 6338 6067
rect 6390 6095 6396 6107
rect 6536 6095 6542 6107
rect 6390 6067 6542 6095
rect 6390 6055 6396 6067
rect 6536 6055 6542 6067
rect 6594 6095 6600 6107
rect 6740 6095 6746 6107
rect 6594 6067 6746 6095
rect 6594 6055 6600 6067
rect 6740 6055 6746 6067
rect 6798 6095 6804 6107
rect 6944 6095 6950 6107
rect 6798 6067 6950 6095
rect 6798 6055 6804 6067
rect 6944 6055 6950 6067
rect 7002 6095 7008 6107
rect 7148 6095 7154 6107
rect 7002 6067 7154 6095
rect 7002 6055 7008 6067
rect 7148 6055 7154 6067
rect 7206 6095 7212 6107
rect 7352 6095 7358 6107
rect 7206 6067 7358 6095
rect 7206 6055 7212 6067
rect 7352 6055 7358 6067
rect 7410 6095 7416 6107
rect 7556 6095 7562 6107
rect 7410 6067 7562 6095
rect 7410 6055 7416 6067
rect 7556 6055 7562 6067
rect 7614 6095 7620 6107
rect 7760 6095 7766 6107
rect 7614 6067 7766 6095
rect 7614 6055 7620 6067
rect 7760 6055 7766 6067
rect 7818 6095 7824 6107
rect 7964 6095 7970 6107
rect 7818 6067 7970 6095
rect 7818 6055 7824 6067
rect 7964 6055 7970 6067
rect 8022 6095 8028 6107
rect 8168 6095 8174 6107
rect 8022 6067 8174 6095
rect 8022 6055 8028 6067
rect 8168 6055 8174 6067
rect 8226 6095 8232 6107
rect 8372 6095 8378 6107
rect 8226 6067 8378 6095
rect 8226 6055 8232 6067
rect 8372 6055 8378 6067
rect 8430 6095 8436 6107
rect 8576 6095 8582 6107
rect 8430 6067 8582 6095
rect 8430 6055 8436 6067
rect 8576 6055 8582 6067
rect 8634 6095 8640 6107
rect 8780 6095 8786 6107
rect 8634 6067 8786 6095
rect 8634 6055 8640 6067
rect 8780 6055 8786 6067
rect 8838 6095 8844 6107
rect 8984 6095 8990 6107
rect 8838 6067 8990 6095
rect 8838 6055 8844 6067
rect 8984 6055 8990 6067
rect 9042 6095 9048 6107
rect 9188 6095 9194 6107
rect 9042 6067 9194 6095
rect 9042 6055 9048 6067
rect 9188 6055 9194 6067
rect 9246 6095 9252 6107
rect 9392 6095 9398 6107
rect 9246 6067 9398 6095
rect 9246 6055 9252 6067
rect 9392 6055 9398 6067
rect 9450 6095 9456 6107
rect 9596 6095 9602 6107
rect 9450 6067 9602 6095
rect 9450 6055 9456 6067
rect 9596 6055 9602 6067
rect 9654 6095 9660 6107
rect 9814 6095 9820 6107
rect 9654 6067 9820 6095
rect 9654 6055 9660 6067
rect 9814 6055 9820 6067
rect 9872 6055 9878 6107
rect 7 5953 59 5959
rect 1 5906 7 5949
rect 1639 5953 1691 5959
rect 59 5941 65 5949
rect 1633 5941 1639 5949
rect 59 5913 1639 5941
rect 59 5906 65 5913
rect 1633 5906 1639 5913
rect 7 5895 59 5901
rect 3271 5953 3323 5959
rect 1691 5941 1697 5949
rect 3265 5941 3271 5949
rect 1691 5913 3271 5941
rect 1691 5906 1697 5913
rect 3265 5906 3271 5913
rect 1639 5895 1691 5901
rect 4903 5953 4955 5959
rect 3323 5941 3329 5949
rect 4897 5941 4903 5949
rect 3323 5913 4903 5941
rect 3323 5906 3329 5913
rect 4897 5906 4903 5913
rect 3271 5895 3323 5901
rect 6535 5953 6587 5959
rect 4955 5941 4961 5949
rect 6529 5941 6535 5949
rect 4955 5913 6535 5941
rect 4955 5906 4961 5913
rect 6529 5906 6535 5913
rect 4903 5895 4955 5901
rect 8167 5953 8219 5959
rect 6587 5941 6593 5949
rect 8161 5941 8167 5949
rect 6587 5913 8167 5941
rect 6587 5906 6593 5913
rect 8161 5906 8167 5913
rect 6535 5895 6587 5901
rect 9799 5953 9851 5959
rect 8219 5941 8225 5949
rect 9793 5941 9799 5949
rect 8219 5913 9799 5941
rect 8219 5906 8225 5913
rect 9793 5906 9799 5913
rect 8167 5895 8219 5901
rect 9851 5906 9857 5949
rect 9799 5895 9851 5901
rect 7 5749 59 5755
rect 1 5702 7 5745
rect 1639 5749 1691 5755
rect 59 5737 65 5745
rect 1633 5737 1639 5745
rect 59 5709 1639 5737
rect 59 5702 65 5709
rect 1633 5702 1639 5709
rect 7 5691 59 5697
rect 3271 5749 3323 5755
rect 1691 5737 1697 5745
rect 3265 5737 3271 5745
rect 1691 5709 3271 5737
rect 1691 5702 1697 5709
rect 3265 5702 3271 5709
rect 1639 5691 1691 5697
rect 4903 5749 4955 5755
rect 3323 5737 3329 5745
rect 4897 5737 4903 5745
rect 3323 5709 4903 5737
rect 3323 5702 3329 5709
rect 4897 5702 4903 5709
rect 3271 5691 3323 5697
rect 6535 5749 6587 5755
rect 4955 5737 4961 5745
rect 6529 5737 6535 5745
rect 4955 5709 6535 5737
rect 4955 5702 4961 5709
rect 6529 5702 6535 5709
rect 4903 5691 4955 5697
rect 8167 5749 8219 5755
rect 6587 5737 6593 5745
rect 8161 5737 8167 5745
rect 6587 5709 8167 5737
rect 6587 5702 6593 5709
rect 8161 5702 8167 5709
rect 6535 5691 6587 5697
rect 9799 5749 9851 5755
rect 8219 5737 8225 5745
rect 9793 5737 9799 5745
rect 8219 5709 9799 5737
rect 8219 5702 8225 5709
rect 9793 5702 9799 5709
rect 8167 5691 8219 5697
rect 9851 5702 9857 5745
rect 9799 5691 9851 5697
rect 7 5545 59 5551
rect 1 5498 7 5541
rect 1639 5545 1691 5551
rect 59 5533 65 5541
rect 1633 5533 1639 5541
rect 59 5505 1639 5533
rect 59 5498 65 5505
rect 1633 5498 1639 5505
rect 7 5487 59 5493
rect 3271 5545 3323 5551
rect 1691 5533 1697 5541
rect 3265 5533 3271 5541
rect 1691 5505 3271 5533
rect 1691 5498 1697 5505
rect 3265 5498 3271 5505
rect 1639 5487 1691 5493
rect 4903 5545 4955 5551
rect 3323 5533 3329 5541
rect 4897 5533 4903 5541
rect 3323 5505 4903 5533
rect 3323 5498 3329 5505
rect 4897 5498 4903 5505
rect 3271 5487 3323 5493
rect 6535 5545 6587 5551
rect 4955 5533 4961 5541
rect 6529 5533 6535 5541
rect 4955 5505 6535 5533
rect 4955 5498 4961 5505
rect 6529 5498 6535 5505
rect 4903 5487 4955 5493
rect 8167 5545 8219 5551
rect 6587 5533 6593 5541
rect 8161 5533 8167 5541
rect 6587 5505 8167 5533
rect 6587 5498 6593 5505
rect 8161 5498 8167 5505
rect 6535 5487 6587 5493
rect 9799 5545 9851 5551
rect 8219 5533 8225 5541
rect 9793 5533 9799 5541
rect 8219 5505 9799 5533
rect 8219 5498 8225 5505
rect 9793 5498 9799 5505
rect 8167 5487 8219 5493
rect 9851 5498 9857 5541
rect 9799 5487 9851 5493
rect 7 5341 59 5347
rect 1 5294 7 5337
rect 1639 5341 1691 5347
rect 59 5329 65 5337
rect 1633 5329 1639 5337
rect 59 5301 1639 5329
rect 59 5294 65 5301
rect 1633 5294 1639 5301
rect 7 5283 59 5289
rect 3271 5341 3323 5347
rect 1691 5329 1697 5337
rect 3265 5329 3271 5337
rect 1691 5301 3271 5329
rect 1691 5294 1697 5301
rect 3265 5294 3271 5301
rect 1639 5283 1691 5289
rect 4903 5341 4955 5347
rect 3323 5329 3329 5337
rect 4897 5329 4903 5337
rect 3323 5301 4903 5329
rect 3323 5294 3329 5301
rect 4897 5294 4903 5301
rect 3271 5283 3323 5289
rect 6535 5341 6587 5347
rect 4955 5329 4961 5337
rect 6529 5329 6535 5337
rect 4955 5301 6535 5329
rect 4955 5294 4961 5301
rect 6529 5294 6535 5301
rect 4903 5283 4955 5289
rect 8167 5341 8219 5347
rect 6587 5329 6593 5337
rect 8161 5329 8167 5337
rect 6587 5301 8167 5329
rect 6587 5294 6593 5301
rect 8161 5294 8167 5301
rect 6535 5283 6587 5289
rect 9799 5341 9851 5347
rect 8219 5329 8225 5337
rect 9793 5329 9799 5337
rect 8219 5301 9799 5329
rect 8219 5294 8225 5301
rect 9793 5294 9799 5301
rect 8167 5283 8219 5289
rect 9851 5294 9857 5337
rect 9799 5283 9851 5289
rect 7 5137 59 5143
rect 1 5090 7 5133
rect 1639 5137 1691 5143
rect 59 5125 65 5133
rect 1633 5125 1639 5133
rect 59 5097 1639 5125
rect 59 5090 65 5097
rect 1633 5090 1639 5097
rect 7 5079 59 5085
rect 3271 5137 3323 5143
rect 1691 5125 1697 5133
rect 3265 5125 3271 5133
rect 1691 5097 3271 5125
rect 1691 5090 1697 5097
rect 3265 5090 3271 5097
rect 1639 5079 1691 5085
rect 4903 5137 4955 5143
rect 3323 5125 3329 5133
rect 4897 5125 4903 5133
rect 3323 5097 4903 5125
rect 3323 5090 3329 5097
rect 4897 5090 4903 5097
rect 3271 5079 3323 5085
rect 6535 5137 6587 5143
rect 4955 5125 4961 5133
rect 6529 5125 6535 5133
rect 4955 5097 6535 5125
rect 4955 5090 4961 5097
rect 6529 5090 6535 5097
rect 4903 5079 4955 5085
rect 8167 5137 8219 5143
rect 6587 5125 6593 5133
rect 8161 5125 8167 5133
rect 6587 5097 8167 5125
rect 6587 5090 6593 5097
rect 8161 5090 8167 5097
rect 6535 5079 6587 5085
rect 9799 5137 9851 5143
rect 8219 5125 8225 5133
rect 9793 5125 9799 5133
rect 8219 5097 9799 5125
rect 8219 5090 8225 5097
rect 9793 5090 9799 5097
rect 8167 5079 8219 5085
rect 9851 5090 9857 5133
rect 9799 5079 9851 5085
rect 7 4933 59 4939
rect 1 4886 7 4929
rect 1639 4933 1691 4939
rect 59 4921 65 4929
rect 1633 4921 1639 4929
rect 59 4893 1639 4921
rect 59 4886 65 4893
rect 1633 4886 1639 4893
rect 7 4875 59 4881
rect 3271 4933 3323 4939
rect 1691 4921 1697 4929
rect 3265 4921 3271 4929
rect 1691 4893 3271 4921
rect 1691 4886 1697 4893
rect 3265 4886 3271 4893
rect 1639 4875 1691 4881
rect 4903 4933 4955 4939
rect 3323 4921 3329 4929
rect 4897 4921 4903 4929
rect 3323 4893 4903 4921
rect 3323 4886 3329 4893
rect 4897 4886 4903 4893
rect 3271 4875 3323 4881
rect 6535 4933 6587 4939
rect 4955 4921 4961 4929
rect 6529 4921 6535 4929
rect 4955 4893 6535 4921
rect 4955 4886 4961 4893
rect 6529 4886 6535 4893
rect 4903 4875 4955 4881
rect 8167 4933 8219 4939
rect 6587 4921 6593 4929
rect 8161 4921 8167 4929
rect 6587 4893 8167 4921
rect 6587 4886 6593 4893
rect 8161 4886 8167 4893
rect 6535 4875 6587 4881
rect 9799 4933 9851 4939
rect 8219 4921 8225 4929
rect 9793 4921 9799 4929
rect 8219 4893 9799 4921
rect 8219 4886 8225 4893
rect 9793 4886 9799 4893
rect 8167 4875 8219 4881
rect 9851 4886 9857 4929
rect 9799 4875 9851 4881
rect 7 4729 59 4735
rect 1 4682 7 4725
rect 1639 4729 1691 4735
rect 59 4717 65 4725
rect 1633 4717 1639 4725
rect 59 4689 1639 4717
rect 59 4682 65 4689
rect 1633 4682 1639 4689
rect 7 4671 59 4677
rect 3271 4729 3323 4735
rect 1691 4717 1697 4725
rect 3265 4717 3271 4725
rect 1691 4689 3271 4717
rect 1691 4682 1697 4689
rect 3265 4682 3271 4689
rect 1639 4671 1691 4677
rect 4903 4729 4955 4735
rect 3323 4717 3329 4725
rect 4897 4717 4903 4725
rect 3323 4689 4903 4717
rect 3323 4682 3329 4689
rect 4897 4682 4903 4689
rect 3271 4671 3323 4677
rect 6535 4729 6587 4735
rect 4955 4717 4961 4725
rect 6529 4717 6535 4725
rect 4955 4689 6535 4717
rect 4955 4682 4961 4689
rect 6529 4682 6535 4689
rect 4903 4671 4955 4677
rect 8167 4729 8219 4735
rect 6587 4717 6593 4725
rect 8161 4717 8167 4725
rect 6587 4689 8167 4717
rect 6587 4682 6593 4689
rect 8161 4682 8167 4689
rect 6535 4671 6587 4677
rect 9799 4729 9851 4735
rect 8219 4717 8225 4725
rect 9793 4717 9799 4725
rect 8219 4689 9799 4717
rect 8219 4682 8225 4689
rect 9793 4682 9799 4689
rect 8167 4671 8219 4677
rect 9851 4682 9857 4725
rect 9799 4671 9851 4677
rect 7 4525 59 4531
rect 1 4478 7 4521
rect 1639 4525 1691 4531
rect 59 4513 65 4521
rect 1633 4513 1639 4521
rect 59 4485 1639 4513
rect 59 4478 65 4485
rect 1633 4478 1639 4485
rect 7 4467 59 4473
rect 3271 4525 3323 4531
rect 1691 4513 1697 4521
rect 3265 4513 3271 4521
rect 1691 4485 3271 4513
rect 1691 4478 1697 4485
rect 3265 4478 3271 4485
rect 1639 4467 1691 4473
rect 4903 4525 4955 4531
rect 3323 4513 3329 4521
rect 4897 4513 4903 4521
rect 3323 4485 4903 4513
rect 3323 4478 3329 4485
rect 4897 4478 4903 4485
rect 3271 4467 3323 4473
rect 6535 4525 6587 4531
rect 4955 4513 4961 4521
rect 6529 4513 6535 4521
rect 4955 4485 6535 4513
rect 4955 4478 4961 4485
rect 6529 4478 6535 4485
rect 4903 4467 4955 4473
rect 8167 4525 8219 4531
rect 6587 4513 6593 4521
rect 8161 4513 8167 4521
rect 6587 4485 8167 4513
rect 6587 4478 6593 4485
rect 8161 4478 8167 4485
rect 6535 4467 6587 4473
rect 9799 4525 9851 4531
rect 8219 4513 8225 4521
rect 9793 4513 9799 4521
rect 8219 4485 9799 4513
rect 8219 4478 8225 4485
rect 9793 4478 9799 4485
rect 8167 4467 8219 4473
rect 9851 4478 9857 4521
rect 9799 4467 9851 4473
rect 212 4319 218 4371
rect 270 4359 276 4371
rect 416 4359 422 4371
rect 270 4331 422 4359
rect 270 4319 276 4331
rect 416 4319 422 4331
rect 474 4359 480 4371
rect 620 4359 626 4371
rect 474 4331 626 4359
rect 474 4319 480 4331
rect 620 4319 626 4331
rect 678 4359 684 4371
rect 824 4359 830 4371
rect 678 4331 830 4359
rect 678 4319 684 4331
rect 824 4319 830 4331
rect 882 4359 888 4371
rect 1028 4359 1034 4371
rect 882 4331 1034 4359
rect 882 4319 888 4331
rect 1028 4319 1034 4331
rect 1086 4359 1092 4371
rect 1232 4359 1238 4371
rect 1086 4331 1238 4359
rect 1086 4319 1092 4331
rect 1232 4319 1238 4331
rect 1290 4359 1296 4371
rect 1436 4359 1442 4371
rect 1290 4331 1442 4359
rect 1290 4319 1296 4331
rect 1436 4319 1442 4331
rect 1494 4359 1500 4371
rect 1640 4359 1646 4371
rect 1494 4331 1646 4359
rect 1494 4319 1500 4331
rect 1640 4319 1646 4331
rect 1698 4359 1704 4371
rect 1844 4359 1850 4371
rect 1698 4331 1850 4359
rect 1698 4319 1704 4331
rect 1844 4319 1850 4331
rect 1902 4359 1908 4371
rect 2048 4359 2054 4371
rect 1902 4331 2054 4359
rect 1902 4319 1908 4331
rect 2048 4319 2054 4331
rect 2106 4359 2112 4371
rect 2252 4359 2258 4371
rect 2106 4331 2258 4359
rect 2106 4319 2112 4331
rect 2252 4319 2258 4331
rect 2310 4359 2316 4371
rect 2456 4359 2462 4371
rect 2310 4331 2462 4359
rect 2310 4319 2316 4331
rect 2456 4319 2462 4331
rect 2514 4359 2520 4371
rect 2660 4359 2666 4371
rect 2514 4331 2666 4359
rect 2514 4319 2520 4331
rect 2660 4319 2666 4331
rect 2718 4359 2724 4371
rect 2864 4359 2870 4371
rect 2718 4331 2870 4359
rect 2718 4319 2724 4331
rect 2864 4319 2870 4331
rect 2922 4359 2928 4371
rect 3068 4359 3074 4371
rect 2922 4331 3074 4359
rect 2922 4319 2928 4331
rect 3068 4319 3074 4331
rect 3126 4359 3132 4371
rect 3272 4359 3278 4371
rect 3126 4331 3278 4359
rect 3126 4319 3132 4331
rect 3272 4319 3278 4331
rect 3330 4359 3336 4371
rect 3476 4359 3482 4371
rect 3330 4331 3482 4359
rect 3330 4319 3336 4331
rect 3476 4319 3482 4331
rect 3534 4359 3540 4371
rect 3680 4359 3686 4371
rect 3534 4331 3686 4359
rect 3534 4319 3540 4331
rect 3680 4319 3686 4331
rect 3738 4359 3744 4371
rect 3884 4359 3890 4371
rect 3738 4331 3890 4359
rect 3738 4319 3744 4331
rect 3884 4319 3890 4331
rect 3942 4359 3948 4371
rect 4088 4359 4094 4371
rect 3942 4331 4094 4359
rect 3942 4319 3948 4331
rect 4088 4319 4094 4331
rect 4146 4359 4152 4371
rect 4292 4359 4298 4371
rect 4146 4331 4298 4359
rect 4146 4319 4152 4331
rect 4292 4319 4298 4331
rect 4350 4359 4356 4371
rect 4496 4359 4502 4371
rect 4350 4331 4502 4359
rect 4350 4319 4356 4331
rect 4496 4319 4502 4331
rect 4554 4359 4560 4371
rect 4700 4359 4706 4371
rect 4554 4331 4706 4359
rect 4554 4319 4560 4331
rect 4700 4319 4706 4331
rect 4758 4359 4764 4371
rect 4904 4359 4910 4371
rect 4758 4331 4910 4359
rect 4758 4319 4764 4331
rect 4904 4319 4910 4331
rect 4962 4359 4968 4371
rect 5108 4359 5114 4371
rect 4962 4331 5114 4359
rect 4962 4319 4968 4331
rect 5108 4319 5114 4331
rect 5166 4359 5172 4371
rect 5312 4359 5318 4371
rect 5166 4331 5318 4359
rect 5166 4319 5172 4331
rect 5312 4319 5318 4331
rect 5370 4359 5376 4371
rect 5516 4359 5522 4371
rect 5370 4331 5522 4359
rect 5370 4319 5376 4331
rect 5516 4319 5522 4331
rect 5574 4359 5580 4371
rect 5720 4359 5726 4371
rect 5574 4331 5726 4359
rect 5574 4319 5580 4331
rect 5720 4319 5726 4331
rect 5778 4359 5784 4371
rect 5924 4359 5930 4371
rect 5778 4331 5930 4359
rect 5778 4319 5784 4331
rect 5924 4319 5930 4331
rect 5982 4359 5988 4371
rect 6128 4359 6134 4371
rect 5982 4331 6134 4359
rect 5982 4319 5988 4331
rect 6128 4319 6134 4331
rect 6186 4359 6192 4371
rect 6332 4359 6338 4371
rect 6186 4331 6338 4359
rect 6186 4319 6192 4331
rect 6332 4319 6338 4331
rect 6390 4359 6396 4371
rect 6536 4359 6542 4371
rect 6390 4331 6542 4359
rect 6390 4319 6396 4331
rect 6536 4319 6542 4331
rect 6594 4359 6600 4371
rect 6740 4359 6746 4371
rect 6594 4331 6746 4359
rect 6594 4319 6600 4331
rect 6740 4319 6746 4331
rect 6798 4359 6804 4371
rect 6944 4359 6950 4371
rect 6798 4331 6950 4359
rect 6798 4319 6804 4331
rect 6944 4319 6950 4331
rect 7002 4359 7008 4371
rect 7148 4359 7154 4371
rect 7002 4331 7154 4359
rect 7002 4319 7008 4331
rect 7148 4319 7154 4331
rect 7206 4359 7212 4371
rect 7352 4359 7358 4371
rect 7206 4331 7358 4359
rect 7206 4319 7212 4331
rect 7352 4319 7358 4331
rect 7410 4359 7416 4371
rect 7556 4359 7562 4371
rect 7410 4331 7562 4359
rect 7410 4319 7416 4331
rect 7556 4319 7562 4331
rect 7614 4359 7620 4371
rect 7760 4359 7766 4371
rect 7614 4331 7766 4359
rect 7614 4319 7620 4331
rect 7760 4319 7766 4331
rect 7818 4359 7824 4371
rect 7964 4359 7970 4371
rect 7818 4331 7970 4359
rect 7818 4319 7824 4331
rect 7964 4319 7970 4331
rect 8022 4359 8028 4371
rect 8168 4359 8174 4371
rect 8022 4331 8174 4359
rect 8022 4319 8028 4331
rect 8168 4319 8174 4331
rect 8226 4359 8232 4371
rect 8372 4359 8378 4371
rect 8226 4331 8378 4359
rect 8226 4319 8232 4331
rect 8372 4319 8378 4331
rect 8430 4359 8436 4371
rect 8576 4359 8582 4371
rect 8430 4331 8582 4359
rect 8430 4319 8436 4331
rect 8576 4319 8582 4331
rect 8634 4359 8640 4371
rect 8780 4359 8786 4371
rect 8634 4331 8786 4359
rect 8634 4319 8640 4331
rect 8780 4319 8786 4331
rect 8838 4359 8844 4371
rect 8984 4359 8990 4371
rect 8838 4331 8990 4359
rect 8838 4319 8844 4331
rect 8984 4319 8990 4331
rect 9042 4359 9048 4371
rect 9188 4359 9194 4371
rect 9042 4331 9194 4359
rect 9042 4319 9048 4331
rect 9188 4319 9194 4331
rect 9246 4359 9252 4371
rect 9392 4359 9398 4371
rect 9246 4331 9398 4359
rect 9246 4319 9252 4331
rect 9392 4319 9398 4331
rect 9450 4359 9456 4371
rect 9596 4359 9602 4371
rect 9450 4331 9602 4359
rect 9450 4319 9456 4331
rect 9596 4319 9602 4331
rect 9654 4359 9660 4371
rect 9814 4359 9820 4371
rect 9654 4331 9820 4359
rect 9654 4319 9660 4331
rect 9814 4319 9820 4331
rect 9872 4319 9878 4371
rect 7 4217 59 4223
rect 1 4170 7 4213
rect 1639 4217 1691 4223
rect 59 4205 65 4213
rect 1633 4205 1639 4213
rect 59 4177 1639 4205
rect 59 4170 65 4177
rect 1633 4170 1639 4177
rect 7 4159 59 4165
rect 3271 4217 3323 4223
rect 1691 4205 1697 4213
rect 3265 4205 3271 4213
rect 1691 4177 3271 4205
rect 1691 4170 1697 4177
rect 3265 4170 3271 4177
rect 1639 4159 1691 4165
rect 4903 4217 4955 4223
rect 3323 4205 3329 4213
rect 4897 4205 4903 4213
rect 3323 4177 4903 4205
rect 3323 4170 3329 4177
rect 4897 4170 4903 4177
rect 3271 4159 3323 4165
rect 6535 4217 6587 4223
rect 4955 4205 4961 4213
rect 6529 4205 6535 4213
rect 4955 4177 6535 4205
rect 4955 4170 4961 4177
rect 6529 4170 6535 4177
rect 4903 4159 4955 4165
rect 8167 4217 8219 4223
rect 6587 4205 6593 4213
rect 8161 4205 8167 4213
rect 6587 4177 8167 4205
rect 6587 4170 6593 4177
rect 8161 4170 8167 4177
rect 6535 4159 6587 4165
rect 9799 4217 9851 4223
rect 8219 4205 8225 4213
rect 9793 4205 9799 4213
rect 8219 4177 9799 4205
rect 8219 4170 8225 4177
rect 9793 4170 9799 4177
rect 8167 4159 8219 4165
rect 9851 4170 9857 4213
rect 9799 4159 9851 4165
rect 7 4013 59 4019
rect 1 3966 7 4009
rect 1639 4013 1691 4019
rect 59 4001 65 4009
rect 1633 4001 1639 4009
rect 59 3973 1639 4001
rect 59 3966 65 3973
rect 1633 3966 1639 3973
rect 7 3955 59 3961
rect 3271 4013 3323 4019
rect 1691 4001 1697 4009
rect 3265 4001 3271 4009
rect 1691 3973 3271 4001
rect 1691 3966 1697 3973
rect 3265 3966 3271 3973
rect 1639 3955 1691 3961
rect 4903 4013 4955 4019
rect 3323 4001 3329 4009
rect 4897 4001 4903 4009
rect 3323 3973 4903 4001
rect 3323 3966 3329 3973
rect 4897 3966 4903 3973
rect 3271 3955 3323 3961
rect 6535 4013 6587 4019
rect 4955 4001 4961 4009
rect 6529 4001 6535 4009
rect 4955 3973 6535 4001
rect 4955 3966 4961 3973
rect 6529 3966 6535 3973
rect 4903 3955 4955 3961
rect 8167 4013 8219 4019
rect 6587 4001 6593 4009
rect 8161 4001 8167 4009
rect 6587 3973 8167 4001
rect 6587 3966 6593 3973
rect 8161 3966 8167 3973
rect 6535 3955 6587 3961
rect 9799 4013 9851 4019
rect 8219 4001 8225 4009
rect 9793 4001 9799 4009
rect 8219 3973 9799 4001
rect 8219 3966 8225 3973
rect 9793 3966 9799 3973
rect 8167 3955 8219 3961
rect 9851 3966 9857 4009
rect 9799 3955 9851 3961
rect 7 3809 59 3815
rect 1 3762 7 3805
rect 1639 3809 1691 3815
rect 59 3797 65 3805
rect 1633 3797 1639 3805
rect 59 3769 1639 3797
rect 59 3762 65 3769
rect 1633 3762 1639 3769
rect 7 3751 59 3757
rect 3271 3809 3323 3815
rect 1691 3797 1697 3805
rect 3265 3797 3271 3805
rect 1691 3769 3271 3797
rect 1691 3762 1697 3769
rect 3265 3762 3271 3769
rect 1639 3751 1691 3757
rect 4903 3809 4955 3815
rect 3323 3797 3329 3805
rect 4897 3797 4903 3805
rect 3323 3769 4903 3797
rect 3323 3762 3329 3769
rect 4897 3762 4903 3769
rect 3271 3751 3323 3757
rect 6535 3809 6587 3815
rect 4955 3797 4961 3805
rect 6529 3797 6535 3805
rect 4955 3769 6535 3797
rect 4955 3762 4961 3769
rect 6529 3762 6535 3769
rect 4903 3751 4955 3757
rect 8167 3809 8219 3815
rect 6587 3797 6593 3805
rect 8161 3797 8167 3805
rect 6587 3769 8167 3797
rect 6587 3762 6593 3769
rect 8161 3762 8167 3769
rect 6535 3751 6587 3757
rect 9799 3809 9851 3815
rect 8219 3797 8225 3805
rect 9793 3797 9799 3805
rect 8219 3769 9799 3797
rect 8219 3762 8225 3769
rect 9793 3762 9799 3769
rect 8167 3751 8219 3757
rect 9851 3762 9857 3805
rect 9799 3751 9851 3757
rect 7 3605 59 3611
rect 1 3558 7 3601
rect 1639 3605 1691 3611
rect 59 3593 65 3601
rect 1633 3593 1639 3601
rect 59 3565 1639 3593
rect 59 3558 65 3565
rect 1633 3558 1639 3565
rect 7 3547 59 3553
rect 3271 3605 3323 3611
rect 1691 3593 1697 3601
rect 3265 3593 3271 3601
rect 1691 3565 3271 3593
rect 1691 3558 1697 3565
rect 3265 3558 3271 3565
rect 1639 3547 1691 3553
rect 4903 3605 4955 3611
rect 3323 3593 3329 3601
rect 4897 3593 4903 3601
rect 3323 3565 4903 3593
rect 3323 3558 3329 3565
rect 4897 3558 4903 3565
rect 3271 3547 3323 3553
rect 6535 3605 6587 3611
rect 4955 3593 4961 3601
rect 6529 3593 6535 3601
rect 4955 3565 6535 3593
rect 4955 3558 4961 3565
rect 6529 3558 6535 3565
rect 4903 3547 4955 3553
rect 8167 3605 8219 3611
rect 6587 3593 6593 3601
rect 8161 3593 8167 3601
rect 6587 3565 8167 3593
rect 6587 3558 6593 3565
rect 8161 3558 8167 3565
rect 6535 3547 6587 3553
rect 9799 3605 9851 3611
rect 8219 3593 8225 3601
rect 9793 3593 9799 3601
rect 8219 3565 9799 3593
rect 8219 3558 8225 3565
rect 9793 3558 9799 3565
rect 8167 3547 8219 3553
rect 9851 3558 9857 3601
rect 9799 3547 9851 3553
rect 7 3401 59 3407
rect 1 3354 7 3397
rect 1639 3401 1691 3407
rect 59 3389 65 3397
rect 1633 3389 1639 3397
rect 59 3361 1639 3389
rect 59 3354 65 3361
rect 1633 3354 1639 3361
rect 7 3343 59 3349
rect 3271 3401 3323 3407
rect 1691 3389 1697 3397
rect 3265 3389 3271 3397
rect 1691 3361 3271 3389
rect 1691 3354 1697 3361
rect 3265 3354 3271 3361
rect 1639 3343 1691 3349
rect 4903 3401 4955 3407
rect 3323 3389 3329 3397
rect 4897 3389 4903 3397
rect 3323 3361 4903 3389
rect 3323 3354 3329 3361
rect 4897 3354 4903 3361
rect 3271 3343 3323 3349
rect 6535 3401 6587 3407
rect 4955 3389 4961 3397
rect 6529 3389 6535 3397
rect 4955 3361 6535 3389
rect 4955 3354 4961 3361
rect 6529 3354 6535 3361
rect 4903 3343 4955 3349
rect 8167 3401 8219 3407
rect 6587 3389 6593 3397
rect 8161 3389 8167 3397
rect 6587 3361 8167 3389
rect 6587 3354 6593 3361
rect 8161 3354 8167 3361
rect 6535 3343 6587 3349
rect 9799 3401 9851 3407
rect 8219 3389 8225 3397
rect 9793 3389 9799 3397
rect 8219 3361 9799 3389
rect 8219 3354 8225 3361
rect 9793 3354 9799 3361
rect 8167 3343 8219 3349
rect 9851 3354 9857 3397
rect 9799 3343 9851 3349
rect 7 3197 59 3203
rect 1 3150 7 3193
rect 1639 3197 1691 3203
rect 59 3185 65 3193
rect 1633 3185 1639 3193
rect 59 3157 1639 3185
rect 59 3150 65 3157
rect 1633 3150 1639 3157
rect 7 3139 59 3145
rect 3271 3197 3323 3203
rect 1691 3185 1697 3193
rect 3265 3185 3271 3193
rect 1691 3157 3271 3185
rect 1691 3150 1697 3157
rect 3265 3150 3271 3157
rect 1639 3139 1691 3145
rect 4903 3197 4955 3203
rect 3323 3185 3329 3193
rect 4897 3185 4903 3193
rect 3323 3157 4903 3185
rect 3323 3150 3329 3157
rect 4897 3150 4903 3157
rect 3271 3139 3323 3145
rect 6535 3197 6587 3203
rect 4955 3185 4961 3193
rect 6529 3185 6535 3193
rect 4955 3157 6535 3185
rect 4955 3150 4961 3157
rect 6529 3150 6535 3157
rect 4903 3139 4955 3145
rect 8167 3197 8219 3203
rect 6587 3185 6593 3193
rect 8161 3185 8167 3193
rect 6587 3157 8167 3185
rect 6587 3150 6593 3157
rect 8161 3150 8167 3157
rect 6535 3139 6587 3145
rect 9799 3197 9851 3203
rect 8219 3185 8225 3193
rect 9793 3185 9799 3193
rect 8219 3157 9799 3185
rect 8219 3150 8225 3157
rect 9793 3150 9799 3157
rect 8167 3139 8219 3145
rect 9851 3150 9857 3193
rect 9799 3139 9851 3145
rect 7 2993 59 2999
rect 1 2946 7 2989
rect 1639 2993 1691 2999
rect 59 2981 65 2989
rect 1633 2981 1639 2989
rect 59 2953 1639 2981
rect 59 2946 65 2953
rect 1633 2946 1639 2953
rect 7 2935 59 2941
rect 3271 2993 3323 2999
rect 1691 2981 1697 2989
rect 3265 2981 3271 2989
rect 1691 2953 3271 2981
rect 1691 2946 1697 2953
rect 3265 2946 3271 2953
rect 1639 2935 1691 2941
rect 4903 2993 4955 2999
rect 3323 2981 3329 2989
rect 4897 2981 4903 2989
rect 3323 2953 4903 2981
rect 3323 2946 3329 2953
rect 4897 2946 4903 2953
rect 3271 2935 3323 2941
rect 6535 2993 6587 2999
rect 4955 2981 4961 2989
rect 6529 2981 6535 2989
rect 4955 2953 6535 2981
rect 4955 2946 4961 2953
rect 6529 2946 6535 2953
rect 4903 2935 4955 2941
rect 8167 2993 8219 2999
rect 6587 2981 6593 2989
rect 8161 2981 8167 2989
rect 6587 2953 8167 2981
rect 6587 2946 6593 2953
rect 8161 2946 8167 2953
rect 6535 2935 6587 2941
rect 9799 2993 9851 2999
rect 8219 2981 8225 2989
rect 9793 2981 9799 2989
rect 8219 2953 9799 2981
rect 8219 2946 8225 2953
rect 9793 2946 9799 2953
rect 8167 2935 8219 2941
rect 9851 2946 9857 2989
rect 9799 2935 9851 2941
rect 7 2789 59 2795
rect 1 2742 7 2785
rect 1639 2789 1691 2795
rect 59 2777 65 2785
rect 1633 2777 1639 2785
rect 59 2749 1639 2777
rect 59 2742 65 2749
rect 1633 2742 1639 2749
rect 7 2731 59 2737
rect 3271 2789 3323 2795
rect 1691 2777 1697 2785
rect 3265 2777 3271 2785
rect 1691 2749 3271 2777
rect 1691 2742 1697 2749
rect 3265 2742 3271 2749
rect 1639 2731 1691 2737
rect 4903 2789 4955 2795
rect 3323 2777 3329 2785
rect 4897 2777 4903 2785
rect 3323 2749 4903 2777
rect 3323 2742 3329 2749
rect 4897 2742 4903 2749
rect 3271 2731 3323 2737
rect 6535 2789 6587 2795
rect 4955 2777 4961 2785
rect 6529 2777 6535 2785
rect 4955 2749 6535 2777
rect 4955 2742 4961 2749
rect 6529 2742 6535 2749
rect 4903 2731 4955 2737
rect 8167 2789 8219 2795
rect 6587 2777 6593 2785
rect 8161 2777 8167 2785
rect 6587 2749 8167 2777
rect 6587 2742 6593 2749
rect 8161 2742 8167 2749
rect 6535 2731 6587 2737
rect 9799 2789 9851 2795
rect 8219 2777 8225 2785
rect 9793 2777 9799 2785
rect 8219 2749 9799 2777
rect 8219 2742 8225 2749
rect 9793 2742 9799 2749
rect 8167 2731 8219 2737
rect 9851 2742 9857 2785
rect 9799 2731 9851 2737
rect 212 2583 218 2635
rect 270 2623 276 2635
rect 416 2623 422 2635
rect 270 2595 422 2623
rect 270 2583 276 2595
rect 416 2583 422 2595
rect 474 2623 480 2635
rect 620 2623 626 2635
rect 474 2595 626 2623
rect 474 2583 480 2595
rect 620 2583 626 2595
rect 678 2623 684 2635
rect 824 2623 830 2635
rect 678 2595 830 2623
rect 678 2583 684 2595
rect 824 2583 830 2595
rect 882 2623 888 2635
rect 1028 2623 1034 2635
rect 882 2595 1034 2623
rect 882 2583 888 2595
rect 1028 2583 1034 2595
rect 1086 2623 1092 2635
rect 1232 2623 1238 2635
rect 1086 2595 1238 2623
rect 1086 2583 1092 2595
rect 1232 2583 1238 2595
rect 1290 2623 1296 2635
rect 1436 2623 1442 2635
rect 1290 2595 1442 2623
rect 1290 2583 1296 2595
rect 1436 2583 1442 2595
rect 1494 2623 1500 2635
rect 1640 2623 1646 2635
rect 1494 2595 1646 2623
rect 1494 2583 1500 2595
rect 1640 2583 1646 2595
rect 1698 2623 1704 2635
rect 1844 2623 1850 2635
rect 1698 2595 1850 2623
rect 1698 2583 1704 2595
rect 1844 2583 1850 2595
rect 1902 2623 1908 2635
rect 2048 2623 2054 2635
rect 1902 2595 2054 2623
rect 1902 2583 1908 2595
rect 2048 2583 2054 2595
rect 2106 2623 2112 2635
rect 2252 2623 2258 2635
rect 2106 2595 2258 2623
rect 2106 2583 2112 2595
rect 2252 2583 2258 2595
rect 2310 2623 2316 2635
rect 2456 2623 2462 2635
rect 2310 2595 2462 2623
rect 2310 2583 2316 2595
rect 2456 2583 2462 2595
rect 2514 2623 2520 2635
rect 2660 2623 2666 2635
rect 2514 2595 2666 2623
rect 2514 2583 2520 2595
rect 2660 2583 2666 2595
rect 2718 2623 2724 2635
rect 2864 2623 2870 2635
rect 2718 2595 2870 2623
rect 2718 2583 2724 2595
rect 2864 2583 2870 2595
rect 2922 2623 2928 2635
rect 3068 2623 3074 2635
rect 2922 2595 3074 2623
rect 2922 2583 2928 2595
rect 3068 2583 3074 2595
rect 3126 2623 3132 2635
rect 3272 2623 3278 2635
rect 3126 2595 3278 2623
rect 3126 2583 3132 2595
rect 3272 2583 3278 2595
rect 3330 2623 3336 2635
rect 3476 2623 3482 2635
rect 3330 2595 3482 2623
rect 3330 2583 3336 2595
rect 3476 2583 3482 2595
rect 3534 2623 3540 2635
rect 3680 2623 3686 2635
rect 3534 2595 3686 2623
rect 3534 2583 3540 2595
rect 3680 2583 3686 2595
rect 3738 2623 3744 2635
rect 3884 2623 3890 2635
rect 3738 2595 3890 2623
rect 3738 2583 3744 2595
rect 3884 2583 3890 2595
rect 3942 2623 3948 2635
rect 4088 2623 4094 2635
rect 3942 2595 4094 2623
rect 3942 2583 3948 2595
rect 4088 2583 4094 2595
rect 4146 2623 4152 2635
rect 4292 2623 4298 2635
rect 4146 2595 4298 2623
rect 4146 2583 4152 2595
rect 4292 2583 4298 2595
rect 4350 2623 4356 2635
rect 4496 2623 4502 2635
rect 4350 2595 4502 2623
rect 4350 2583 4356 2595
rect 4496 2583 4502 2595
rect 4554 2623 4560 2635
rect 4700 2623 4706 2635
rect 4554 2595 4706 2623
rect 4554 2583 4560 2595
rect 4700 2583 4706 2595
rect 4758 2623 4764 2635
rect 4904 2623 4910 2635
rect 4758 2595 4910 2623
rect 4758 2583 4764 2595
rect 4904 2583 4910 2595
rect 4962 2623 4968 2635
rect 5108 2623 5114 2635
rect 4962 2595 5114 2623
rect 4962 2583 4968 2595
rect 5108 2583 5114 2595
rect 5166 2623 5172 2635
rect 5312 2623 5318 2635
rect 5166 2595 5318 2623
rect 5166 2583 5172 2595
rect 5312 2583 5318 2595
rect 5370 2623 5376 2635
rect 5516 2623 5522 2635
rect 5370 2595 5522 2623
rect 5370 2583 5376 2595
rect 5516 2583 5522 2595
rect 5574 2623 5580 2635
rect 5720 2623 5726 2635
rect 5574 2595 5726 2623
rect 5574 2583 5580 2595
rect 5720 2583 5726 2595
rect 5778 2623 5784 2635
rect 5924 2623 5930 2635
rect 5778 2595 5930 2623
rect 5778 2583 5784 2595
rect 5924 2583 5930 2595
rect 5982 2623 5988 2635
rect 6128 2623 6134 2635
rect 5982 2595 6134 2623
rect 5982 2583 5988 2595
rect 6128 2583 6134 2595
rect 6186 2623 6192 2635
rect 6332 2623 6338 2635
rect 6186 2595 6338 2623
rect 6186 2583 6192 2595
rect 6332 2583 6338 2595
rect 6390 2623 6396 2635
rect 6536 2623 6542 2635
rect 6390 2595 6542 2623
rect 6390 2583 6396 2595
rect 6536 2583 6542 2595
rect 6594 2623 6600 2635
rect 6740 2623 6746 2635
rect 6594 2595 6746 2623
rect 6594 2583 6600 2595
rect 6740 2583 6746 2595
rect 6798 2623 6804 2635
rect 6944 2623 6950 2635
rect 6798 2595 6950 2623
rect 6798 2583 6804 2595
rect 6944 2583 6950 2595
rect 7002 2623 7008 2635
rect 7148 2623 7154 2635
rect 7002 2595 7154 2623
rect 7002 2583 7008 2595
rect 7148 2583 7154 2595
rect 7206 2623 7212 2635
rect 7352 2623 7358 2635
rect 7206 2595 7358 2623
rect 7206 2583 7212 2595
rect 7352 2583 7358 2595
rect 7410 2623 7416 2635
rect 7556 2623 7562 2635
rect 7410 2595 7562 2623
rect 7410 2583 7416 2595
rect 7556 2583 7562 2595
rect 7614 2623 7620 2635
rect 7760 2623 7766 2635
rect 7614 2595 7766 2623
rect 7614 2583 7620 2595
rect 7760 2583 7766 2595
rect 7818 2623 7824 2635
rect 7964 2623 7970 2635
rect 7818 2595 7970 2623
rect 7818 2583 7824 2595
rect 7964 2583 7970 2595
rect 8022 2623 8028 2635
rect 8168 2623 8174 2635
rect 8022 2595 8174 2623
rect 8022 2583 8028 2595
rect 8168 2583 8174 2595
rect 8226 2623 8232 2635
rect 8372 2623 8378 2635
rect 8226 2595 8378 2623
rect 8226 2583 8232 2595
rect 8372 2583 8378 2595
rect 8430 2623 8436 2635
rect 8576 2623 8582 2635
rect 8430 2595 8582 2623
rect 8430 2583 8436 2595
rect 8576 2583 8582 2595
rect 8634 2623 8640 2635
rect 8780 2623 8786 2635
rect 8634 2595 8786 2623
rect 8634 2583 8640 2595
rect 8780 2583 8786 2595
rect 8838 2623 8844 2635
rect 8984 2623 8990 2635
rect 8838 2595 8990 2623
rect 8838 2583 8844 2595
rect 8984 2583 8990 2595
rect 9042 2623 9048 2635
rect 9188 2623 9194 2635
rect 9042 2595 9194 2623
rect 9042 2583 9048 2595
rect 9188 2583 9194 2595
rect 9246 2623 9252 2635
rect 9392 2623 9398 2635
rect 9246 2595 9398 2623
rect 9246 2583 9252 2595
rect 9392 2583 9398 2595
rect 9450 2623 9456 2635
rect 9596 2623 9602 2635
rect 9450 2595 9602 2623
rect 9450 2583 9456 2595
rect 9596 2583 9602 2595
rect 9654 2623 9660 2635
rect 9814 2623 9820 2635
rect 9654 2595 9820 2623
rect 9654 2583 9660 2595
rect 9814 2583 9820 2595
rect 9872 2583 9878 2635
rect 7 2481 59 2487
rect 1 2434 7 2477
rect 1639 2481 1691 2487
rect 59 2469 65 2477
rect 1633 2469 1639 2477
rect 59 2441 1639 2469
rect 59 2434 65 2441
rect 1633 2434 1639 2441
rect 7 2423 59 2429
rect 3271 2481 3323 2487
rect 1691 2469 1697 2477
rect 3265 2469 3271 2477
rect 1691 2441 3271 2469
rect 1691 2434 1697 2441
rect 3265 2434 3271 2441
rect 1639 2423 1691 2429
rect 4903 2481 4955 2487
rect 3323 2469 3329 2477
rect 4897 2469 4903 2477
rect 3323 2441 4903 2469
rect 3323 2434 3329 2441
rect 4897 2434 4903 2441
rect 3271 2423 3323 2429
rect 6535 2481 6587 2487
rect 4955 2469 4961 2477
rect 6529 2469 6535 2477
rect 4955 2441 6535 2469
rect 4955 2434 4961 2441
rect 6529 2434 6535 2441
rect 4903 2423 4955 2429
rect 8167 2481 8219 2487
rect 6587 2469 6593 2477
rect 8161 2469 8167 2477
rect 6587 2441 8167 2469
rect 6587 2434 6593 2441
rect 8161 2434 8167 2441
rect 6535 2423 6587 2429
rect 9799 2481 9851 2487
rect 8219 2469 8225 2477
rect 9793 2469 9799 2477
rect 8219 2441 9799 2469
rect 8219 2434 8225 2441
rect 9793 2434 9799 2441
rect 8167 2423 8219 2429
rect 9851 2434 9857 2477
rect 9799 2423 9851 2429
rect 7 2277 59 2283
rect 1 2230 7 2273
rect 1639 2277 1691 2283
rect 59 2265 65 2273
rect 1633 2265 1639 2273
rect 59 2237 1639 2265
rect 59 2230 65 2237
rect 1633 2230 1639 2237
rect 7 2219 59 2225
rect 3271 2277 3323 2283
rect 1691 2265 1697 2273
rect 3265 2265 3271 2273
rect 1691 2237 3271 2265
rect 1691 2230 1697 2237
rect 3265 2230 3271 2237
rect 1639 2219 1691 2225
rect 4903 2277 4955 2283
rect 3323 2265 3329 2273
rect 4897 2265 4903 2273
rect 3323 2237 4903 2265
rect 3323 2230 3329 2237
rect 4897 2230 4903 2237
rect 3271 2219 3323 2225
rect 6535 2277 6587 2283
rect 4955 2265 4961 2273
rect 6529 2265 6535 2273
rect 4955 2237 6535 2265
rect 4955 2230 4961 2237
rect 6529 2230 6535 2237
rect 4903 2219 4955 2225
rect 8167 2277 8219 2283
rect 6587 2265 6593 2273
rect 8161 2265 8167 2273
rect 6587 2237 8167 2265
rect 6587 2230 6593 2237
rect 8161 2230 8167 2237
rect 6535 2219 6587 2225
rect 9799 2277 9851 2283
rect 8219 2265 8225 2273
rect 9793 2265 9799 2273
rect 8219 2237 9799 2265
rect 8219 2230 8225 2237
rect 9793 2230 9799 2237
rect 8167 2219 8219 2225
rect 9851 2230 9857 2273
rect 9799 2219 9851 2225
rect 7 2073 59 2079
rect 1 2026 7 2069
rect 1639 2073 1691 2079
rect 59 2061 65 2069
rect 1633 2061 1639 2069
rect 59 2033 1639 2061
rect 59 2026 65 2033
rect 1633 2026 1639 2033
rect 7 2015 59 2021
rect 3271 2073 3323 2079
rect 1691 2061 1697 2069
rect 3265 2061 3271 2069
rect 1691 2033 3271 2061
rect 1691 2026 1697 2033
rect 3265 2026 3271 2033
rect 1639 2015 1691 2021
rect 4903 2073 4955 2079
rect 3323 2061 3329 2069
rect 4897 2061 4903 2069
rect 3323 2033 4903 2061
rect 3323 2026 3329 2033
rect 4897 2026 4903 2033
rect 3271 2015 3323 2021
rect 6535 2073 6587 2079
rect 4955 2061 4961 2069
rect 6529 2061 6535 2069
rect 4955 2033 6535 2061
rect 4955 2026 4961 2033
rect 6529 2026 6535 2033
rect 4903 2015 4955 2021
rect 8167 2073 8219 2079
rect 6587 2061 6593 2069
rect 8161 2061 8167 2069
rect 6587 2033 8167 2061
rect 6587 2026 6593 2033
rect 8161 2026 8167 2033
rect 6535 2015 6587 2021
rect 9799 2073 9851 2079
rect 8219 2061 8225 2069
rect 9793 2061 9799 2069
rect 8219 2033 9799 2061
rect 8219 2026 8225 2033
rect 9793 2026 9799 2033
rect 8167 2015 8219 2021
rect 9851 2026 9857 2069
rect 9799 2015 9851 2021
rect 7 1869 59 1875
rect 1 1822 7 1865
rect 1639 1869 1691 1875
rect 59 1857 65 1865
rect 1633 1857 1639 1865
rect 59 1829 1639 1857
rect 59 1822 65 1829
rect 1633 1822 1639 1829
rect 7 1811 59 1817
rect 3271 1869 3323 1875
rect 1691 1857 1697 1865
rect 3265 1857 3271 1865
rect 1691 1829 3271 1857
rect 1691 1822 1697 1829
rect 3265 1822 3271 1829
rect 1639 1811 1691 1817
rect 4903 1869 4955 1875
rect 3323 1857 3329 1865
rect 4897 1857 4903 1865
rect 3323 1829 4903 1857
rect 3323 1822 3329 1829
rect 4897 1822 4903 1829
rect 3271 1811 3323 1817
rect 6535 1869 6587 1875
rect 4955 1857 4961 1865
rect 6529 1857 6535 1865
rect 4955 1829 6535 1857
rect 4955 1822 4961 1829
rect 6529 1822 6535 1829
rect 4903 1811 4955 1817
rect 8167 1869 8219 1875
rect 6587 1857 6593 1865
rect 8161 1857 8167 1865
rect 6587 1829 8167 1857
rect 6587 1822 6593 1829
rect 8161 1822 8167 1829
rect 6535 1811 6587 1817
rect 9799 1869 9851 1875
rect 8219 1857 8225 1865
rect 9793 1857 9799 1865
rect 8219 1829 9799 1857
rect 8219 1822 8225 1829
rect 9793 1822 9799 1829
rect 8167 1811 8219 1817
rect 9851 1822 9857 1865
rect 9799 1811 9851 1817
rect 7 1665 59 1671
rect 1 1618 7 1661
rect 1639 1665 1691 1671
rect 59 1653 65 1661
rect 1633 1653 1639 1661
rect 59 1625 1639 1653
rect 59 1618 65 1625
rect 1633 1618 1639 1625
rect 7 1607 59 1613
rect 3271 1665 3323 1671
rect 1691 1653 1697 1661
rect 3265 1653 3271 1661
rect 1691 1625 3271 1653
rect 1691 1618 1697 1625
rect 3265 1618 3271 1625
rect 1639 1607 1691 1613
rect 4903 1665 4955 1671
rect 3323 1653 3329 1661
rect 4897 1653 4903 1661
rect 3323 1625 4903 1653
rect 3323 1618 3329 1625
rect 4897 1618 4903 1625
rect 3271 1607 3323 1613
rect 6535 1665 6587 1671
rect 4955 1653 4961 1661
rect 6529 1653 6535 1661
rect 4955 1625 6535 1653
rect 4955 1618 4961 1625
rect 6529 1618 6535 1625
rect 4903 1607 4955 1613
rect 8167 1665 8219 1671
rect 6587 1653 6593 1661
rect 8161 1653 8167 1661
rect 6587 1625 8167 1653
rect 6587 1618 6593 1625
rect 8161 1618 8167 1625
rect 6535 1607 6587 1613
rect 9799 1665 9851 1671
rect 8219 1653 8225 1661
rect 9793 1653 9799 1661
rect 8219 1625 9799 1653
rect 8219 1618 8225 1625
rect 9793 1618 9799 1625
rect 8167 1607 8219 1613
rect 9851 1618 9857 1661
rect 9799 1607 9851 1613
rect 7 1461 59 1467
rect 1 1414 7 1457
rect 1639 1461 1691 1467
rect 59 1449 65 1457
rect 1633 1449 1639 1457
rect 59 1421 1639 1449
rect 59 1414 65 1421
rect 1633 1414 1639 1421
rect 7 1403 59 1409
rect 3271 1461 3323 1467
rect 1691 1449 1697 1457
rect 3265 1449 3271 1457
rect 1691 1421 3271 1449
rect 1691 1414 1697 1421
rect 3265 1414 3271 1421
rect 1639 1403 1691 1409
rect 4903 1461 4955 1467
rect 3323 1449 3329 1457
rect 4897 1449 4903 1457
rect 3323 1421 4903 1449
rect 3323 1414 3329 1421
rect 4897 1414 4903 1421
rect 3271 1403 3323 1409
rect 6535 1461 6587 1467
rect 4955 1449 4961 1457
rect 6529 1449 6535 1457
rect 4955 1421 6535 1449
rect 4955 1414 4961 1421
rect 6529 1414 6535 1421
rect 4903 1403 4955 1409
rect 8167 1461 8219 1467
rect 6587 1449 6593 1457
rect 8161 1449 8167 1457
rect 6587 1421 8167 1449
rect 6587 1414 6593 1421
rect 8161 1414 8167 1421
rect 6535 1403 6587 1409
rect 9799 1461 9851 1467
rect 8219 1449 8225 1457
rect 9793 1449 9799 1457
rect 8219 1421 9799 1449
rect 8219 1414 8225 1421
rect 9793 1414 9799 1421
rect 8167 1403 8219 1409
rect 9851 1414 9857 1457
rect 9799 1403 9851 1409
rect 7 1257 59 1263
rect 1 1210 7 1253
rect 1639 1257 1691 1263
rect 59 1245 65 1253
rect 1633 1245 1639 1253
rect 59 1217 1639 1245
rect 59 1210 65 1217
rect 1633 1210 1639 1217
rect 7 1199 59 1205
rect 3271 1257 3323 1263
rect 1691 1245 1697 1253
rect 3265 1245 3271 1253
rect 1691 1217 3271 1245
rect 1691 1210 1697 1217
rect 3265 1210 3271 1217
rect 1639 1199 1691 1205
rect 4903 1257 4955 1263
rect 3323 1245 3329 1253
rect 4897 1245 4903 1253
rect 3323 1217 4903 1245
rect 3323 1210 3329 1217
rect 4897 1210 4903 1217
rect 3271 1199 3323 1205
rect 6535 1257 6587 1263
rect 4955 1245 4961 1253
rect 6529 1245 6535 1253
rect 4955 1217 6535 1245
rect 4955 1210 4961 1217
rect 6529 1210 6535 1217
rect 4903 1199 4955 1205
rect 8167 1257 8219 1263
rect 6587 1245 6593 1253
rect 8161 1245 8167 1253
rect 6587 1217 8167 1245
rect 6587 1210 6593 1217
rect 8161 1210 8167 1217
rect 6535 1199 6587 1205
rect 9799 1257 9851 1263
rect 8219 1245 8225 1253
rect 9793 1245 9799 1253
rect 8219 1217 9799 1245
rect 8219 1210 8225 1217
rect 9793 1210 9799 1217
rect 8167 1199 8219 1205
rect 9851 1210 9857 1253
rect 9799 1199 9851 1205
rect 7 1053 59 1059
rect 1 1006 7 1049
rect 1639 1053 1691 1059
rect 59 1041 65 1049
rect 1633 1041 1639 1049
rect 59 1013 1639 1041
rect 59 1006 65 1013
rect 1633 1006 1639 1013
rect 7 995 59 1001
rect 3271 1053 3323 1059
rect 1691 1041 1697 1049
rect 3265 1041 3271 1049
rect 1691 1013 3271 1041
rect 1691 1006 1697 1013
rect 3265 1006 3271 1013
rect 1639 995 1691 1001
rect 4903 1053 4955 1059
rect 3323 1041 3329 1049
rect 4897 1041 4903 1049
rect 3323 1013 4903 1041
rect 3323 1006 3329 1013
rect 4897 1006 4903 1013
rect 3271 995 3323 1001
rect 6535 1053 6587 1059
rect 4955 1041 4961 1049
rect 6529 1041 6535 1049
rect 4955 1013 6535 1041
rect 4955 1006 4961 1013
rect 6529 1006 6535 1013
rect 4903 995 4955 1001
rect 8167 1053 8219 1059
rect 6587 1041 6593 1049
rect 8161 1041 8167 1049
rect 6587 1013 8167 1041
rect 6587 1006 6593 1013
rect 8161 1006 8167 1013
rect 6535 995 6587 1001
rect 9799 1053 9851 1059
rect 8219 1041 8225 1049
rect 9793 1041 9799 1049
rect 8219 1013 9799 1041
rect 8219 1006 8225 1013
rect 9793 1006 9799 1013
rect 8167 995 8219 1001
rect 9851 1006 9857 1049
rect 9799 995 9851 1001
rect 212 847 218 899
rect 270 887 276 899
rect 416 887 422 899
rect 270 859 422 887
rect 270 847 276 859
rect 416 847 422 859
rect 474 887 480 899
rect 620 887 626 899
rect 474 859 626 887
rect 474 847 480 859
rect 620 847 626 859
rect 678 887 684 899
rect 824 887 830 899
rect 678 859 830 887
rect 678 847 684 859
rect 824 847 830 859
rect 882 887 888 899
rect 1028 887 1034 899
rect 882 859 1034 887
rect 882 847 888 859
rect 1028 847 1034 859
rect 1086 887 1092 899
rect 1232 887 1238 899
rect 1086 859 1238 887
rect 1086 847 1092 859
rect 1232 847 1238 859
rect 1290 887 1296 899
rect 1436 887 1442 899
rect 1290 859 1442 887
rect 1290 847 1296 859
rect 1436 847 1442 859
rect 1494 887 1500 899
rect 1640 887 1646 899
rect 1494 859 1646 887
rect 1494 847 1500 859
rect 1640 847 1646 859
rect 1698 887 1704 899
rect 1844 887 1850 899
rect 1698 859 1850 887
rect 1698 847 1704 859
rect 1844 847 1850 859
rect 1902 887 1908 899
rect 2048 887 2054 899
rect 1902 859 2054 887
rect 1902 847 1908 859
rect 2048 847 2054 859
rect 2106 887 2112 899
rect 2252 887 2258 899
rect 2106 859 2258 887
rect 2106 847 2112 859
rect 2252 847 2258 859
rect 2310 887 2316 899
rect 2456 887 2462 899
rect 2310 859 2462 887
rect 2310 847 2316 859
rect 2456 847 2462 859
rect 2514 887 2520 899
rect 2660 887 2666 899
rect 2514 859 2666 887
rect 2514 847 2520 859
rect 2660 847 2666 859
rect 2718 887 2724 899
rect 2864 887 2870 899
rect 2718 859 2870 887
rect 2718 847 2724 859
rect 2864 847 2870 859
rect 2922 887 2928 899
rect 3068 887 3074 899
rect 2922 859 3074 887
rect 2922 847 2928 859
rect 3068 847 3074 859
rect 3126 887 3132 899
rect 3272 887 3278 899
rect 3126 859 3278 887
rect 3126 847 3132 859
rect 3272 847 3278 859
rect 3330 887 3336 899
rect 3476 887 3482 899
rect 3330 859 3482 887
rect 3330 847 3336 859
rect 3476 847 3482 859
rect 3534 887 3540 899
rect 3680 887 3686 899
rect 3534 859 3686 887
rect 3534 847 3540 859
rect 3680 847 3686 859
rect 3738 887 3744 899
rect 3884 887 3890 899
rect 3738 859 3890 887
rect 3738 847 3744 859
rect 3884 847 3890 859
rect 3942 887 3948 899
rect 4088 887 4094 899
rect 3942 859 4094 887
rect 3942 847 3948 859
rect 4088 847 4094 859
rect 4146 887 4152 899
rect 4292 887 4298 899
rect 4146 859 4298 887
rect 4146 847 4152 859
rect 4292 847 4298 859
rect 4350 887 4356 899
rect 4496 887 4502 899
rect 4350 859 4502 887
rect 4350 847 4356 859
rect 4496 847 4502 859
rect 4554 887 4560 899
rect 4700 887 4706 899
rect 4554 859 4706 887
rect 4554 847 4560 859
rect 4700 847 4706 859
rect 4758 887 4764 899
rect 4904 887 4910 899
rect 4758 859 4910 887
rect 4758 847 4764 859
rect 4904 847 4910 859
rect 4962 887 4968 899
rect 5108 887 5114 899
rect 4962 859 5114 887
rect 4962 847 4968 859
rect 5108 847 5114 859
rect 5166 887 5172 899
rect 5312 887 5318 899
rect 5166 859 5318 887
rect 5166 847 5172 859
rect 5312 847 5318 859
rect 5370 887 5376 899
rect 5516 887 5522 899
rect 5370 859 5522 887
rect 5370 847 5376 859
rect 5516 847 5522 859
rect 5574 887 5580 899
rect 5720 887 5726 899
rect 5574 859 5726 887
rect 5574 847 5580 859
rect 5720 847 5726 859
rect 5778 887 5784 899
rect 5924 887 5930 899
rect 5778 859 5930 887
rect 5778 847 5784 859
rect 5924 847 5930 859
rect 5982 887 5988 899
rect 6128 887 6134 899
rect 5982 859 6134 887
rect 5982 847 5988 859
rect 6128 847 6134 859
rect 6186 887 6192 899
rect 6332 887 6338 899
rect 6186 859 6338 887
rect 6186 847 6192 859
rect 6332 847 6338 859
rect 6390 887 6396 899
rect 6536 887 6542 899
rect 6390 859 6542 887
rect 6390 847 6396 859
rect 6536 847 6542 859
rect 6594 887 6600 899
rect 6740 887 6746 899
rect 6594 859 6746 887
rect 6594 847 6600 859
rect 6740 847 6746 859
rect 6798 887 6804 899
rect 6944 887 6950 899
rect 6798 859 6950 887
rect 6798 847 6804 859
rect 6944 847 6950 859
rect 7002 887 7008 899
rect 7148 887 7154 899
rect 7002 859 7154 887
rect 7002 847 7008 859
rect 7148 847 7154 859
rect 7206 887 7212 899
rect 7352 887 7358 899
rect 7206 859 7358 887
rect 7206 847 7212 859
rect 7352 847 7358 859
rect 7410 887 7416 899
rect 7556 887 7562 899
rect 7410 859 7562 887
rect 7410 847 7416 859
rect 7556 847 7562 859
rect 7614 887 7620 899
rect 7760 887 7766 899
rect 7614 859 7766 887
rect 7614 847 7620 859
rect 7760 847 7766 859
rect 7818 887 7824 899
rect 7964 887 7970 899
rect 7818 859 7970 887
rect 7818 847 7824 859
rect 7964 847 7970 859
rect 8022 887 8028 899
rect 8168 887 8174 899
rect 8022 859 8174 887
rect 8022 847 8028 859
rect 8168 847 8174 859
rect 8226 887 8232 899
rect 8372 887 8378 899
rect 8226 859 8378 887
rect 8226 847 8232 859
rect 8372 847 8378 859
rect 8430 887 8436 899
rect 8576 887 8582 899
rect 8430 859 8582 887
rect 8430 847 8436 859
rect 8576 847 8582 859
rect 8634 887 8640 899
rect 8780 887 8786 899
rect 8634 859 8786 887
rect 8634 847 8640 859
rect 8780 847 8786 859
rect 8838 887 8844 899
rect 8984 887 8990 899
rect 8838 859 8990 887
rect 8838 847 8844 859
rect 8984 847 8990 859
rect 9042 887 9048 899
rect 9188 887 9194 899
rect 9042 859 9194 887
rect 9042 847 9048 859
rect 9188 847 9194 859
rect 9246 887 9252 899
rect 9392 887 9398 899
rect 9246 859 9398 887
rect 9246 847 9252 859
rect 9392 847 9398 859
rect 9450 887 9456 899
rect 9596 887 9602 899
rect 9450 859 9602 887
rect 9450 847 9456 859
rect 9596 847 9602 859
rect 9654 887 9660 899
rect 9814 887 9820 899
rect 9654 859 9820 887
rect 9654 847 9660 859
rect 9814 847 9820 859
rect 9872 847 9878 899
rect 61 368 89 396
rect 12 -32 40 32
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_0
timestamp 1581321262
transform 1 0 9588 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1
timestamp 1581321262
transform 1 0 9384 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_2
timestamp 1581321262
transform 1 0 9180 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_3
timestamp 1581321262
transform 1 0 8976 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_4
timestamp 1581321262
transform 1 0 8772 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_5
timestamp 1581321262
transform 1 0 8568 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_6
timestamp 1581321262
transform 1 0 8364 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_7
timestamp 1581321262
transform 1 0 8160 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_8
timestamp 1581321262
transform 1 0 7956 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_9
timestamp 1581321262
transform 1 0 7752 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_10
timestamp 1581321262
transform 1 0 7548 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_11
timestamp 1581321262
transform 1 0 7344 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_12
timestamp 1581321262
transform 1 0 7140 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_13
timestamp 1581321262
transform 1 0 6936 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_14
timestamp 1581321262
transform 1 0 6732 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_15
timestamp 1581321262
transform 1 0 6528 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_16
timestamp 1581321262
transform 1 0 6324 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_17
timestamp 1581321262
transform 1 0 6120 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_18
timestamp 1581321262
transform 1 0 5916 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_19
timestamp 1581321262
transform 1 0 5712 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_20
timestamp 1581321262
transform 1 0 5508 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_21
timestamp 1581321262
transform 1 0 5304 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_22
timestamp 1581321262
transform 1 0 5100 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_23
timestamp 1581321262
transform 1 0 4896 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_24
timestamp 1581321262
transform 1 0 4692 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_25
timestamp 1581321262
transform 1 0 4488 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_26
timestamp 1581321262
transform 1 0 4284 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_27
timestamp 1581321262
transform 1 0 4080 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_28
timestamp 1581321262
transform 1 0 3876 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_29
timestamp 1581321262
transform 1 0 3672 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_30
timestamp 1581321262
transform 1 0 3468 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_31
timestamp 1581321262
transform 1 0 3264 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_32
timestamp 1581321262
transform 1 0 3060 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_33
timestamp 1581321262
transform 1 0 2856 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_34
timestamp 1581321262
transform 1 0 2652 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_35
timestamp 1581321262
transform 1 0 2448 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_36
timestamp 1581321262
transform 1 0 2244 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_37
timestamp 1581321262
transform 1 0 2040 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_38
timestamp 1581321262
transform 1 0 1836 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_39
timestamp 1581321262
transform 1 0 1632 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_40
timestamp 1581321262
transform 1 0 1428 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_41
timestamp 1581321262
transform 1 0 1224 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_42
timestamp 1581321262
transform 1 0 1020 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_43
timestamp 1581321262
transform 1 0 816 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_44
timestamp 1581321262
transform 1 0 612 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_45
timestamp 1581321262
transform 1 0 408 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_46
timestamp 1581321262
transform 1 0 204 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_47
timestamp 1581321262
transform 1 0 0 0 1 10065
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_48
timestamp 1581321262
transform 1 0 9588 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_49
timestamp 1581321262
transform 1 0 9384 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_50
timestamp 1581321262
transform 1 0 9180 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_51
timestamp 1581321262
transform 1 0 8976 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_52
timestamp 1581321262
transform 1 0 8568 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_53
timestamp 1581321262
transform 1 0 8364 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_54
timestamp 1581321262
transform 1 0 7548 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_55
timestamp 1581321262
transform 1 0 7344 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_56
timestamp 1581321262
transform 1 0 7140 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_57
timestamp 1581321262
transform 1 0 6936 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_58
timestamp 1581321262
transform 1 0 6528 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_59
timestamp 1581321262
transform 1 0 6324 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_60
timestamp 1581321262
transform 1 0 6120 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_61
timestamp 1581321262
transform 1 0 5916 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_62
timestamp 1581321262
transform 1 0 5712 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_63
timestamp 1581321262
transform 1 0 5508 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_64
timestamp 1581321262
transform 1 0 5304 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_65
timestamp 1581321262
transform 1 0 5100 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_66
timestamp 1581321262
transform 1 0 4896 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_67
timestamp 1581321262
transform 1 0 4692 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_68
timestamp 1581321262
transform 1 0 4080 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_69
timestamp 1581321262
transform 1 0 3876 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_70
timestamp 1581321262
transform 1 0 3264 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_71
timestamp 1581321262
transform 1 0 3060 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_72
timestamp 1581321262
transform 1 0 2652 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_73
timestamp 1581321262
transform 1 0 2448 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_74
timestamp 1581321262
transform 1 0 2040 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_75
timestamp 1581321262
transform 1 0 1632 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_76
timestamp 1581321262
transform 1 0 1428 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_77
timestamp 1581321262
transform 1 0 1224 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_78
timestamp 1581321262
transform 1 0 612 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_79
timestamp 1581321262
transform 1 0 408 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_80
timestamp 1581321262
transform 1 0 204 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_81
timestamp 1581321262
transform 1 0 8772 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_82
timestamp 1581321262
transform 1 0 8568 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_83
timestamp 1581321262
transform 1 0 7956 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_84
timestamp 1581321262
transform 1 0 7548 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_85
timestamp 1581321262
transform 1 0 7344 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_86
timestamp 1581321262
transform 1 0 7140 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_87
timestamp 1581321262
transform 1 0 6936 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_88
timestamp 1581321262
transform 1 0 6732 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_89
timestamp 1581321262
transform 1 0 6324 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_90
timestamp 1581321262
transform 1 0 6120 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_91
timestamp 1581321262
transform 1 0 5916 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_92
timestamp 1581321262
transform 1 0 5712 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_93
timestamp 1581321262
transform 1 0 5100 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_94
timestamp 1581321262
transform 1 0 4896 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_95
timestamp 1581321262
transform 1 0 4488 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_96
timestamp 1581321262
transform 1 0 3876 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_97
timestamp 1581321262
transform 1 0 3468 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_98
timestamp 1581321262
transform 1 0 3264 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_99
timestamp 1581321262
transform 1 0 2652 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_100
timestamp 1581321262
transform 1 0 2040 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_101
timestamp 1581321262
transform 1 0 1836 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_102
timestamp 1581321262
transform 1 0 1632 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_103
timestamp 1581321262
transform 1 0 1428 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_104
timestamp 1581321262
transform 1 0 816 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_105
timestamp 1581321262
transform 1 0 408 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_106
timestamp 1581321262
transform 1 0 204 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_107
timestamp 1581321262
transform 1 0 0 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_108
timestamp 1581321262
transform 1 0 9384 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_109
timestamp 1581321262
transform 1 0 8772 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_110
timestamp 1581321262
transform 1 0 8160 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_111
timestamp 1581321262
transform 1 0 7956 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_112
timestamp 1581321262
transform 1 0 7752 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_113
timestamp 1581321262
transform 1 0 6732 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_114
timestamp 1581321262
transform 1 0 5712 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_115
timestamp 1581321262
transform 1 0 5100 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_116
timestamp 1581321262
transform 1 0 4080 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_117
timestamp 1581321262
transform 1 0 3264 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_118
timestamp 1581321262
transform 1 0 2652 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_119
timestamp 1581321262
transform 1 0 2448 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_120
timestamp 1581321262
transform 1 0 1836 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_121
timestamp 1581321262
transform 1 0 1224 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_122
timestamp 1581321262
transform 1 0 612 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_123
timestamp 1581321262
transform 1 0 204 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_124
timestamp 1581321262
transform 1 0 9384 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_125
timestamp 1581321262
transform 1 0 9180 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_126
timestamp 1581321262
transform 1 0 8772 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_127
timestamp 1581321262
transform 1 0 8160 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_128
timestamp 1581321262
transform 1 0 7956 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_129
timestamp 1581321262
transform 1 0 7752 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_130
timestamp 1581321262
transform 1 0 7548 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_131
timestamp 1581321262
transform 1 0 6324 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_132
timestamp 1581321262
transform 1 0 6120 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_133
timestamp 1581321262
transform 1 0 5916 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_134
timestamp 1581321262
transform 1 0 5712 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_135
timestamp 1581321262
transform 1 0 5304 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_136
timestamp 1581321262
transform 1 0 4896 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_137
timestamp 1581321262
transform 1 0 4488 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_138
timestamp 1581321262
transform 1 0 3876 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_139
timestamp 1581321262
transform 1 0 3468 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_140
timestamp 1581321262
transform 1 0 2448 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_141
timestamp 1581321262
transform 1 0 1836 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_142
timestamp 1581321262
transform 1 0 1428 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_143
timestamp 1581321262
transform 1 0 1224 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_144
timestamp 1581321262
transform 1 0 816 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_145
timestamp 1581321262
transform 1 0 612 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_146
timestamp 1581321262
transform 1 0 408 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_147
timestamp 1581321262
transform 1 0 9384 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_148
timestamp 1581321262
transform 1 0 9180 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_149
timestamp 1581321262
transform 1 0 8976 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_150
timestamp 1581321262
transform 1 0 8772 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_151
timestamp 1581321262
transform 1 0 8568 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_152
timestamp 1581321262
transform 1 0 8364 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_153
timestamp 1581321262
transform 1 0 8160 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_154
timestamp 1581321262
transform 1 0 7752 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_155
timestamp 1581321262
transform 1 0 7548 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_156
timestamp 1581321262
transform 1 0 6732 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_157
timestamp 1581321262
transform 1 0 6528 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_158
timestamp 1581321262
transform 1 0 6120 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_159
timestamp 1581321262
transform 1 0 5916 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_160
timestamp 1581321262
transform 1 0 5508 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_161
timestamp 1581321262
transform 1 0 5304 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_162
timestamp 1581321262
transform 1 0 5100 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_163
timestamp 1581321262
transform 1 0 4896 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_164
timestamp 1581321262
transform 1 0 4284 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_165
timestamp 1581321262
transform 1 0 4080 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_166
timestamp 1581321262
transform 1 0 3672 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_167
timestamp 1581321262
transform 1 0 3264 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_168
timestamp 1581321262
transform 1 0 3060 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_169
timestamp 1581321262
transform 1 0 2448 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_170
timestamp 1581321262
transform 1 0 2040 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_171
timestamp 1581321262
transform 1 0 1428 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_172
timestamp 1581321262
transform 1 0 1224 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_173
timestamp 1581321262
transform 1 0 816 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_174
timestamp 1581321262
transform 1 0 612 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_175
timestamp 1581321262
transform 1 0 408 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_176
timestamp 1581321262
transform 1 0 9384 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_177
timestamp 1581321262
transform 1 0 8976 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_178
timestamp 1581321262
transform 1 0 8772 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_179
timestamp 1581321262
transform 1 0 8364 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_180
timestamp 1581321262
transform 1 0 8160 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_181
timestamp 1581321262
transform 1 0 7956 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_182
timestamp 1581321262
transform 1 0 7752 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_183
timestamp 1581321262
transform 1 0 7548 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_184
timestamp 1581321262
transform 1 0 7344 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_185
timestamp 1581321262
transform 1 0 6732 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_186
timestamp 1581321262
transform 1 0 6528 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_187
timestamp 1581321262
transform 1 0 5712 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_188
timestamp 1581321262
transform 1 0 4896 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_189
timestamp 1581321262
transform 1 0 4284 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_190
timestamp 1581321262
transform 1 0 3876 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_191
timestamp 1581321262
transform 1 0 3672 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_192
timestamp 1581321262
transform 1 0 2856 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_193
timestamp 1581321262
transform 1 0 2652 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_194
timestamp 1581321262
transform 1 0 2448 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_195
timestamp 1581321262
transform 1 0 1836 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_196
timestamp 1581321262
transform 1 0 1632 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_197
timestamp 1581321262
transform 1 0 1020 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_198
timestamp 1581321262
transform 1 0 816 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_199
timestamp 1581321262
transform 1 0 612 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_200
timestamp 1581321262
transform 1 0 204 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_201
timestamp 1581321262
transform 1 0 9180 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_202
timestamp 1581321262
transform 1 0 8976 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_203
timestamp 1581321262
transform 1 0 8568 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_204
timestamp 1581321262
transform 1 0 7752 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_205
timestamp 1581321262
transform 1 0 7548 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_206
timestamp 1581321262
transform 1 0 6936 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_207
timestamp 1581321262
transform 1 0 6732 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_208
timestamp 1581321262
transform 1 0 6120 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_209
timestamp 1581321262
transform 1 0 5916 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_210
timestamp 1581321262
transform 1 0 5712 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_211
timestamp 1581321262
transform 1 0 5100 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_212
timestamp 1581321262
transform 1 0 4896 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_213
timestamp 1581321262
transform 1 0 4080 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_214
timestamp 1581321262
transform 1 0 3876 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_215
timestamp 1581321262
transform 1 0 3264 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_216
timestamp 1581321262
transform 1 0 3060 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_217
timestamp 1581321262
transform 1 0 2856 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_218
timestamp 1581321262
transform 1 0 2652 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_219
timestamp 1581321262
transform 1 0 2448 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_220
timestamp 1581321262
transform 1 0 1632 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_221
timestamp 1581321262
transform 1 0 816 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_222
timestamp 1581321262
transform 1 0 408 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_223
timestamp 1581321262
transform 1 0 9384 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_224
timestamp 1581321262
transform 1 0 8364 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_225
timestamp 1581321262
transform 1 0 8160 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_226
timestamp 1581321262
transform 1 0 7752 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_227
timestamp 1581321262
transform 1 0 7140 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_228
timestamp 1581321262
transform 1 0 6936 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_229
timestamp 1581321262
transform 1 0 6732 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_230
timestamp 1581321262
transform 1 0 6324 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_231
timestamp 1581321262
transform 1 0 6120 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_232
timestamp 1581321262
transform 1 0 5100 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_233
timestamp 1581321262
transform 1 0 4896 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_234
timestamp 1581321262
transform 1 0 4692 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_235
timestamp 1581321262
transform 1 0 3264 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_236
timestamp 1581321262
transform 1 0 3060 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_237
timestamp 1581321262
transform 1 0 2856 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_238
timestamp 1581321262
transform 1 0 2652 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_239
timestamp 1581321262
transform 1 0 2244 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_240
timestamp 1581321262
transform 1 0 2040 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_241
timestamp 1581321262
transform 1 0 1836 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_242
timestamp 1581321262
transform 1 0 1632 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_243
timestamp 1581321262
transform 1 0 1428 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_244
timestamp 1581321262
transform 1 0 1224 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_245
timestamp 1581321262
transform 1 0 204 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_246
timestamp 1581321262
transform 1 0 8364 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_247
timestamp 1581321262
transform 1 0 7752 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_248
timestamp 1581321262
transform 1 0 7548 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_249
timestamp 1581321262
transform 1 0 7344 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_250
timestamp 1581321262
transform 1 0 5916 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_251
timestamp 1581321262
transform 1 0 5712 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_252
timestamp 1581321262
transform 1 0 4692 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_253
timestamp 1581321262
transform 1 0 4488 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_254
timestamp 1581321262
transform 1 0 4080 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_255
timestamp 1581321262
transform 1 0 3876 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_256
timestamp 1581321262
transform 1 0 3468 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_257
timestamp 1581321262
transform 1 0 3264 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_258
timestamp 1581321262
transform 1 0 3060 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_259
timestamp 1581321262
transform 1 0 2448 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_260
timestamp 1581321262
transform 1 0 2244 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_261
timestamp 1581321262
transform 1 0 1632 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_262
timestamp 1581321262
transform 1 0 1428 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_263
timestamp 1581321262
transform 1 0 1224 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_264
timestamp 1581321262
transform 1 0 1020 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_265
timestamp 1581321262
transform 1 0 612 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_266
timestamp 1581321262
transform 1 0 9588 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_267
timestamp 1581321262
transform 1 0 8976 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_268
timestamp 1581321262
transform 1 0 8772 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_269
timestamp 1581321262
transform 1 0 8364 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_270
timestamp 1581321262
transform 1 0 8160 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_271
timestamp 1581321262
transform 1 0 7956 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_272
timestamp 1581321262
transform 1 0 7140 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_273
timestamp 1581321262
transform 1 0 6936 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_274
timestamp 1581321262
transform 1 0 6528 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_275
timestamp 1581321262
transform 1 0 6120 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_276
timestamp 1581321262
transform 1 0 4896 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_277
timestamp 1581321262
transform 1 0 4488 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_278
timestamp 1581321262
transform 1 0 4284 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_279
timestamp 1581321262
transform 1 0 4080 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_280
timestamp 1581321262
transform 1 0 3468 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_281
timestamp 1581321262
transform 1 0 2856 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_282
timestamp 1581321262
transform 1 0 2448 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_283
timestamp 1581321262
transform 1 0 2244 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_284
timestamp 1581321262
transform 1 0 1836 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_285
timestamp 1581321262
transform 1 0 816 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_286
timestamp 1581321262
transform 1 0 204 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_287
timestamp 1581321262
transform 1 0 9180 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_288
timestamp 1581321262
transform 1 0 8772 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_289
timestamp 1581321262
transform 1 0 7956 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_290
timestamp 1581321262
transform 1 0 7548 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_291
timestamp 1581321262
transform 1 0 7140 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_292
timestamp 1581321262
transform 1 0 6528 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_293
timestamp 1581321262
transform 1 0 6324 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_294
timestamp 1581321262
transform 1 0 5916 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_295
timestamp 1581321262
transform 1 0 5712 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_296
timestamp 1581321262
transform 1 0 4896 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_297
timestamp 1581321262
transform 1 0 4284 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_298
timestamp 1581321262
transform 1 0 3060 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_299
timestamp 1581321262
transform 1 0 2040 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_300
timestamp 1581321262
transform 1 0 1836 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_301
timestamp 1581321262
transform 1 0 1632 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_302
timestamp 1581321262
transform 1 0 1224 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_303
timestamp 1581321262
transform 1 0 408 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_304
timestamp 1581321262
transform 1 0 9180 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_305
timestamp 1581321262
transform 1 0 8976 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_306
timestamp 1581321262
transform 1 0 8364 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_307
timestamp 1581321262
transform 1 0 8160 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_308
timestamp 1581321262
transform 1 0 7752 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_309
timestamp 1581321262
transform 1 0 7344 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_310
timestamp 1581321262
transform 1 0 6732 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_311
timestamp 1581321262
transform 1 0 6324 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_312
timestamp 1581321262
transform 1 0 4896 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_313
timestamp 1581321262
transform 1 0 3876 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_314
timestamp 1581321262
transform 1 0 3672 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_315
timestamp 1581321262
transform 1 0 3468 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_316
timestamp 1581321262
transform 1 0 3264 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_317
timestamp 1581321262
transform 1 0 3060 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_318
timestamp 1581321262
transform 1 0 2244 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_319
timestamp 1581321262
transform 1 0 1836 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_320
timestamp 1581321262
transform 1 0 1632 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_321
timestamp 1581321262
transform 1 0 1020 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_322
timestamp 1581321262
transform 1 0 612 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_323
timestamp 1581321262
transform 1 0 408 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_324
timestamp 1581321262
transform 1 0 0 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_325
timestamp 1581321262
transform 1 0 9588 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_326
timestamp 1581321262
transform 1 0 9180 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_327
timestamp 1581321262
transform 1 0 8772 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_328
timestamp 1581321262
transform 1 0 8568 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_329
timestamp 1581321262
transform 1 0 7752 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_330
timestamp 1581321262
transform 1 0 7140 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_331
timestamp 1581321262
transform 1 0 6936 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_332
timestamp 1581321262
transform 1 0 6120 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_333
timestamp 1581321262
transform 1 0 5100 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_334
timestamp 1581321262
transform 1 0 4896 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_335
timestamp 1581321262
transform 1 0 4488 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_336
timestamp 1581321262
transform 1 0 4284 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_337
timestamp 1581321262
transform 1 0 2856 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_338
timestamp 1581321262
transform 1 0 2040 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_339
timestamp 1581321262
transform 1 0 1836 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_340
timestamp 1581321262
transform 1 0 1632 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_341
timestamp 1581321262
transform 1 0 1020 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_342
timestamp 1581321262
transform 1 0 816 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_343
timestamp 1581321262
transform 1 0 612 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_344
timestamp 1581321262
transform 1 0 408 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_345
timestamp 1581321262
transform 1 0 204 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_346
timestamp 1581321262
transform 1 0 9180 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_347
timestamp 1581321262
transform 1 0 8568 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_348
timestamp 1581321262
transform 1 0 8364 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_349
timestamp 1581321262
transform 1 0 7752 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_350
timestamp 1581321262
transform 1 0 7344 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_351
timestamp 1581321262
transform 1 0 6936 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_352
timestamp 1581321262
transform 1 0 6528 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_353
timestamp 1581321262
transform 1 0 6324 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_354
timestamp 1581321262
transform 1 0 5916 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_355
timestamp 1581321262
transform 1 0 5712 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_356
timestamp 1581321262
transform 1 0 5508 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_357
timestamp 1581321262
transform 1 0 4692 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_358
timestamp 1581321262
transform 1 0 4488 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_359
timestamp 1581321262
transform 1 0 4080 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_360
timestamp 1581321262
transform 1 0 3876 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_361
timestamp 1581321262
transform 1 0 3672 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_362
timestamp 1581321262
transform 1 0 3468 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_363
timestamp 1581321262
transform 1 0 2652 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_364
timestamp 1581321262
transform 1 0 1020 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_365
timestamp 1581321262
transform 1 0 612 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_366
timestamp 1581321262
transform 1 0 408 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_367
timestamp 1581321262
transform 1 0 204 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_368
timestamp 1581321262
transform 1 0 0 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_369
timestamp 1581321262
transform 1 0 9588 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_370
timestamp 1581321262
transform 1 0 9180 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_371
timestamp 1581321262
transform 1 0 8976 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_372
timestamp 1581321262
transform 1 0 8772 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_373
timestamp 1581321262
transform 1 0 7752 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_374
timestamp 1581321262
transform 1 0 7548 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_375
timestamp 1581321262
transform 1 0 6936 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_376
timestamp 1581321262
transform 1 0 6120 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_377
timestamp 1581321262
transform 1 0 5916 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_378
timestamp 1581321262
transform 1 0 4896 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_379
timestamp 1581321262
transform 1 0 4080 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_380
timestamp 1581321262
transform 1 0 3468 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_381
timestamp 1581321262
transform 1 0 2652 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_382
timestamp 1581321262
transform 1 0 2448 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_383
timestamp 1581321262
transform 1 0 1632 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_384
timestamp 1581321262
transform 1 0 1428 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_385
timestamp 1581321262
transform 1 0 1224 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_386
timestamp 1581321262
transform 1 0 1020 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_387
timestamp 1581321262
transform 1 0 612 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_388
timestamp 1581321262
transform 1 0 204 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_389
timestamp 1581321262
transform 1 0 0 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_390
timestamp 1581321262
transform 1 0 9588 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_391
timestamp 1581321262
transform 1 0 9384 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_392
timestamp 1581321262
transform 1 0 8976 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_393
timestamp 1581321262
transform 1 0 8568 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_394
timestamp 1581321262
transform 1 0 8364 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_395
timestamp 1581321262
transform 1 0 8160 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_396
timestamp 1581321262
transform 1 0 7752 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_397
timestamp 1581321262
transform 1 0 7140 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_398
timestamp 1581321262
transform 1 0 6732 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_399
timestamp 1581321262
transform 1 0 6528 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_400
timestamp 1581321262
transform 1 0 6120 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_401
timestamp 1581321262
transform 1 0 5508 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_402
timestamp 1581321262
transform 1 0 5304 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_403
timestamp 1581321262
transform 1 0 5100 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_404
timestamp 1581321262
transform 1 0 4080 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_405
timestamp 1581321262
transform 1 0 3672 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_406
timestamp 1581321262
transform 1 0 3264 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_407
timestamp 1581321262
transform 1 0 2652 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_408
timestamp 1581321262
transform 1 0 1836 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_409
timestamp 1581321262
transform 1 0 1632 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_410
timestamp 1581321262
transform 1 0 1428 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_411
timestamp 1581321262
transform 1 0 408 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_412
timestamp 1581321262
transform 1 0 0 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_413
timestamp 1581321262
transform 1 0 9180 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_414
timestamp 1581321262
transform 1 0 8976 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_415
timestamp 1581321262
transform 1 0 8772 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_416
timestamp 1581321262
transform 1 0 8568 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_417
timestamp 1581321262
transform 1 0 8364 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_418
timestamp 1581321262
transform 1 0 7752 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_419
timestamp 1581321262
transform 1 0 7344 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_420
timestamp 1581321262
transform 1 0 6732 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_421
timestamp 1581321262
transform 1 0 6528 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_422
timestamp 1581321262
transform 1 0 6120 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_423
timestamp 1581321262
transform 1 0 5712 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_424
timestamp 1581321262
transform 1 0 5100 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_425
timestamp 1581321262
transform 1 0 4896 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_426
timestamp 1581321262
transform 1 0 4692 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_427
timestamp 1581321262
transform 1 0 4488 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_428
timestamp 1581321262
transform 1 0 3672 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_429
timestamp 1581321262
transform 1 0 2856 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_430
timestamp 1581321262
transform 1 0 2448 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_431
timestamp 1581321262
transform 1 0 1020 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_432
timestamp 1581321262
transform 1 0 408 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_433
timestamp 1581321262
transform 1 0 204 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_434
timestamp 1581321262
transform 1 0 8976 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_435
timestamp 1581321262
transform 1 0 8568 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_436
timestamp 1581321262
transform 1 0 8160 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_437
timestamp 1581321262
transform 1 0 7752 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_438
timestamp 1581321262
transform 1 0 7344 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_439
timestamp 1581321262
transform 1 0 6936 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_440
timestamp 1581321262
transform 1 0 6528 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_441
timestamp 1581321262
transform 1 0 5916 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_442
timestamp 1581321262
transform 1 0 5712 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_443
timestamp 1581321262
transform 1 0 4488 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_444
timestamp 1581321262
transform 1 0 4284 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_445
timestamp 1581321262
transform 1 0 4080 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_446
timestamp 1581321262
transform 1 0 3876 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_447
timestamp 1581321262
transform 1 0 3468 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_448
timestamp 1581321262
transform 1 0 3060 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_449
timestamp 1581321262
transform 1 0 2244 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_450
timestamp 1581321262
transform 1 0 2040 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_451
timestamp 1581321262
transform 1 0 1632 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_452
timestamp 1581321262
transform 1 0 1428 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_453
timestamp 1581321262
transform 1 0 1224 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_454
timestamp 1581321262
transform 1 0 1020 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_455
timestamp 1581321262
transform 1 0 816 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_456
timestamp 1581321262
transform 1 0 612 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_457
timestamp 1581321262
transform 1 0 9588 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_458
timestamp 1581321262
transform 1 0 8976 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_459
timestamp 1581321262
transform 1 0 7956 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_460
timestamp 1581321262
transform 1 0 7548 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_461
timestamp 1581321262
transform 1 0 7344 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_462
timestamp 1581321262
transform 1 0 7140 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_463
timestamp 1581321262
transform 1 0 6936 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_464
timestamp 1581321262
transform 1 0 6732 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_465
timestamp 1581321262
transform 1 0 6324 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_466
timestamp 1581321262
transform 1 0 6120 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_467
timestamp 1581321262
transform 1 0 5508 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_468
timestamp 1581321262
transform 1 0 4896 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_469
timestamp 1581321262
transform 1 0 4692 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_470
timestamp 1581321262
transform 1 0 4488 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_471
timestamp 1581321262
transform 1 0 4284 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_472
timestamp 1581321262
transform 1 0 3876 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_473
timestamp 1581321262
transform 1 0 3468 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_474
timestamp 1581321262
transform 1 0 3060 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_475
timestamp 1581321262
transform 1 0 2856 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_476
timestamp 1581321262
transform 1 0 2448 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_477
timestamp 1581321262
transform 1 0 2040 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_478
timestamp 1581321262
transform 1 0 1224 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_479
timestamp 1581321262
transform 1 0 816 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_480
timestamp 1581321262
transform 1 0 612 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_481
timestamp 1581321262
transform 1 0 9180 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_482
timestamp 1581321262
transform 1 0 8568 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_483
timestamp 1581321262
transform 1 0 8364 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_484
timestamp 1581321262
transform 1 0 7752 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_485
timestamp 1581321262
transform 1 0 7548 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_486
timestamp 1581321262
transform 1 0 7344 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_487
timestamp 1581321262
transform 1 0 6936 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_488
timestamp 1581321262
transform 1 0 6732 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_489
timestamp 1581321262
transform 1 0 6528 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_490
timestamp 1581321262
transform 1 0 6324 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_491
timestamp 1581321262
transform 1 0 4692 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_492
timestamp 1581321262
transform 1 0 4488 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_493
timestamp 1581321262
transform 1 0 3672 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_494
timestamp 1581321262
transform 1 0 3468 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_495
timestamp 1581321262
transform 1 0 3060 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_496
timestamp 1581321262
transform 1 0 2856 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_497
timestamp 1581321262
transform 1 0 2448 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_498
timestamp 1581321262
transform 1 0 1428 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_499
timestamp 1581321262
transform 1 0 1224 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_500
timestamp 1581321262
transform 1 0 1020 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_501
timestamp 1581321262
transform 1 0 9588 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_502
timestamp 1581321262
transform 1 0 9384 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_503
timestamp 1581321262
transform 1 0 9180 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_504
timestamp 1581321262
transform 1 0 8772 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_505
timestamp 1581321262
transform 1 0 8568 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_506
timestamp 1581321262
transform 1 0 8364 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_507
timestamp 1581321262
transform 1 0 8160 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_508
timestamp 1581321262
transform 1 0 7956 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_509
timestamp 1581321262
transform 1 0 6936 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_510
timestamp 1581321262
transform 1 0 6324 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_511
timestamp 1581321262
transform 1 0 6120 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_512
timestamp 1581321262
transform 1 0 5508 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_513
timestamp 1581321262
transform 1 0 5304 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_514
timestamp 1581321262
transform 1 0 5100 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_515
timestamp 1581321262
transform 1 0 4488 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_516
timestamp 1581321262
transform 1 0 4284 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_517
timestamp 1581321262
transform 1 0 4080 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_518
timestamp 1581321262
transform 1 0 3876 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_519
timestamp 1581321262
transform 1 0 3264 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_520
timestamp 1581321262
transform 1 0 2856 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_521
timestamp 1581321262
transform 1 0 2448 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_522
timestamp 1581321262
transform 1 0 1428 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_523
timestamp 1581321262
transform 1 0 1224 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_524
timestamp 1581321262
transform 1 0 9588 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_525
timestamp 1581321262
transform 1 0 9384 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_526
timestamp 1581321262
transform 1 0 8568 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_527
timestamp 1581321262
transform 1 0 7752 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_528
timestamp 1581321262
transform 1 0 7344 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_529
timestamp 1581321262
transform 1 0 6936 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_530
timestamp 1581321262
transform 1 0 6528 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_531
timestamp 1581321262
transform 1 0 5712 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_532
timestamp 1581321262
transform 1 0 5508 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_533
timestamp 1581321262
transform 1 0 4896 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_534
timestamp 1581321262
transform 1 0 4488 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_535
timestamp 1581321262
transform 1 0 3876 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_536
timestamp 1581321262
transform 1 0 3672 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_537
timestamp 1581321262
transform 1 0 3468 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_538
timestamp 1581321262
transform 1 0 3060 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_539
timestamp 1581321262
transform 1 0 2244 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_540
timestamp 1581321262
transform 1 0 1428 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_541
timestamp 1581321262
transform 1 0 816 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_542
timestamp 1581321262
transform 1 0 9588 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_543
timestamp 1581321262
transform 1 0 9384 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_544
timestamp 1581321262
transform 1 0 9180 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_545
timestamp 1581321262
transform 1 0 8976 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_546
timestamp 1581321262
transform 1 0 8772 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_547
timestamp 1581321262
transform 1 0 8568 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_548
timestamp 1581321262
transform 1 0 8364 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_549
timestamp 1581321262
transform 1 0 8160 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_550
timestamp 1581321262
transform 1 0 6732 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_551
timestamp 1581321262
transform 1 0 6324 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_552
timestamp 1581321262
transform 1 0 6120 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_553
timestamp 1581321262
transform 1 0 5916 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_554
timestamp 1581321262
transform 1 0 5508 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_555
timestamp 1581321262
transform 1 0 5100 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_556
timestamp 1581321262
transform 1 0 4896 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_557
timestamp 1581321262
transform 1 0 4692 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_558
timestamp 1581321262
transform 1 0 4488 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_559
timestamp 1581321262
transform 1 0 4284 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_560
timestamp 1581321262
transform 1 0 3672 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_561
timestamp 1581321262
transform 1 0 3264 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_562
timestamp 1581321262
transform 1 0 2448 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_563
timestamp 1581321262
transform 1 0 2244 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_564
timestamp 1581321262
transform 1 0 2040 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_565
timestamp 1581321262
transform 1 0 816 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_566
timestamp 1581321262
transform 1 0 408 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_567
timestamp 1581321262
transform 1 0 204 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_568
timestamp 1581321262
transform 1 0 9384 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_569
timestamp 1581321262
transform 1 0 9180 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_570
timestamp 1581321262
transform 1 0 8772 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_571
timestamp 1581321262
transform 1 0 8160 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_572
timestamp 1581321262
transform 1 0 7344 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_573
timestamp 1581321262
transform 1 0 6732 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_574
timestamp 1581321262
transform 1 0 6528 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_575
timestamp 1581321262
transform 1 0 5916 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_576
timestamp 1581321262
transform 1 0 5712 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_577
timestamp 1581321262
transform 1 0 5508 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_578
timestamp 1581321262
transform 1 0 5304 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_579
timestamp 1581321262
transform 1 0 5100 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_580
timestamp 1581321262
transform 1 0 4488 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_581
timestamp 1581321262
transform 1 0 4284 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_582
timestamp 1581321262
transform 1 0 4080 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_583
timestamp 1581321262
transform 1 0 3876 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_584
timestamp 1581321262
transform 1 0 3672 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_585
timestamp 1581321262
transform 1 0 3468 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_586
timestamp 1581321262
transform 1 0 3264 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_587
timestamp 1581321262
transform 1 0 3060 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_588
timestamp 1581321262
transform 1 0 2652 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_589
timestamp 1581321262
transform 1 0 2448 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_590
timestamp 1581321262
transform 1 0 2040 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_591
timestamp 1581321262
transform 1 0 1836 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_592
timestamp 1581321262
transform 1 0 1428 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_593
timestamp 1581321262
transform 1 0 1224 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_594
timestamp 1581321262
transform 1 0 1020 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_595
timestamp 1581321262
transform 1 0 816 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_596
timestamp 1581321262
transform 1 0 408 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_597
timestamp 1581321262
transform 1 0 0 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_598
timestamp 1581321262
transform 1 0 9384 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_599
timestamp 1581321262
transform 1 0 9180 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_600
timestamp 1581321262
transform 1 0 8772 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_601
timestamp 1581321262
transform 1 0 7956 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_602
timestamp 1581321262
transform 1 0 7752 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_603
timestamp 1581321262
transform 1 0 7344 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_604
timestamp 1581321262
transform 1 0 6120 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_605
timestamp 1581321262
transform 1 0 5916 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_606
timestamp 1581321262
transform 1 0 5508 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_607
timestamp 1581321262
transform 1 0 5304 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_608
timestamp 1581321262
transform 1 0 4692 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_609
timestamp 1581321262
transform 1 0 4080 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_610
timestamp 1581321262
transform 1 0 3672 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_611
timestamp 1581321262
transform 1 0 3468 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_612
timestamp 1581321262
transform 1 0 3060 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_613
timestamp 1581321262
transform 1 0 2040 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_614
timestamp 1581321262
transform 1 0 1632 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_615
timestamp 1581321262
transform 1 0 1428 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_616
timestamp 1581321262
transform 1 0 612 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_617
timestamp 1581321262
transform 1 0 204 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_618
timestamp 1581321262
transform 1 0 0 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_619
timestamp 1581321262
transform 1 0 9588 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_620
timestamp 1581321262
transform 1 0 8772 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_621
timestamp 1581321262
transform 1 0 8568 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_622
timestamp 1581321262
transform 1 0 7956 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_623
timestamp 1581321262
transform 1 0 7344 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_624
timestamp 1581321262
transform 1 0 7140 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_625
timestamp 1581321262
transform 1 0 6936 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_626
timestamp 1581321262
transform 1 0 6732 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_627
timestamp 1581321262
transform 1 0 6528 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_628
timestamp 1581321262
transform 1 0 6120 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_629
timestamp 1581321262
transform 1 0 5712 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_630
timestamp 1581321262
transform 1 0 4488 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_631
timestamp 1581321262
transform 1 0 2856 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_632
timestamp 1581321262
transform 1 0 2448 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_633
timestamp 1581321262
transform 1 0 2040 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_634
timestamp 1581321262
transform 1 0 1836 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_635
timestamp 1581321262
transform 1 0 1632 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_636
timestamp 1581321262
transform 1 0 816 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_637
timestamp 1581321262
transform 1 0 408 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_638
timestamp 1581321262
transform 1 0 0 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_639
timestamp 1581321262
transform 1 0 9384 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_640
timestamp 1581321262
transform 1 0 8976 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_641
timestamp 1581321262
transform 1 0 7956 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_642
timestamp 1581321262
transform 1 0 7752 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_643
timestamp 1581321262
transform 1 0 7548 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_644
timestamp 1581321262
transform 1 0 7344 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_645
timestamp 1581321262
transform 1 0 7140 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_646
timestamp 1581321262
transform 1 0 6936 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_647
timestamp 1581321262
transform 1 0 6732 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_648
timestamp 1581321262
transform 1 0 6324 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_649
timestamp 1581321262
transform 1 0 5916 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_650
timestamp 1581321262
transform 1 0 5712 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_651
timestamp 1581321262
transform 1 0 5508 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_652
timestamp 1581321262
transform 1 0 5304 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_653
timestamp 1581321262
transform 1 0 5100 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_654
timestamp 1581321262
transform 1 0 4896 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_655
timestamp 1581321262
transform 1 0 4284 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_656
timestamp 1581321262
transform 1 0 3876 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_657
timestamp 1581321262
transform 1 0 3264 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_658
timestamp 1581321262
transform 1 0 2856 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_659
timestamp 1581321262
transform 1 0 2448 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_660
timestamp 1581321262
transform 1 0 2040 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_661
timestamp 1581321262
transform 1 0 1428 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_662
timestamp 1581321262
transform 1 0 1224 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_663
timestamp 1581321262
transform 1 0 816 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_664
timestamp 1581321262
transform 1 0 408 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_665
timestamp 1581321262
transform 1 0 0 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_666
timestamp 1581321262
transform 1 0 8772 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_667
timestamp 1581321262
transform 1 0 7956 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_668
timestamp 1581321262
transform 1 0 7548 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_669
timestamp 1581321262
transform 1 0 7140 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_670
timestamp 1581321262
transform 1 0 6732 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_671
timestamp 1581321262
transform 1 0 6528 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_672
timestamp 1581321262
transform 1 0 6324 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_673
timestamp 1581321262
transform 1 0 6120 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_674
timestamp 1581321262
transform 1 0 5508 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_675
timestamp 1581321262
transform 1 0 5304 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_676
timestamp 1581321262
transform 1 0 5100 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_677
timestamp 1581321262
transform 1 0 3672 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_678
timestamp 1581321262
transform 1 0 3468 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_679
timestamp 1581321262
transform 1 0 3264 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_680
timestamp 1581321262
transform 1 0 2856 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_681
timestamp 1581321262
transform 1 0 2448 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_682
timestamp 1581321262
transform 1 0 2244 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_683
timestamp 1581321262
transform 1 0 1020 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_684
timestamp 1581321262
transform 1 0 612 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_685
timestamp 1581321262
transform 1 0 204 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_686
timestamp 1581321262
transform 1 0 9588 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_687
timestamp 1581321262
transform 1 0 9384 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_688
timestamp 1581321262
transform 1 0 8976 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_689
timestamp 1581321262
transform 1 0 8364 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_690
timestamp 1581321262
transform 1 0 7956 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_691
timestamp 1581321262
transform 1 0 7752 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_692
timestamp 1581321262
transform 1 0 7548 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_693
timestamp 1581321262
transform 1 0 7344 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_694
timestamp 1581321262
transform 1 0 6528 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_695
timestamp 1581321262
transform 1 0 6324 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_696
timestamp 1581321262
transform 1 0 5916 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_697
timestamp 1581321262
transform 1 0 5712 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_698
timestamp 1581321262
transform 1 0 5508 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_699
timestamp 1581321262
transform 1 0 5100 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_700
timestamp 1581321262
transform 1 0 4896 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_701
timestamp 1581321262
transform 1 0 4488 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_702
timestamp 1581321262
transform 1 0 4284 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_703
timestamp 1581321262
transform 1 0 3468 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_704
timestamp 1581321262
transform 1 0 3264 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_705
timestamp 1581321262
transform 1 0 2856 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_706
timestamp 1581321262
transform 1 0 2652 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_707
timestamp 1581321262
transform 1 0 1632 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_708
timestamp 1581321262
transform 1 0 1428 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_709
timestamp 1581321262
transform 1 0 1224 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_710
timestamp 1581321262
transform 1 0 0 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_711
timestamp 1581321262
transform 1 0 9180 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_712
timestamp 1581321262
transform 1 0 8772 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_713
timestamp 1581321262
transform 1 0 8364 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_714
timestamp 1581321262
transform 1 0 8160 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_715
timestamp 1581321262
transform 1 0 7752 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_716
timestamp 1581321262
transform 1 0 5712 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_717
timestamp 1581321262
transform 1 0 5508 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_718
timestamp 1581321262
transform 1 0 5100 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_719
timestamp 1581321262
transform 1 0 4896 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_720
timestamp 1581321262
transform 1 0 4488 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_721
timestamp 1581321262
transform 1 0 4284 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_722
timestamp 1581321262
transform 1 0 3672 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_723
timestamp 1581321262
transform 1 0 3468 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_724
timestamp 1581321262
transform 1 0 3264 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_725
timestamp 1581321262
transform 1 0 3060 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_726
timestamp 1581321262
transform 1 0 2652 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_727
timestamp 1581321262
transform 1 0 2448 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_728
timestamp 1581321262
transform 1 0 2040 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_729
timestamp 1581321262
transform 1 0 1632 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_730
timestamp 1581321262
transform 1 0 204 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_731
timestamp 1581321262
transform 1 0 9180 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_732
timestamp 1581321262
transform 1 0 8976 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_733
timestamp 1581321262
transform 1 0 8772 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_734
timestamp 1581321262
transform 1 0 8364 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_735
timestamp 1581321262
transform 1 0 8160 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_736
timestamp 1581321262
transform 1 0 7548 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_737
timestamp 1581321262
transform 1 0 6936 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_738
timestamp 1581321262
transform 1 0 6324 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_739
timestamp 1581321262
transform 1 0 5508 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_740
timestamp 1581321262
transform 1 0 5304 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_741
timestamp 1581321262
transform 1 0 5100 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_742
timestamp 1581321262
transform 1 0 4896 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_743
timestamp 1581321262
transform 1 0 4692 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_744
timestamp 1581321262
transform 1 0 4488 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_745
timestamp 1581321262
transform 1 0 4284 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_746
timestamp 1581321262
transform 1 0 4080 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_747
timestamp 1581321262
transform 1 0 3876 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_748
timestamp 1581321262
transform 1 0 3468 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_749
timestamp 1581321262
transform 1 0 3264 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_750
timestamp 1581321262
transform 1 0 2652 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_751
timestamp 1581321262
transform 1 0 2448 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_752
timestamp 1581321262
transform 1 0 1428 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_753
timestamp 1581321262
transform 1 0 1224 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_754
timestamp 1581321262
transform 1 0 1020 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_755
timestamp 1581321262
transform 1 0 816 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_756
timestamp 1581321262
transform 1 0 612 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_757
timestamp 1581321262
transform 1 0 204 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_758
timestamp 1581321262
transform 1 0 9588 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_759
timestamp 1581321262
transform 1 0 9180 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_760
timestamp 1581321262
transform 1 0 8976 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_761
timestamp 1581321262
transform 1 0 8568 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_762
timestamp 1581321262
transform 1 0 8160 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_763
timestamp 1581321262
transform 1 0 7752 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_764
timestamp 1581321262
transform 1 0 7344 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_765
timestamp 1581321262
transform 1 0 7140 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_766
timestamp 1581321262
transform 1 0 6936 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_767
timestamp 1581321262
transform 1 0 6732 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_768
timestamp 1581321262
transform 1 0 6324 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_769
timestamp 1581321262
transform 1 0 5712 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_770
timestamp 1581321262
transform 1 0 5304 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_771
timestamp 1581321262
transform 1 0 4896 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_772
timestamp 1581321262
transform 1 0 4488 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_773
timestamp 1581321262
transform 1 0 4284 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_774
timestamp 1581321262
transform 1 0 3468 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_775
timestamp 1581321262
transform 1 0 2040 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_776
timestamp 1581321262
transform 1 0 1632 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_777
timestamp 1581321262
transform 1 0 1428 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_778
timestamp 1581321262
transform 1 0 1020 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_779
timestamp 1581321262
transform 1 0 816 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_780
timestamp 1581321262
transform 1 0 612 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_781
timestamp 1581321262
transform 1 0 408 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_782
timestamp 1581321262
transform 1 0 204 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_783
timestamp 1581321262
transform 1 0 0 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_784
timestamp 1581321262
transform 1 0 9588 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_785
timestamp 1581321262
transform 1 0 8976 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_786
timestamp 1581321262
transform 1 0 8568 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_787
timestamp 1581321262
transform 1 0 8364 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_788
timestamp 1581321262
transform 1 0 8160 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_789
timestamp 1581321262
transform 1 0 7956 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_790
timestamp 1581321262
transform 1 0 7548 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_791
timestamp 1581321262
transform 1 0 7344 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_792
timestamp 1581321262
transform 1 0 6936 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_793
timestamp 1581321262
transform 1 0 6732 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_794
timestamp 1581321262
transform 1 0 6528 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_795
timestamp 1581321262
transform 1 0 6120 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_796
timestamp 1581321262
transform 1 0 5712 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_797
timestamp 1581321262
transform 1 0 5508 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_798
timestamp 1581321262
transform 1 0 5304 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_799
timestamp 1581321262
transform 1 0 5100 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_800
timestamp 1581321262
transform 1 0 4896 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_801
timestamp 1581321262
transform 1 0 4488 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_802
timestamp 1581321262
transform 1 0 4284 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_803
timestamp 1581321262
transform 1 0 4080 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_804
timestamp 1581321262
transform 1 0 3876 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_805
timestamp 1581321262
transform 1 0 3468 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_806
timestamp 1581321262
transform 1 0 2652 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_807
timestamp 1581321262
transform 1 0 2040 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_808
timestamp 1581321262
transform 1 0 1836 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_809
timestamp 1581321262
transform 1 0 1224 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_810
timestamp 1581321262
transform 1 0 204 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_811
timestamp 1581321262
transform 1 0 0 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_812
timestamp 1581321262
transform 1 0 8976 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_813
timestamp 1581321262
transform 1 0 8568 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_814
timestamp 1581321262
transform 1 0 8364 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_815
timestamp 1581321262
transform 1 0 8160 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_816
timestamp 1581321262
transform 1 0 7956 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_817
timestamp 1581321262
transform 1 0 7752 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_818
timestamp 1581321262
transform 1 0 7344 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_819
timestamp 1581321262
transform 1 0 7140 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_820
timestamp 1581321262
transform 1 0 6936 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_821
timestamp 1581321262
transform 1 0 6732 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_822
timestamp 1581321262
transform 1 0 6324 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_823
timestamp 1581321262
transform 1 0 6120 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_824
timestamp 1581321262
transform 1 0 5916 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_825
timestamp 1581321262
transform 1 0 5712 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_826
timestamp 1581321262
transform 1 0 5304 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_827
timestamp 1581321262
transform 1 0 4896 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_828
timestamp 1581321262
transform 1 0 4488 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_829
timestamp 1581321262
transform 1 0 3672 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_830
timestamp 1581321262
transform 1 0 3264 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_831
timestamp 1581321262
transform 1 0 2652 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_832
timestamp 1581321262
transform 1 0 2040 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_833
timestamp 1581321262
transform 1 0 1836 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_834
timestamp 1581321262
transform 1 0 1224 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_835
timestamp 1581321262
transform 1 0 816 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_836
timestamp 1581321262
transform 1 0 612 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_837
timestamp 1581321262
transform 1 0 408 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_838
timestamp 1581321262
transform 1 0 9588 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_839
timestamp 1581321262
transform 1 0 8976 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_840
timestamp 1581321262
transform 1 0 8568 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_841
timestamp 1581321262
transform 1 0 8160 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_842
timestamp 1581321262
transform 1 0 7956 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_843
timestamp 1581321262
transform 1 0 7548 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_844
timestamp 1581321262
transform 1 0 7344 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_845
timestamp 1581321262
transform 1 0 6732 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_846
timestamp 1581321262
transform 1 0 6120 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_847
timestamp 1581321262
transform 1 0 5916 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_848
timestamp 1581321262
transform 1 0 5304 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_849
timestamp 1581321262
transform 1 0 4896 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_850
timestamp 1581321262
transform 1 0 4692 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_851
timestamp 1581321262
transform 1 0 4488 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_852
timestamp 1581321262
transform 1 0 4284 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_853
timestamp 1581321262
transform 1 0 3468 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_854
timestamp 1581321262
transform 1 0 3264 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_855
timestamp 1581321262
transform 1 0 3060 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_856
timestamp 1581321262
transform 1 0 2856 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_857
timestamp 1581321262
transform 1 0 2244 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_858
timestamp 1581321262
transform 1 0 2040 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_859
timestamp 1581321262
transform 1 0 1632 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_860
timestamp 1581321262
transform 1 0 1020 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_861
timestamp 1581321262
transform 1 0 816 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_862
timestamp 1581321262
transform 1 0 0 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_863
timestamp 1581321262
transform 1 0 9588 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_864
timestamp 1581321262
transform 1 0 9384 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_865
timestamp 1581321262
transform 1 0 9180 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_866
timestamp 1581321262
transform 1 0 8568 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_867
timestamp 1581321262
transform 1 0 7140 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_868
timestamp 1581321262
transform 1 0 6528 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_869
timestamp 1581321262
transform 1 0 4896 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_870
timestamp 1581321262
transform 1 0 4488 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_871
timestamp 1581321262
transform 1 0 3876 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_872
timestamp 1581321262
transform 1 0 3672 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_873
timestamp 1581321262
transform 1 0 3468 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_874
timestamp 1581321262
transform 1 0 2652 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_875
timestamp 1581321262
transform 1 0 2040 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_876
timestamp 1581321262
transform 1 0 1836 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_877
timestamp 1581321262
transform 1 0 1632 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_878
timestamp 1581321262
transform 1 0 816 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_879
timestamp 1581321262
transform 1 0 9384 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_880
timestamp 1581321262
transform 1 0 9180 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_881
timestamp 1581321262
transform 1 0 8772 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_882
timestamp 1581321262
transform 1 0 8160 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_883
timestamp 1581321262
transform 1 0 7956 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_884
timestamp 1581321262
transform 1 0 7752 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_885
timestamp 1581321262
transform 1 0 7140 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_886
timestamp 1581321262
transform 1 0 6732 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_887
timestamp 1581321262
transform 1 0 5508 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_888
timestamp 1581321262
transform 1 0 5304 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_889
timestamp 1581321262
transform 1 0 4896 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_890
timestamp 1581321262
transform 1 0 4080 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_891
timestamp 1581321262
transform 1 0 3672 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_892
timestamp 1581321262
transform 1 0 3060 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_893
timestamp 1581321262
transform 1 0 2856 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_894
timestamp 1581321262
transform 1 0 2652 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_895
timestamp 1581321262
transform 1 0 2448 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_896
timestamp 1581321262
transform 1 0 2040 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_897
timestamp 1581321262
transform 1 0 1836 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_898
timestamp 1581321262
transform 1 0 1632 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_899
timestamp 1581321262
transform 1 0 816 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_900
timestamp 1581321262
transform 1 0 612 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_901
timestamp 1581321262
transform 1 0 408 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_902
timestamp 1581321262
transform 1 0 204 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_903
timestamp 1581321262
transform 1 0 9180 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_904
timestamp 1581321262
transform 1 0 8568 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_905
timestamp 1581321262
transform 1 0 8364 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_906
timestamp 1581321262
transform 1 0 8160 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_907
timestamp 1581321262
transform 1 0 7956 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_908
timestamp 1581321262
transform 1 0 7752 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_909
timestamp 1581321262
transform 1 0 7344 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_910
timestamp 1581321262
transform 1 0 7140 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_911
timestamp 1581321262
transform 1 0 6732 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_912
timestamp 1581321262
transform 1 0 6324 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_913
timestamp 1581321262
transform 1 0 6120 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_914
timestamp 1581321262
transform 1 0 5100 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_915
timestamp 1581321262
transform 1 0 4692 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_916
timestamp 1581321262
transform 1 0 4080 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_917
timestamp 1581321262
transform 1 0 3876 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_918
timestamp 1581321262
transform 1 0 3672 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_919
timestamp 1581321262
transform 1 0 2856 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_920
timestamp 1581321262
transform 1 0 1836 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_921
timestamp 1581321262
transform 1 0 1632 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_922
timestamp 1581321262
transform 1 0 408 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_923
timestamp 1581321262
transform 1 0 204 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_924
timestamp 1581321262
transform 1 0 0 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_925
timestamp 1581321262
transform 1 0 9588 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_926
timestamp 1581321262
transform 1 0 9384 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_927
timestamp 1581321262
transform 1 0 9180 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_928
timestamp 1581321262
transform 1 0 8568 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_929
timestamp 1581321262
transform 1 0 7344 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_930
timestamp 1581321262
transform 1 0 7140 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_931
timestamp 1581321262
transform 1 0 6936 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_932
timestamp 1581321262
transform 1 0 6732 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_933
timestamp 1581321262
transform 1 0 6528 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_934
timestamp 1581321262
transform 1 0 6324 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_935
timestamp 1581321262
transform 1 0 5916 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_936
timestamp 1581321262
transform 1 0 5712 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_937
timestamp 1581321262
transform 1 0 5508 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_938
timestamp 1581321262
transform 1 0 5304 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_939
timestamp 1581321262
transform 1 0 5100 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_940
timestamp 1581321262
transform 1 0 4692 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_941
timestamp 1581321262
transform 1 0 4488 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_942
timestamp 1581321262
transform 1 0 3672 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_943
timestamp 1581321262
transform 1 0 2652 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_944
timestamp 1581321262
transform 1 0 2244 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_945
timestamp 1581321262
transform 1 0 2040 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_946
timestamp 1581321262
transform 1 0 816 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_947
timestamp 1581321262
transform 1 0 612 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_948
timestamp 1581321262
transform 1 0 0 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_949
timestamp 1581321262
transform 1 0 9384 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_950
timestamp 1581321262
transform 1 0 9180 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_951
timestamp 1581321262
transform 1 0 8976 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_952
timestamp 1581321262
transform 1 0 8364 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_953
timestamp 1581321262
transform 1 0 8160 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_954
timestamp 1581321262
transform 1 0 7956 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_955
timestamp 1581321262
transform 1 0 7140 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_956
timestamp 1581321262
transform 1 0 6732 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_957
timestamp 1581321262
transform 1 0 6324 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_958
timestamp 1581321262
transform 1 0 6120 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_959
timestamp 1581321262
transform 1 0 5916 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_960
timestamp 1581321262
transform 1 0 5100 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_961
timestamp 1581321262
transform 1 0 4896 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_962
timestamp 1581321262
transform 1 0 4692 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_963
timestamp 1581321262
transform 1 0 4488 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_964
timestamp 1581321262
transform 1 0 4284 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_965
timestamp 1581321262
transform 1 0 3876 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_966
timestamp 1581321262
transform 1 0 2856 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_967
timestamp 1581321262
transform 1 0 2652 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_968
timestamp 1581321262
transform 1 0 2448 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_969
timestamp 1581321262
transform 1 0 2244 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_970
timestamp 1581321262
transform 1 0 2040 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_971
timestamp 1581321262
transform 1 0 1632 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_972
timestamp 1581321262
transform 1 0 1224 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_973
timestamp 1581321262
transform 1 0 816 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_974
timestamp 1581321262
transform 1 0 612 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_975
timestamp 1581321262
transform 1 0 204 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_976
timestamp 1581321262
transform 1 0 0 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_977
timestamp 1581321262
transform 1 0 9588 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_978
timestamp 1581321262
transform 1 0 9180 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_979
timestamp 1581321262
transform 1 0 8976 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_980
timestamp 1581321262
transform 1 0 8364 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_981
timestamp 1581321262
transform 1 0 7752 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_982
timestamp 1581321262
transform 1 0 6732 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_983
timestamp 1581321262
transform 1 0 5916 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_984
timestamp 1581321262
transform 1 0 5712 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_985
timestamp 1581321262
transform 1 0 5304 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_986
timestamp 1581321262
transform 1 0 5100 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_987
timestamp 1581321262
transform 1 0 4896 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_988
timestamp 1581321262
transform 1 0 4692 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_989
timestamp 1581321262
transform 1 0 4488 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_990
timestamp 1581321262
transform 1 0 4080 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_991
timestamp 1581321262
transform 1 0 3264 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_992
timestamp 1581321262
transform 1 0 3060 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_993
timestamp 1581321262
transform 1 0 2856 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_994
timestamp 1581321262
transform 1 0 2244 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_995
timestamp 1581321262
transform 1 0 2040 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_996
timestamp 1581321262
transform 1 0 1632 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_997
timestamp 1581321262
transform 1 0 1428 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_998
timestamp 1581321262
transform 1 0 1020 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_999
timestamp 1581321262
transform 1 0 612 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1000
timestamp 1581321262
transform 1 0 408 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1001
timestamp 1581321262
transform 1 0 204 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1002
timestamp 1581321262
transform 1 0 9588 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1003
timestamp 1581321262
transform 1 0 8976 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1004
timestamp 1581321262
transform 1 0 8568 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1005
timestamp 1581321262
transform 1 0 8364 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1006
timestamp 1581321262
transform 1 0 7548 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1007
timestamp 1581321262
transform 1 0 7344 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1008
timestamp 1581321262
transform 1 0 7140 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1009
timestamp 1581321262
transform 1 0 6936 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1010
timestamp 1581321262
transform 1 0 6528 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1011
timestamp 1581321262
transform 1 0 5100 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1012
timestamp 1581321262
transform 1 0 4896 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1013
timestamp 1581321262
transform 1 0 4692 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1014
timestamp 1581321262
transform 1 0 4488 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1015
timestamp 1581321262
transform 1 0 3876 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1016
timestamp 1581321262
transform 1 0 3672 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1017
timestamp 1581321262
transform 1 0 3264 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1018
timestamp 1581321262
transform 1 0 2652 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1019
timestamp 1581321262
transform 1 0 2244 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1020
timestamp 1581321262
transform 1 0 1632 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1021
timestamp 1581321262
transform 1 0 1428 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1022
timestamp 1581321262
transform 1 0 1020 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_one_cell  sky130_rom_krom_rom_base_one_cell_1023
timestamp 1581321262
transform 1 0 612 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_0
timestamp 1581321262
transform 1 0 8772 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1
timestamp 1581321262
transform 1 0 8160 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_2
timestamp 1581321262
transform 1 0 7956 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_3
timestamp 1581321262
transform 1 0 7752 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_4
timestamp 1581321262
transform 1 0 6732 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_5
timestamp 1581321262
transform 1 0 4488 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_6
timestamp 1581321262
transform 1 0 4284 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_7
timestamp 1581321262
transform 1 0 3672 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_8
timestamp 1581321262
transform 1 0 3468 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_9
timestamp 1581321262
transform 1 0 2856 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_10
timestamp 1581321262
transform 1 0 2244 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_11
timestamp 1581321262
transform 1 0 1836 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_12
timestamp 1581321262
transform 1 0 1020 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_13
timestamp 1581321262
transform 1 0 816 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_14
timestamp 1581321262
transform 1 0 0 0 1 9861
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_15
timestamp 1581321262
transform 1 0 9588 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_16
timestamp 1581321262
transform 1 0 9384 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_17
timestamp 1581321262
transform 1 0 9180 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_18
timestamp 1581321262
transform 1 0 8976 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_19
timestamp 1581321262
transform 1 0 8364 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_20
timestamp 1581321262
transform 1 0 8160 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_21
timestamp 1581321262
transform 1 0 7752 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_22
timestamp 1581321262
transform 1 0 6528 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_23
timestamp 1581321262
transform 1 0 5508 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_24
timestamp 1581321262
transform 1 0 5304 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_25
timestamp 1581321262
transform 1 0 4692 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_26
timestamp 1581321262
transform 1 0 4284 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_27
timestamp 1581321262
transform 1 0 4080 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_28
timestamp 1581321262
transform 1 0 3672 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_29
timestamp 1581321262
transform 1 0 3060 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_30
timestamp 1581321262
transform 1 0 2856 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_31
timestamp 1581321262
transform 1 0 2448 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_32
timestamp 1581321262
transform 1 0 2244 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_33
timestamp 1581321262
transform 1 0 1224 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_34
timestamp 1581321262
transform 1 0 1020 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_35
timestamp 1581321262
transform 1 0 612 0 1 9657
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_36
timestamp 1581321262
transform 1 0 9588 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_37
timestamp 1581321262
transform 1 0 9180 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_38
timestamp 1581321262
transform 1 0 8976 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_39
timestamp 1581321262
transform 1 0 8568 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_40
timestamp 1581321262
transform 1 0 8364 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_41
timestamp 1581321262
transform 1 0 7548 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_42
timestamp 1581321262
transform 1 0 7344 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_43
timestamp 1581321262
transform 1 0 7140 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_44
timestamp 1581321262
transform 1 0 6936 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_45
timestamp 1581321262
transform 1 0 6528 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_46
timestamp 1581321262
transform 1 0 6324 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_47
timestamp 1581321262
transform 1 0 6120 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_48
timestamp 1581321262
transform 1 0 5916 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_49
timestamp 1581321262
transform 1 0 5508 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_50
timestamp 1581321262
transform 1 0 5304 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_51
timestamp 1581321262
transform 1 0 4896 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_52
timestamp 1581321262
transform 1 0 4692 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_53
timestamp 1581321262
transform 1 0 4488 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_54
timestamp 1581321262
transform 1 0 4284 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_55
timestamp 1581321262
transform 1 0 3876 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_56
timestamp 1581321262
transform 1 0 3672 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_57
timestamp 1581321262
transform 1 0 3468 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_58
timestamp 1581321262
transform 1 0 3060 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_59
timestamp 1581321262
transform 1 0 2856 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_60
timestamp 1581321262
transform 1 0 2244 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_61
timestamp 1581321262
transform 1 0 2040 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_62
timestamp 1581321262
transform 1 0 1632 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_63
timestamp 1581321262
transform 1 0 1428 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_64
timestamp 1581321262
transform 1 0 1020 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_65
timestamp 1581321262
transform 1 0 816 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_66
timestamp 1581321262
transform 1 0 408 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_67
timestamp 1581321262
transform 1 0 0 0 1 9349
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_68
timestamp 1581321262
transform 1 0 9588 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_69
timestamp 1581321262
transform 1 0 8976 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_70
timestamp 1581321262
transform 1 0 8568 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_71
timestamp 1581321262
transform 1 0 8364 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_72
timestamp 1581321262
transform 1 0 7344 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_73
timestamp 1581321262
transform 1 0 7140 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_74
timestamp 1581321262
transform 1 0 6936 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_75
timestamp 1581321262
transform 1 0 6732 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_76
timestamp 1581321262
transform 1 0 6528 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_77
timestamp 1581321262
transform 1 0 5508 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_78
timestamp 1581321262
transform 1 0 5100 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_79
timestamp 1581321262
transform 1 0 4692 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_80
timestamp 1581321262
transform 1 0 4284 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_81
timestamp 1581321262
transform 1 0 4080 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_82
timestamp 1581321262
transform 1 0 3672 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_83
timestamp 1581321262
transform 1 0 3264 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_84
timestamp 1581321262
transform 1 0 3060 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_85
timestamp 1581321262
transform 1 0 2856 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_86
timestamp 1581321262
transform 1 0 2652 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_87
timestamp 1581321262
transform 1 0 2244 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_88
timestamp 1581321262
transform 1 0 2040 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_89
timestamp 1581321262
transform 1 0 1632 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_90
timestamp 1581321262
transform 1 0 1020 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_91
timestamp 1581321262
transform 1 0 204 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_92
timestamp 1581321262
transform 1 0 0 0 1 9145
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_93
timestamp 1581321262
transform 1 0 9588 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_94
timestamp 1581321262
transform 1 0 7956 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_95
timestamp 1581321262
transform 1 0 7344 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_96
timestamp 1581321262
transform 1 0 7140 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_97
timestamp 1581321262
transform 1 0 6936 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_98
timestamp 1581321262
transform 1 0 6324 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_99
timestamp 1581321262
transform 1 0 5712 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_100
timestamp 1581321262
transform 1 0 4692 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_101
timestamp 1581321262
transform 1 0 4488 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_102
timestamp 1581321262
transform 1 0 3876 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_103
timestamp 1581321262
transform 1 0 3468 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_104
timestamp 1581321262
transform 1 0 2856 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_105
timestamp 1581321262
transform 1 0 2652 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_106
timestamp 1581321262
transform 1 0 2244 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_107
timestamp 1581321262
transform 1 0 1836 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_108
timestamp 1581321262
transform 1 0 1632 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_109
timestamp 1581321262
transform 1 0 1020 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_110
timestamp 1581321262
transform 1 0 204 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_111
timestamp 1581321262
transform 1 0 0 0 1 8941
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_112
timestamp 1581321262
transform 1 0 9588 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_113
timestamp 1581321262
transform 1 0 9180 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_114
timestamp 1581321262
transform 1 0 8568 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_115
timestamp 1581321262
transform 1 0 7140 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_116
timestamp 1581321262
transform 1 0 6936 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_117
timestamp 1581321262
transform 1 0 6324 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_118
timestamp 1581321262
transform 1 0 6120 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_119
timestamp 1581321262
transform 1 0 5916 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_120
timestamp 1581321262
transform 1 0 5508 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_121
timestamp 1581321262
transform 1 0 5304 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_122
timestamp 1581321262
transform 1 0 5100 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_123
timestamp 1581321262
transform 1 0 4692 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_124
timestamp 1581321262
transform 1 0 4488 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_125
timestamp 1581321262
transform 1 0 4080 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_126
timestamp 1581321262
transform 1 0 3468 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_127
timestamp 1581321262
transform 1 0 3264 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_128
timestamp 1581321262
transform 1 0 3060 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_129
timestamp 1581321262
transform 1 0 2244 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_130
timestamp 1581321262
transform 1 0 2040 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_131
timestamp 1581321262
transform 1 0 1428 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_132
timestamp 1581321262
transform 1 0 1224 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_133
timestamp 1581321262
transform 1 0 408 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_134
timestamp 1581321262
transform 1 0 0 0 1 8737
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_135
timestamp 1581321262
transform 1 0 9588 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_136
timestamp 1581321262
transform 1 0 9384 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_137
timestamp 1581321262
transform 1 0 8772 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_138
timestamp 1581321262
transform 1 0 8364 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_139
timestamp 1581321262
transform 1 0 8160 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_140
timestamp 1581321262
transform 1 0 7956 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_141
timestamp 1581321262
transform 1 0 7344 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_142
timestamp 1581321262
transform 1 0 7140 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_143
timestamp 1581321262
transform 1 0 6528 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_144
timestamp 1581321262
transform 1 0 6324 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_145
timestamp 1581321262
transform 1 0 5508 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_146
timestamp 1581321262
transform 1 0 5304 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_147
timestamp 1581321262
transform 1 0 4692 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_148
timestamp 1581321262
transform 1 0 4488 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_149
timestamp 1581321262
transform 1 0 4284 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_150
timestamp 1581321262
transform 1 0 3672 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_151
timestamp 1581321262
transform 1 0 3468 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_152
timestamp 1581321262
transform 1 0 2244 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_153
timestamp 1581321262
transform 1 0 2040 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_154
timestamp 1581321262
transform 1 0 1836 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_155
timestamp 1581321262
transform 1 0 1428 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_156
timestamp 1581321262
transform 1 0 1224 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_157
timestamp 1581321262
transform 1 0 1020 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_158
timestamp 1581321262
transform 1 0 612 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_159
timestamp 1581321262
transform 1 0 204 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_160
timestamp 1581321262
transform 1 0 0 0 1 8533
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_161
timestamp 1581321262
transform 1 0 9588 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_162
timestamp 1581321262
transform 1 0 9180 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_163
timestamp 1581321262
transform 1 0 8976 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_164
timestamp 1581321262
transform 1 0 8772 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_165
timestamp 1581321262
transform 1 0 8568 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_166
timestamp 1581321262
transform 1 0 7956 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_167
timestamp 1581321262
transform 1 0 7548 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_168
timestamp 1581321262
transform 1 0 7344 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_169
timestamp 1581321262
transform 1 0 6528 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_170
timestamp 1581321262
transform 1 0 5916 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_171
timestamp 1581321262
transform 1 0 5712 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_172
timestamp 1581321262
transform 1 0 5508 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_173
timestamp 1581321262
transform 1 0 5304 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_174
timestamp 1581321262
transform 1 0 4488 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_175
timestamp 1581321262
transform 1 0 4284 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_176
timestamp 1581321262
transform 1 0 4080 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_177
timestamp 1581321262
transform 1 0 3876 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_178
timestamp 1581321262
transform 1 0 3672 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_179
timestamp 1581321262
transform 1 0 3468 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_180
timestamp 1581321262
transform 1 0 2448 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_181
timestamp 1581321262
transform 1 0 1020 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_182
timestamp 1581321262
transform 1 0 816 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_183
timestamp 1581321262
transform 1 0 612 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_184
timestamp 1581321262
transform 1 0 408 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_185
timestamp 1581321262
transform 1 0 0 0 1 8329
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_186
timestamp 1581321262
transform 1 0 9588 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_187
timestamp 1581321262
transform 1 0 9384 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_188
timestamp 1581321262
transform 1 0 9180 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_189
timestamp 1581321262
transform 1 0 8976 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_190
timestamp 1581321262
transform 1 0 8772 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_191
timestamp 1581321262
transform 1 0 8568 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_192
timestamp 1581321262
transform 1 0 8160 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_193
timestamp 1581321262
transform 1 0 7956 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_194
timestamp 1581321262
transform 1 0 7140 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_195
timestamp 1581321262
transform 1 0 6936 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_196
timestamp 1581321262
transform 1 0 6732 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_197
timestamp 1581321262
transform 1 0 6528 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_198
timestamp 1581321262
transform 1 0 6324 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_199
timestamp 1581321262
transform 1 0 6120 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_200
timestamp 1581321262
transform 1 0 5508 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_201
timestamp 1581321262
transform 1 0 5304 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_202
timestamp 1581321262
transform 1 0 5100 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_203
timestamp 1581321262
transform 1 0 4896 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_204
timestamp 1581321262
transform 1 0 4284 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_205
timestamp 1581321262
transform 1 0 3672 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_206
timestamp 1581321262
transform 1 0 2856 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_207
timestamp 1581321262
transform 1 0 2652 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_208
timestamp 1581321262
transform 1 0 2040 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_209
timestamp 1581321262
transform 1 0 1836 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_210
timestamp 1581321262
transform 1 0 816 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_211
timestamp 1581321262
transform 1 0 408 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_212
timestamp 1581321262
transform 1 0 204 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_213
timestamp 1581321262
transform 1 0 0 0 1 8125
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_214
timestamp 1581321262
transform 1 0 9384 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_215
timestamp 1581321262
transform 1 0 9180 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_216
timestamp 1581321262
transform 1 0 8568 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_217
timestamp 1581321262
transform 1 0 7752 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_218
timestamp 1581321262
transform 1 0 7548 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_219
timestamp 1581321262
transform 1 0 7344 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_220
timestamp 1581321262
transform 1 0 6732 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_221
timestamp 1581321262
transform 1 0 6324 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_222
timestamp 1581321262
transform 1 0 5916 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_223
timestamp 1581321262
transform 1 0 5712 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_224
timestamp 1581321262
transform 1 0 5508 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_225
timestamp 1581321262
transform 1 0 5304 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_226
timestamp 1581321262
transform 1 0 5100 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_227
timestamp 1581321262
transform 1 0 4692 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_228
timestamp 1581321262
transform 1 0 3876 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_229
timestamp 1581321262
transform 1 0 3672 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_230
timestamp 1581321262
transform 1 0 3264 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_231
timestamp 1581321262
transform 1 0 3060 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_232
timestamp 1581321262
transform 1 0 2652 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_233
timestamp 1581321262
transform 1 0 2040 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_234
timestamp 1581321262
transform 1 0 1632 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_235
timestamp 1581321262
transform 1 0 1428 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_236
timestamp 1581321262
transform 1 0 1224 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_237
timestamp 1581321262
transform 1 0 1020 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_238
timestamp 1581321262
transform 1 0 612 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_239
timestamp 1581321262
transform 1 0 408 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_240
timestamp 1581321262
transform 1 0 0 0 1 7921
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_241
timestamp 1581321262
transform 1 0 9588 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_242
timestamp 1581321262
transform 1 0 9384 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_243
timestamp 1581321262
transform 1 0 8976 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_244
timestamp 1581321262
transform 1 0 8568 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_245
timestamp 1581321262
transform 1 0 8364 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_246
timestamp 1581321262
transform 1 0 8160 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_247
timestamp 1581321262
transform 1 0 7752 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_248
timestamp 1581321262
transform 1 0 7344 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_249
timestamp 1581321262
transform 1 0 6936 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_250
timestamp 1581321262
transform 1 0 6732 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_251
timestamp 1581321262
transform 1 0 6120 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_252
timestamp 1581321262
transform 1 0 5508 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_253
timestamp 1581321262
transform 1 0 5304 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_254
timestamp 1581321262
transform 1 0 5100 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_255
timestamp 1581321262
transform 1 0 4692 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_256
timestamp 1581321262
transform 1 0 4488 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_257
timestamp 1581321262
transform 1 0 4080 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_258
timestamp 1581321262
transform 1 0 3876 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_259
timestamp 1581321262
transform 1 0 3672 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_260
timestamp 1581321262
transform 1 0 3468 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_261
timestamp 1581321262
transform 1 0 3264 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_262
timestamp 1581321262
transform 1 0 2856 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_263
timestamp 1581321262
transform 1 0 2652 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_264
timestamp 1581321262
transform 1 0 2448 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_265
timestamp 1581321262
transform 1 0 2244 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_266
timestamp 1581321262
transform 1 0 1428 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_267
timestamp 1581321262
transform 1 0 1020 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_268
timestamp 1581321262
transform 1 0 816 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_269
timestamp 1581321262
transform 1 0 612 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_270
timestamp 1581321262
transform 1 0 204 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_271
timestamp 1581321262
transform 1 0 0 0 1 7613
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_272
timestamp 1581321262
transform 1 0 9588 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_273
timestamp 1581321262
transform 1 0 9384 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_274
timestamp 1581321262
transform 1 0 8772 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_275
timestamp 1581321262
transform 1 0 8568 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_276
timestamp 1581321262
transform 1 0 7956 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_277
timestamp 1581321262
transform 1 0 7548 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_278
timestamp 1581321262
transform 1 0 7140 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_279
timestamp 1581321262
transform 1 0 6936 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_280
timestamp 1581321262
transform 1 0 6528 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_281
timestamp 1581321262
transform 1 0 6120 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_282
timestamp 1581321262
transform 1 0 5916 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_283
timestamp 1581321262
transform 1 0 5712 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_284
timestamp 1581321262
transform 1 0 5508 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_285
timestamp 1581321262
transform 1 0 5304 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_286
timestamp 1581321262
transform 1 0 5100 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_287
timestamp 1581321262
transform 1 0 4692 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_288
timestamp 1581321262
transform 1 0 4488 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_289
timestamp 1581321262
transform 1 0 4284 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_290
timestamp 1581321262
transform 1 0 4080 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_291
timestamp 1581321262
transform 1 0 2856 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_292
timestamp 1581321262
transform 1 0 2652 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_293
timestamp 1581321262
transform 1 0 2448 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_294
timestamp 1581321262
transform 1 0 2040 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_295
timestamp 1581321262
transform 1 0 1428 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_296
timestamp 1581321262
transform 1 0 1224 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_297
timestamp 1581321262
transform 1 0 816 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_298
timestamp 1581321262
transform 1 0 204 0 1 7409
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_299
timestamp 1581321262
transform 1 0 9384 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_300
timestamp 1581321262
transform 1 0 8976 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_301
timestamp 1581321262
transform 1 0 8364 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_302
timestamp 1581321262
transform 1 0 8160 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_303
timestamp 1581321262
transform 1 0 7956 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_304
timestamp 1581321262
transform 1 0 7548 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_305
timestamp 1581321262
transform 1 0 7344 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_306
timestamp 1581321262
transform 1 0 6732 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_307
timestamp 1581321262
transform 1 0 6528 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_308
timestamp 1581321262
transform 1 0 6324 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_309
timestamp 1581321262
transform 1 0 5916 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_310
timestamp 1581321262
transform 1 0 5712 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_311
timestamp 1581321262
transform 1 0 5508 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_312
timestamp 1581321262
transform 1 0 5304 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_313
timestamp 1581321262
transform 1 0 4692 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_314
timestamp 1581321262
transform 1 0 4080 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_315
timestamp 1581321262
transform 1 0 3876 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_316
timestamp 1581321262
transform 1 0 3672 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_317
timestamp 1581321262
transform 1 0 3468 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_318
timestamp 1581321262
transform 1 0 3264 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_319
timestamp 1581321262
transform 1 0 3060 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_320
timestamp 1581321262
transform 1 0 2652 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_321
timestamp 1581321262
transform 1 0 2448 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_322
timestamp 1581321262
transform 1 0 2244 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_323
timestamp 1581321262
transform 1 0 1428 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_324
timestamp 1581321262
transform 1 0 1224 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_325
timestamp 1581321262
transform 1 0 0 0 1 7205
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_326
timestamp 1581321262
transform 1 0 9588 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_327
timestamp 1581321262
transform 1 0 9384 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_328
timestamp 1581321262
transform 1 0 8976 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_329
timestamp 1581321262
transform 1 0 8772 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_330
timestamp 1581321262
transform 1 0 8160 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_331
timestamp 1581321262
transform 1 0 7956 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_332
timestamp 1581321262
transform 1 0 7548 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_333
timestamp 1581321262
transform 1 0 7140 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_334
timestamp 1581321262
transform 1 0 6732 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_335
timestamp 1581321262
transform 1 0 6120 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_336
timestamp 1581321262
transform 1 0 5304 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_337
timestamp 1581321262
transform 1 0 5100 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_338
timestamp 1581321262
transform 1 0 4896 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_339
timestamp 1581321262
transform 1 0 4284 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_340
timestamp 1581321262
transform 1 0 3264 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_341
timestamp 1581321262
transform 1 0 3060 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_342
timestamp 1581321262
transform 1 0 2856 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_343
timestamp 1581321262
transform 1 0 2448 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_344
timestamp 1581321262
transform 1 0 2244 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_345
timestamp 1581321262
transform 1 0 2040 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_346
timestamp 1581321262
transform 1 0 1836 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_347
timestamp 1581321262
transform 1 0 1632 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_348
timestamp 1581321262
transform 1 0 1428 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_349
timestamp 1581321262
transform 1 0 1224 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_350
timestamp 1581321262
transform 1 0 816 0 1 7001
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_351
timestamp 1581321262
transform 1 0 9384 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_352
timestamp 1581321262
transform 1 0 8568 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_353
timestamp 1581321262
transform 1 0 8364 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_354
timestamp 1581321262
transform 1 0 8160 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_355
timestamp 1581321262
transform 1 0 7956 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_356
timestamp 1581321262
transform 1 0 7344 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_357
timestamp 1581321262
transform 1 0 7140 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_358
timestamp 1581321262
transform 1 0 6732 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_359
timestamp 1581321262
transform 1 0 6528 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_360
timestamp 1581321262
transform 1 0 6324 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_361
timestamp 1581321262
transform 1 0 5712 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_362
timestamp 1581321262
transform 1 0 5508 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_363
timestamp 1581321262
transform 1 0 5304 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_364
timestamp 1581321262
transform 1 0 5100 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_365
timestamp 1581321262
transform 1 0 4692 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_366
timestamp 1581321262
transform 1 0 4488 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_367
timestamp 1581321262
transform 1 0 4284 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_368
timestamp 1581321262
transform 1 0 3876 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_369
timestamp 1581321262
transform 1 0 3672 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_370
timestamp 1581321262
transform 1 0 3264 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_371
timestamp 1581321262
transform 1 0 3060 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_372
timestamp 1581321262
transform 1 0 2856 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_373
timestamp 1581321262
transform 1 0 2244 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_374
timestamp 1581321262
transform 1 0 2040 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_375
timestamp 1581321262
transform 1 0 1836 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_376
timestamp 1581321262
transform 1 0 816 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_377
timestamp 1581321262
transform 1 0 408 0 1 6797
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_378
timestamp 1581321262
transform 1 0 9180 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_379
timestamp 1581321262
transform 1 0 8772 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_380
timestamp 1581321262
transform 1 0 7956 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_381
timestamp 1581321262
transform 1 0 7548 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_382
timestamp 1581321262
transform 1 0 7344 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_383
timestamp 1581321262
transform 1 0 6936 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_384
timestamp 1581321262
transform 1 0 6324 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_385
timestamp 1581321262
transform 1 0 5916 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_386
timestamp 1581321262
transform 1 0 5712 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_387
timestamp 1581321262
transform 1 0 4896 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_388
timestamp 1581321262
transform 1 0 4692 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_389
timestamp 1581321262
transform 1 0 4488 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_390
timestamp 1581321262
transform 1 0 4284 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_391
timestamp 1581321262
transform 1 0 3876 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_392
timestamp 1581321262
transform 1 0 3468 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_393
timestamp 1581321262
transform 1 0 3060 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_394
timestamp 1581321262
transform 1 0 2856 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_395
timestamp 1581321262
transform 1 0 2448 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_396
timestamp 1581321262
transform 1 0 2244 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_397
timestamp 1581321262
transform 1 0 2040 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_398
timestamp 1581321262
transform 1 0 1224 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_399
timestamp 1581321262
transform 1 0 1020 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_400
timestamp 1581321262
transform 1 0 816 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_401
timestamp 1581321262
transform 1 0 612 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_402
timestamp 1581321262
transform 1 0 204 0 1 6593
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_403
timestamp 1581321262
transform 1 0 9588 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_404
timestamp 1581321262
transform 1 0 9384 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_405
timestamp 1581321262
transform 1 0 8160 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_406
timestamp 1581321262
transform 1 0 7956 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_407
timestamp 1581321262
transform 1 0 7548 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_408
timestamp 1581321262
transform 1 0 7140 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_409
timestamp 1581321262
transform 1 0 6936 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_410
timestamp 1581321262
transform 1 0 6324 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_411
timestamp 1581321262
transform 1 0 5916 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_412
timestamp 1581321262
transform 1 0 5508 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_413
timestamp 1581321262
transform 1 0 5304 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_414
timestamp 1581321262
transform 1 0 4284 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_415
timestamp 1581321262
transform 1 0 4080 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_416
timestamp 1581321262
transform 1 0 3876 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_417
timestamp 1581321262
transform 1 0 3468 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_418
timestamp 1581321262
transform 1 0 3264 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_419
timestamp 1581321262
transform 1 0 3060 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_420
timestamp 1581321262
transform 1 0 2652 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_421
timestamp 1581321262
transform 1 0 2244 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_422
timestamp 1581321262
transform 1 0 2040 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_423
timestamp 1581321262
transform 1 0 1836 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_424
timestamp 1581321262
transform 1 0 1632 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_425
timestamp 1581321262
transform 1 0 1428 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_426
timestamp 1581321262
transform 1 0 1224 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_427
timestamp 1581321262
transform 1 0 816 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_428
timestamp 1581321262
transform 1 0 612 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_429
timestamp 1581321262
transform 1 0 0 0 1 6389
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_430
timestamp 1581321262
transform 1 0 9588 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_431
timestamp 1581321262
transform 1 0 9384 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_432
timestamp 1581321262
transform 1 0 9180 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_433
timestamp 1581321262
transform 1 0 8772 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_434
timestamp 1581321262
transform 1 0 8364 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_435
timestamp 1581321262
transform 1 0 7956 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_436
timestamp 1581321262
transform 1 0 7548 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_437
timestamp 1581321262
transform 1 0 7140 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_438
timestamp 1581321262
transform 1 0 6732 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_439
timestamp 1581321262
transform 1 0 6324 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_440
timestamp 1581321262
transform 1 0 6120 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_441
timestamp 1581321262
transform 1 0 5508 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_442
timestamp 1581321262
transform 1 0 5304 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_443
timestamp 1581321262
transform 1 0 5100 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_444
timestamp 1581321262
transform 1 0 4896 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_445
timestamp 1581321262
transform 1 0 4692 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_446
timestamp 1581321262
transform 1 0 3672 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_447
timestamp 1581321262
transform 1 0 3264 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_448
timestamp 1581321262
transform 1 0 2856 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_449
timestamp 1581321262
transform 1 0 2652 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_450
timestamp 1581321262
transform 1 0 2448 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_451
timestamp 1581321262
transform 1 0 1836 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_452
timestamp 1581321262
transform 1 0 408 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_453
timestamp 1581321262
transform 1 0 204 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_454
timestamp 1581321262
transform 1 0 0 0 1 6185
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_455
timestamp 1581321262
transform 1 0 9384 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_456
timestamp 1581321262
transform 1 0 9180 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_457
timestamp 1581321262
transform 1 0 8772 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_458
timestamp 1581321262
transform 1 0 8568 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_459
timestamp 1581321262
transform 1 0 8364 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_460
timestamp 1581321262
transform 1 0 8160 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_461
timestamp 1581321262
transform 1 0 7752 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_462
timestamp 1581321262
transform 1 0 6528 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_463
timestamp 1581321262
transform 1 0 5916 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_464
timestamp 1581321262
transform 1 0 5712 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_465
timestamp 1581321262
transform 1 0 5304 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_466
timestamp 1581321262
transform 1 0 5100 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_467
timestamp 1581321262
transform 1 0 4080 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_468
timestamp 1581321262
transform 1 0 3672 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_469
timestamp 1581321262
transform 1 0 3264 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_470
timestamp 1581321262
transform 1 0 2652 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_471
timestamp 1581321262
transform 1 0 2244 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_472
timestamp 1581321262
transform 1 0 1836 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_473
timestamp 1581321262
transform 1 0 1632 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_474
timestamp 1581321262
transform 1 0 1428 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_475
timestamp 1581321262
transform 1 0 1020 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_476
timestamp 1581321262
transform 1 0 408 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_477
timestamp 1581321262
transform 1 0 204 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_478
timestamp 1581321262
transform 1 0 0 0 1 5877
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_479
timestamp 1581321262
transform 1 0 9588 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_480
timestamp 1581321262
transform 1 0 9384 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_481
timestamp 1581321262
transform 1 0 8976 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_482
timestamp 1581321262
transform 1 0 8772 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_483
timestamp 1581321262
transform 1 0 8160 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_484
timestamp 1581321262
transform 1 0 7956 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_485
timestamp 1581321262
transform 1 0 7140 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_486
timestamp 1581321262
transform 1 0 6120 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_487
timestamp 1581321262
transform 1 0 5916 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_488
timestamp 1581321262
transform 1 0 5712 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_489
timestamp 1581321262
transform 1 0 5508 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_490
timestamp 1581321262
transform 1 0 5304 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_491
timestamp 1581321262
transform 1 0 5100 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_492
timestamp 1581321262
transform 1 0 4896 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_493
timestamp 1581321262
transform 1 0 4284 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_494
timestamp 1581321262
transform 1 0 4080 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_495
timestamp 1581321262
transform 1 0 3876 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_496
timestamp 1581321262
transform 1 0 3264 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_497
timestamp 1581321262
transform 1 0 2652 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_498
timestamp 1581321262
transform 1 0 2244 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_499
timestamp 1581321262
transform 1 0 2040 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_500
timestamp 1581321262
transform 1 0 1836 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_501
timestamp 1581321262
transform 1 0 1632 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_502
timestamp 1581321262
transform 1 0 816 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_503
timestamp 1581321262
transform 1 0 612 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_504
timestamp 1581321262
transform 1 0 408 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_505
timestamp 1581321262
transform 1 0 204 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_506
timestamp 1581321262
transform 1 0 0 0 1 5673
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_507
timestamp 1581321262
transform 1 0 8976 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_508
timestamp 1581321262
transform 1 0 7752 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_509
timestamp 1581321262
transform 1 0 7548 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_510
timestamp 1581321262
transform 1 0 7344 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_511
timestamp 1581321262
transform 1 0 7140 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_512
timestamp 1581321262
transform 1 0 6732 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_513
timestamp 1581321262
transform 1 0 6528 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_514
timestamp 1581321262
transform 1 0 5916 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_515
timestamp 1581321262
transform 1 0 5712 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_516
timestamp 1581321262
transform 1 0 4896 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_517
timestamp 1581321262
transform 1 0 4692 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_518
timestamp 1581321262
transform 1 0 3672 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_519
timestamp 1581321262
transform 1 0 3468 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_520
timestamp 1581321262
transform 1 0 3060 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_521
timestamp 1581321262
transform 1 0 2652 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_522
timestamp 1581321262
transform 1 0 2244 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_523
timestamp 1581321262
transform 1 0 2040 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_524
timestamp 1581321262
transform 1 0 1836 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_525
timestamp 1581321262
transform 1 0 1632 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_526
timestamp 1581321262
transform 1 0 1020 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_527
timestamp 1581321262
transform 1 0 816 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_528
timestamp 1581321262
transform 1 0 612 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_529
timestamp 1581321262
transform 1 0 408 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_530
timestamp 1581321262
transform 1 0 204 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_531
timestamp 1581321262
transform 1 0 0 0 1 5469
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_532
timestamp 1581321262
transform 1 0 9180 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_533
timestamp 1581321262
transform 1 0 8976 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_534
timestamp 1581321262
transform 1 0 8772 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_535
timestamp 1581321262
transform 1 0 8364 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_536
timestamp 1581321262
transform 1 0 8160 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_537
timestamp 1581321262
transform 1 0 7956 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_538
timestamp 1581321262
transform 1 0 7548 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_539
timestamp 1581321262
transform 1 0 7140 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_540
timestamp 1581321262
transform 1 0 6732 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_541
timestamp 1581321262
transform 1 0 6324 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_542
timestamp 1581321262
transform 1 0 6120 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_543
timestamp 1581321262
transform 1 0 5916 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_544
timestamp 1581321262
transform 1 0 5304 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_545
timestamp 1581321262
transform 1 0 5100 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_546
timestamp 1581321262
transform 1 0 4692 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_547
timestamp 1581321262
transform 1 0 4284 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_548
timestamp 1581321262
transform 1 0 4080 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_549
timestamp 1581321262
transform 1 0 3264 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_550
timestamp 1581321262
transform 1 0 2856 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_551
timestamp 1581321262
transform 1 0 2652 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_552
timestamp 1581321262
transform 1 0 2448 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_553
timestamp 1581321262
transform 1 0 2040 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_554
timestamp 1581321262
transform 1 0 1836 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_555
timestamp 1581321262
transform 1 0 1632 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_556
timestamp 1581321262
transform 1 0 1224 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_557
timestamp 1581321262
transform 1 0 1020 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_558
timestamp 1581321262
transform 1 0 612 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_559
timestamp 1581321262
transform 1 0 408 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_560
timestamp 1581321262
transform 1 0 204 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_561
timestamp 1581321262
transform 1 0 0 0 1 5265
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_562
timestamp 1581321262
transform 1 0 7956 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_563
timestamp 1581321262
transform 1 0 7752 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_564
timestamp 1581321262
transform 1 0 7548 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_565
timestamp 1581321262
transform 1 0 7344 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_566
timestamp 1581321262
transform 1 0 7140 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_567
timestamp 1581321262
transform 1 0 6936 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_568
timestamp 1581321262
transform 1 0 6528 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_569
timestamp 1581321262
transform 1 0 5712 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_570
timestamp 1581321262
transform 1 0 5304 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_571
timestamp 1581321262
transform 1 0 4080 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_572
timestamp 1581321262
transform 1 0 3876 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_573
timestamp 1581321262
transform 1 0 3468 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_574
timestamp 1581321262
transform 1 0 3060 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_575
timestamp 1581321262
transform 1 0 2856 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_576
timestamp 1581321262
transform 1 0 2652 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_577
timestamp 1581321262
transform 1 0 1836 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_578
timestamp 1581321262
transform 1 0 1632 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_579
timestamp 1581321262
transform 1 0 1428 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_580
timestamp 1581321262
transform 1 0 1224 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_581
timestamp 1581321262
transform 1 0 1020 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_582
timestamp 1581321262
transform 1 0 612 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_583
timestamp 1581321262
transform 1 0 0 0 1 5061
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_584
timestamp 1581321262
transform 1 0 9588 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_585
timestamp 1581321262
transform 1 0 8976 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_586
timestamp 1581321262
transform 1 0 8568 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_587
timestamp 1581321262
transform 1 0 8364 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_588
timestamp 1581321262
transform 1 0 7956 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_589
timestamp 1581321262
transform 1 0 7752 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_590
timestamp 1581321262
transform 1 0 7548 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_591
timestamp 1581321262
transform 1 0 7140 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_592
timestamp 1581321262
transform 1 0 6936 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_593
timestamp 1581321262
transform 1 0 6324 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_594
timestamp 1581321262
transform 1 0 6120 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_595
timestamp 1581321262
transform 1 0 4896 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_596
timestamp 1581321262
transform 1 0 4692 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_597
timestamp 1581321262
transform 1 0 2856 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_598
timestamp 1581321262
transform 1 0 2244 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_599
timestamp 1581321262
transform 1 0 1632 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_600
timestamp 1581321262
transform 1 0 612 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_601
timestamp 1581321262
transform 1 0 204 0 1 4857
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_602
timestamp 1581321262
transform 1 0 9588 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_603
timestamp 1581321262
transform 1 0 8976 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_604
timestamp 1581321262
transform 1 0 8568 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_605
timestamp 1581321262
transform 1 0 8364 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_606
timestamp 1581321262
transform 1 0 8160 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_607
timestamp 1581321262
transform 1 0 7548 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_608
timestamp 1581321262
transform 1 0 7140 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_609
timestamp 1581321262
transform 1 0 6936 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_610
timestamp 1581321262
transform 1 0 6732 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_611
timestamp 1581321262
transform 1 0 6528 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_612
timestamp 1581321262
transform 1 0 6324 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_613
timestamp 1581321262
transform 1 0 5712 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_614
timestamp 1581321262
transform 1 0 5100 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_615
timestamp 1581321262
transform 1 0 4896 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_616
timestamp 1581321262
transform 1 0 4488 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_617
timestamp 1581321262
transform 1 0 4284 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_618
timestamp 1581321262
transform 1 0 3876 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_619
timestamp 1581321262
transform 1 0 3264 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_620
timestamp 1581321262
transform 1 0 2856 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_621
timestamp 1581321262
transform 1 0 2652 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_622
timestamp 1581321262
transform 1 0 2448 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_623
timestamp 1581321262
transform 1 0 2244 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_624
timestamp 1581321262
transform 1 0 1836 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_625
timestamp 1581321262
transform 1 0 1224 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_626
timestamp 1581321262
transform 1 0 1020 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_627
timestamp 1581321262
transform 1 0 816 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_628
timestamp 1581321262
transform 1 0 408 0 1 4653
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_629
timestamp 1581321262
transform 1 0 9384 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_630
timestamp 1581321262
transform 1 0 9180 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_631
timestamp 1581321262
transform 1 0 8976 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_632
timestamp 1581321262
transform 1 0 8364 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_633
timestamp 1581321262
transform 1 0 8160 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_634
timestamp 1581321262
transform 1 0 7752 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_635
timestamp 1581321262
transform 1 0 7548 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_636
timestamp 1581321262
transform 1 0 6324 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_637
timestamp 1581321262
transform 1 0 5916 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_638
timestamp 1581321262
transform 1 0 5508 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_639
timestamp 1581321262
transform 1 0 5304 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_640
timestamp 1581321262
transform 1 0 5100 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_641
timestamp 1581321262
transform 1 0 4896 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_642
timestamp 1581321262
transform 1 0 4692 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_643
timestamp 1581321262
transform 1 0 4284 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_644
timestamp 1581321262
transform 1 0 4080 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_645
timestamp 1581321262
transform 1 0 3876 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_646
timestamp 1581321262
transform 1 0 3672 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_647
timestamp 1581321262
transform 1 0 3468 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_648
timestamp 1581321262
transform 1 0 3264 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_649
timestamp 1581321262
transform 1 0 3060 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_650
timestamp 1581321262
transform 1 0 2652 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_651
timestamp 1581321262
transform 1 0 2244 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_652
timestamp 1581321262
transform 1 0 1428 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_653
timestamp 1581321262
transform 1 0 1224 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_654
timestamp 1581321262
transform 1 0 1020 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_655
timestamp 1581321262
transform 1 0 612 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_656
timestamp 1581321262
transform 1 0 204 0 1 4449
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_657
timestamp 1581321262
transform 1 0 9588 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_658
timestamp 1581321262
transform 1 0 9180 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_659
timestamp 1581321262
transform 1 0 8772 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_660
timestamp 1581321262
transform 1 0 8568 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_661
timestamp 1581321262
transform 1 0 8364 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_662
timestamp 1581321262
transform 1 0 8160 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_663
timestamp 1581321262
transform 1 0 6528 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_664
timestamp 1581321262
transform 1 0 6120 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_665
timestamp 1581321262
transform 1 0 4692 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_666
timestamp 1581321262
transform 1 0 4488 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_667
timestamp 1581321262
transform 1 0 4080 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_668
timestamp 1581321262
transform 1 0 3672 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_669
timestamp 1581321262
transform 1 0 3468 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_670
timestamp 1581321262
transform 1 0 3060 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_671
timestamp 1581321262
transform 1 0 2652 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_672
timestamp 1581321262
transform 1 0 2244 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_673
timestamp 1581321262
transform 1 0 1836 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_674
timestamp 1581321262
transform 1 0 1632 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_675
timestamp 1581321262
transform 1 0 1020 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_676
timestamp 1581321262
transform 1 0 612 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_677
timestamp 1581321262
transform 1 0 204 0 1 4141
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_678
timestamp 1581321262
transform 1 0 9588 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_679
timestamp 1581321262
transform 1 0 9384 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_680
timestamp 1581321262
transform 1 0 9180 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_681
timestamp 1581321262
transform 1 0 8976 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_682
timestamp 1581321262
transform 1 0 8568 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_683
timestamp 1581321262
transform 1 0 8364 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_684
timestamp 1581321262
transform 1 0 8160 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_685
timestamp 1581321262
transform 1 0 7752 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_686
timestamp 1581321262
transform 1 0 7344 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_687
timestamp 1581321262
transform 1 0 6936 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_688
timestamp 1581321262
transform 1 0 5916 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_689
timestamp 1581321262
transform 1 0 5712 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_690
timestamp 1581321262
transform 1 0 4896 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_691
timestamp 1581321262
transform 1 0 4692 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_692
timestamp 1581321262
transform 1 0 4488 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_693
timestamp 1581321262
transform 1 0 4284 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_694
timestamp 1581321262
transform 1 0 4080 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_695
timestamp 1581321262
transform 1 0 3876 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_696
timestamp 1581321262
transform 1 0 3060 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_697
timestamp 1581321262
transform 1 0 2652 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_698
timestamp 1581321262
transform 1 0 2040 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_699
timestamp 1581321262
transform 1 0 1836 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_700
timestamp 1581321262
transform 1 0 1632 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_701
timestamp 1581321262
transform 1 0 1428 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_702
timestamp 1581321262
transform 1 0 1224 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_703
timestamp 1581321262
transform 1 0 816 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_704
timestamp 1581321262
transform 1 0 408 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_705
timestamp 1581321262
transform 1 0 0 0 1 3937
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_706
timestamp 1581321262
transform 1 0 9180 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_707
timestamp 1581321262
transform 1 0 8772 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_708
timestamp 1581321262
transform 1 0 8568 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_709
timestamp 1581321262
transform 1 0 8160 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_710
timestamp 1581321262
transform 1 0 7140 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_711
timestamp 1581321262
transform 1 0 6936 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_712
timestamp 1581321262
transform 1 0 6732 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_713
timestamp 1581321262
transform 1 0 6120 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_714
timestamp 1581321262
transform 1 0 5304 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_715
timestamp 1581321262
transform 1 0 4692 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_716
timestamp 1581321262
transform 1 0 4080 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_717
timestamp 1581321262
transform 1 0 3876 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_718
timestamp 1581321262
transform 1 0 3672 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_719
timestamp 1581321262
transform 1 0 3060 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_720
timestamp 1581321262
transform 1 0 2448 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_721
timestamp 1581321262
transform 1 0 2244 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_722
timestamp 1581321262
transform 1 0 2040 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_723
timestamp 1581321262
transform 1 0 1836 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_724
timestamp 1581321262
transform 1 0 1020 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_725
timestamp 1581321262
transform 1 0 816 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_726
timestamp 1581321262
transform 1 0 612 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_727
timestamp 1581321262
transform 1 0 408 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_728
timestamp 1581321262
transform 1 0 204 0 1 3733
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_729
timestamp 1581321262
transform 1 0 9588 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_730
timestamp 1581321262
transform 1 0 9384 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_731
timestamp 1581321262
transform 1 0 8976 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_732
timestamp 1581321262
transform 1 0 8568 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_733
timestamp 1581321262
transform 1 0 7956 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_734
timestamp 1581321262
transform 1 0 7548 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_735
timestamp 1581321262
transform 1 0 7344 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_736
timestamp 1581321262
transform 1 0 7140 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_737
timestamp 1581321262
transform 1 0 6936 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_738
timestamp 1581321262
transform 1 0 6732 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_739
timestamp 1581321262
transform 1 0 6528 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_740
timestamp 1581321262
transform 1 0 6324 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_741
timestamp 1581321262
transform 1 0 6120 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_742
timestamp 1581321262
transform 1 0 5916 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_743
timestamp 1581321262
transform 1 0 5304 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_744
timestamp 1581321262
transform 1 0 4692 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_745
timestamp 1581321262
transform 1 0 4080 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_746
timestamp 1581321262
transform 1 0 3876 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_747
timestamp 1581321262
transform 1 0 2856 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_748
timestamp 1581321262
transform 1 0 2244 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_749
timestamp 1581321262
transform 1 0 1836 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_750
timestamp 1581321262
transform 1 0 1428 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_751
timestamp 1581321262
transform 1 0 1224 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_752
timestamp 1581321262
transform 1 0 1020 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_753
timestamp 1581321262
transform 1 0 816 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_754
timestamp 1581321262
transform 1 0 612 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_755
timestamp 1581321262
transform 1 0 408 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_756
timestamp 1581321262
transform 1 0 0 0 1 3529
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_757
timestamp 1581321262
transform 1 0 9588 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_758
timestamp 1581321262
transform 1 0 9384 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_759
timestamp 1581321262
transform 1 0 8568 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_760
timestamp 1581321262
transform 1 0 7956 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_761
timestamp 1581321262
transform 1 0 7752 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_762
timestamp 1581321262
transform 1 0 7344 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_763
timestamp 1581321262
transform 1 0 7140 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_764
timestamp 1581321262
transform 1 0 6732 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_765
timestamp 1581321262
transform 1 0 6528 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_766
timestamp 1581321262
transform 1 0 6120 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_767
timestamp 1581321262
transform 1 0 5916 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_768
timestamp 1581321262
transform 1 0 5712 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_769
timestamp 1581321262
transform 1 0 3672 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_770
timestamp 1581321262
transform 1 0 3060 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_771
timestamp 1581321262
transform 1 0 2856 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_772
timestamp 1581321262
transform 1 0 2244 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_773
timestamp 1581321262
transform 1 0 2040 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_774
timestamp 1581321262
transform 1 0 1836 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_775
timestamp 1581321262
transform 1 0 1632 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_776
timestamp 1581321262
transform 1 0 408 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_777
timestamp 1581321262
transform 1 0 0 0 1 3325
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_778
timestamp 1581321262
transform 1 0 9384 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_779
timestamp 1581321262
transform 1 0 8772 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_780
timestamp 1581321262
transform 1 0 8364 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_781
timestamp 1581321262
transform 1 0 7956 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_782
timestamp 1581321262
transform 1 0 7548 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_783
timestamp 1581321262
transform 1 0 6528 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_784
timestamp 1581321262
transform 1 0 6120 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_785
timestamp 1581321262
transform 1 0 5916 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_786
timestamp 1581321262
transform 1 0 5508 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_787
timestamp 1581321262
transform 1 0 5100 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_788
timestamp 1581321262
transform 1 0 4692 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_789
timestamp 1581321262
transform 1 0 4080 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_790
timestamp 1581321262
transform 1 0 3876 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_791
timestamp 1581321262
transform 1 0 3672 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_792
timestamp 1581321262
transform 1 0 3264 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_793
timestamp 1581321262
transform 1 0 3060 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_794
timestamp 1581321262
transform 1 0 2856 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_795
timestamp 1581321262
transform 1 0 2652 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_796
timestamp 1581321262
transform 1 0 2448 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_797
timestamp 1581321262
transform 1 0 2244 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_798
timestamp 1581321262
transform 1 0 1836 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_799
timestamp 1581321262
transform 1 0 1224 0 1 3121
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_800
timestamp 1581321262
transform 1 0 9384 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_801
timestamp 1581321262
transform 1 0 9180 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_802
timestamp 1581321262
transform 1 0 8772 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_803
timestamp 1581321262
transform 1 0 7752 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_804
timestamp 1581321262
transform 1 0 7140 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_805
timestamp 1581321262
transform 1 0 6324 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_806
timestamp 1581321262
transform 1 0 5916 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_807
timestamp 1581321262
transform 1 0 4692 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_808
timestamp 1581321262
transform 1 0 3672 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_809
timestamp 1581321262
transform 1 0 3264 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_810
timestamp 1581321262
transform 1 0 3060 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_811
timestamp 1581321262
transform 1 0 2856 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_812
timestamp 1581321262
transform 1 0 2448 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_813
timestamp 1581321262
transform 1 0 2244 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_814
timestamp 1581321262
transform 1 0 1632 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_815
timestamp 1581321262
transform 1 0 1428 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_816
timestamp 1581321262
transform 1 0 1020 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_817
timestamp 1581321262
transform 1 0 816 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_818
timestamp 1581321262
transform 1 0 612 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_819
timestamp 1581321262
transform 1 0 408 0 1 2917
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_820
timestamp 1581321262
transform 1 0 9588 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_821
timestamp 1581321262
transform 1 0 9384 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_822
timestamp 1581321262
transform 1 0 9180 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_823
timestamp 1581321262
transform 1 0 8772 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_824
timestamp 1581321262
transform 1 0 7548 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_825
timestamp 1581321262
transform 1 0 6528 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_826
timestamp 1581321262
transform 1 0 5508 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_827
timestamp 1581321262
transform 1 0 5100 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_828
timestamp 1581321262
transform 1 0 4692 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_829
timestamp 1581321262
transform 1 0 4284 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_830
timestamp 1581321262
transform 1 0 4080 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_831
timestamp 1581321262
transform 1 0 3876 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_832
timestamp 1581321262
transform 1 0 3468 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_833
timestamp 1581321262
transform 1 0 3060 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_834
timestamp 1581321262
transform 1 0 2856 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_835
timestamp 1581321262
transform 1 0 2448 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_836
timestamp 1581321262
transform 1 0 2244 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_837
timestamp 1581321262
transform 1 0 1632 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_838
timestamp 1581321262
transform 1 0 1428 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_839
timestamp 1581321262
transform 1 0 1020 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_840
timestamp 1581321262
transform 1 0 204 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_841
timestamp 1581321262
transform 1 0 0 0 1 2713
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_842
timestamp 1581321262
transform 1 0 9384 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_843
timestamp 1581321262
transform 1 0 9180 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_844
timestamp 1581321262
transform 1 0 8772 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_845
timestamp 1581321262
transform 1 0 8364 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_846
timestamp 1581321262
transform 1 0 7752 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_847
timestamp 1581321262
transform 1 0 7140 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_848
timestamp 1581321262
transform 1 0 6936 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_849
timestamp 1581321262
transform 1 0 6528 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_850
timestamp 1581321262
transform 1 0 6324 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_851
timestamp 1581321262
transform 1 0 5712 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_852
timestamp 1581321262
transform 1 0 5508 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_853
timestamp 1581321262
transform 1 0 5100 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_854
timestamp 1581321262
transform 1 0 4080 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_855
timestamp 1581321262
transform 1 0 3876 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_856
timestamp 1581321262
transform 1 0 3672 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_857
timestamp 1581321262
transform 1 0 2652 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_858
timestamp 1581321262
transform 1 0 2448 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_859
timestamp 1581321262
transform 1 0 1836 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_860
timestamp 1581321262
transform 1 0 1428 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_861
timestamp 1581321262
transform 1 0 1224 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_862
timestamp 1581321262
transform 1 0 612 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_863
timestamp 1581321262
transform 1 0 408 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_864
timestamp 1581321262
transform 1 0 204 0 1 2405
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_865
timestamp 1581321262
transform 1 0 8976 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_866
timestamp 1581321262
transform 1 0 8772 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_867
timestamp 1581321262
transform 1 0 8364 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_868
timestamp 1581321262
transform 1 0 8160 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_869
timestamp 1581321262
transform 1 0 7956 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_870
timestamp 1581321262
transform 1 0 7752 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_871
timestamp 1581321262
transform 1 0 7548 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_872
timestamp 1581321262
transform 1 0 7344 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_873
timestamp 1581321262
transform 1 0 6936 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_874
timestamp 1581321262
transform 1 0 6732 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_875
timestamp 1581321262
transform 1 0 6324 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_876
timestamp 1581321262
transform 1 0 6120 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_877
timestamp 1581321262
transform 1 0 5916 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_878
timestamp 1581321262
transform 1 0 5712 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_879
timestamp 1581321262
transform 1 0 5508 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_880
timestamp 1581321262
transform 1 0 5304 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_881
timestamp 1581321262
transform 1 0 5100 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_882
timestamp 1581321262
transform 1 0 4692 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_883
timestamp 1581321262
transform 1 0 4284 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_884
timestamp 1581321262
transform 1 0 4080 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_885
timestamp 1581321262
transform 1 0 3264 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_886
timestamp 1581321262
transform 1 0 3060 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_887
timestamp 1581321262
transform 1 0 2856 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_888
timestamp 1581321262
transform 1 0 2448 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_889
timestamp 1581321262
transform 1 0 2244 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_890
timestamp 1581321262
transform 1 0 1428 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_891
timestamp 1581321262
transform 1 0 1224 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_892
timestamp 1581321262
transform 1 0 1020 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_893
timestamp 1581321262
transform 1 0 612 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_894
timestamp 1581321262
transform 1 0 408 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_895
timestamp 1581321262
transform 1 0 204 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_896
timestamp 1581321262
transform 1 0 0 0 1 2201
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_897
timestamp 1581321262
transform 1 0 9588 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_898
timestamp 1581321262
transform 1 0 8976 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_899
timestamp 1581321262
transform 1 0 8568 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_900
timestamp 1581321262
transform 1 0 8364 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_901
timestamp 1581321262
transform 1 0 7548 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_902
timestamp 1581321262
transform 1 0 7344 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_903
timestamp 1581321262
transform 1 0 6936 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_904
timestamp 1581321262
transform 1 0 6528 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_905
timestamp 1581321262
transform 1 0 6324 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_906
timestamp 1581321262
transform 1 0 6120 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_907
timestamp 1581321262
transform 1 0 5916 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_908
timestamp 1581321262
transform 1 0 5712 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_909
timestamp 1581321262
transform 1 0 5100 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_910
timestamp 1581321262
transform 1 0 4692 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_911
timestamp 1581321262
transform 1 0 4488 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_912
timestamp 1581321262
transform 1 0 4284 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_913
timestamp 1581321262
transform 1 0 3876 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_914
timestamp 1581321262
transform 1 0 3468 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_915
timestamp 1581321262
transform 1 0 3264 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_916
timestamp 1581321262
transform 1 0 2244 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_917
timestamp 1581321262
transform 1 0 1428 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_918
timestamp 1581321262
transform 1 0 1224 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_919
timestamp 1581321262
transform 1 0 1020 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_920
timestamp 1581321262
transform 1 0 0 0 1 1997
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_921
timestamp 1581321262
transform 1 0 9588 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_922
timestamp 1581321262
transform 1 0 9384 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_923
timestamp 1581321262
transform 1 0 8976 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_924
timestamp 1581321262
transform 1 0 8772 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_925
timestamp 1581321262
transform 1 0 7548 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_926
timestamp 1581321262
transform 1 0 6936 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_927
timestamp 1581321262
transform 1 0 6528 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_928
timestamp 1581321262
transform 1 0 5916 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_929
timestamp 1581321262
transform 1 0 5712 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_930
timestamp 1581321262
transform 1 0 5508 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_931
timestamp 1581321262
transform 1 0 5304 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_932
timestamp 1581321262
transform 1 0 4896 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_933
timestamp 1581321262
transform 1 0 4488 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_934
timestamp 1581321262
transform 1 0 4284 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_935
timestamp 1581321262
transform 1 0 3468 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_936
timestamp 1581321262
transform 1 0 3264 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_937
timestamp 1581321262
transform 1 0 3060 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_938
timestamp 1581321262
transform 1 0 2652 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_939
timestamp 1581321262
transform 1 0 2448 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_940
timestamp 1581321262
transform 1 0 2244 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_941
timestamp 1581321262
transform 1 0 2040 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_942
timestamp 1581321262
transform 1 0 1428 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_943
timestamp 1581321262
transform 1 0 1224 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_944
timestamp 1581321262
transform 1 0 1020 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_945
timestamp 1581321262
transform 1 0 816 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_946
timestamp 1581321262
transform 1 0 612 0 1 1793
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_947
timestamp 1581321262
transform 1 0 8976 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_948
timestamp 1581321262
transform 1 0 8772 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_949
timestamp 1581321262
transform 1 0 8364 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_950
timestamp 1581321262
transform 1 0 8160 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_951
timestamp 1581321262
transform 1 0 7956 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_952
timestamp 1581321262
transform 1 0 7752 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_953
timestamp 1581321262
transform 1 0 7548 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_954
timestamp 1581321262
transform 1 0 6120 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_955
timestamp 1581321262
transform 1 0 4896 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_956
timestamp 1581321262
transform 1 0 4284 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_957
timestamp 1581321262
transform 1 0 4080 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_958
timestamp 1581321262
transform 1 0 3876 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_959
timestamp 1581321262
transform 1 0 3468 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_960
timestamp 1581321262
transform 1 0 3264 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_961
timestamp 1581321262
transform 1 0 3060 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_962
timestamp 1581321262
transform 1 0 2856 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_963
timestamp 1581321262
transform 1 0 2448 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_964
timestamp 1581321262
transform 1 0 1836 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_965
timestamp 1581321262
transform 1 0 1632 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_966
timestamp 1581321262
transform 1 0 1428 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_967
timestamp 1581321262
transform 1 0 1224 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_968
timestamp 1581321262
transform 1 0 1020 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_969
timestamp 1581321262
transform 1 0 408 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_970
timestamp 1581321262
transform 1 0 204 0 1 1589
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_971
timestamp 1581321262
transform 1 0 9588 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_972
timestamp 1581321262
transform 1 0 8772 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_973
timestamp 1581321262
transform 1 0 8568 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_974
timestamp 1581321262
transform 1 0 7752 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_975
timestamp 1581321262
transform 1 0 7548 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_976
timestamp 1581321262
transform 1 0 7344 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_977
timestamp 1581321262
transform 1 0 6936 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_978
timestamp 1581321262
transform 1 0 6528 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_979
timestamp 1581321262
transform 1 0 5712 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_980
timestamp 1581321262
transform 1 0 5508 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_981
timestamp 1581321262
transform 1 0 5304 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_982
timestamp 1581321262
transform 1 0 4080 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_983
timestamp 1581321262
transform 1 0 3672 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_984
timestamp 1581321262
transform 1 0 3468 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_985
timestamp 1581321262
transform 1 0 3264 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_986
timestamp 1581321262
transform 1 0 3060 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_987
timestamp 1581321262
transform 1 0 1836 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_988
timestamp 1581321262
transform 1 0 1428 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_989
timestamp 1581321262
transform 1 0 1020 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_990
timestamp 1581321262
transform 1 0 408 0 1 1385
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_991
timestamp 1581321262
transform 1 0 9384 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_992
timestamp 1581321262
transform 1 0 8772 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_993
timestamp 1581321262
transform 1 0 8568 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_994
timestamp 1581321262
transform 1 0 8160 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_995
timestamp 1581321262
transform 1 0 7956 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_996
timestamp 1581321262
transform 1 0 7548 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_997
timestamp 1581321262
transform 1 0 7344 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_998
timestamp 1581321262
transform 1 0 7140 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_999
timestamp 1581321262
transform 1 0 6936 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1000
timestamp 1581321262
transform 1 0 6528 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1001
timestamp 1581321262
transform 1 0 6324 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1002
timestamp 1581321262
transform 1 0 6120 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1003
timestamp 1581321262
transform 1 0 5508 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1004
timestamp 1581321262
transform 1 0 4284 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1005
timestamp 1581321262
transform 1 0 3876 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1006
timestamp 1581321262
transform 1 0 3672 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1007
timestamp 1581321262
transform 1 0 3468 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1008
timestamp 1581321262
transform 1 0 2652 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1009
timestamp 1581321262
transform 1 0 2448 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1010
timestamp 1581321262
transform 1 0 1836 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1011
timestamp 1581321262
transform 1 0 1224 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1012
timestamp 1581321262
transform 1 0 816 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1013
timestamp 1581321262
transform 1 0 0 0 1 1181
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1014
timestamp 1581321262
transform 1 0 9384 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1015
timestamp 1581321262
transform 1 0 9180 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1016
timestamp 1581321262
transform 1 0 8772 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1017
timestamp 1581321262
transform 1 0 8160 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1018
timestamp 1581321262
transform 1 0 7956 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1019
timestamp 1581321262
transform 1 0 7752 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1020
timestamp 1581321262
transform 1 0 6732 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1021
timestamp 1581321262
transform 1 0 6324 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1022
timestamp 1581321262
transform 1 0 6120 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1023
timestamp 1581321262
transform 1 0 5916 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1024
timestamp 1581321262
transform 1 0 5712 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1025
timestamp 1581321262
transform 1 0 5508 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1026
timestamp 1581321262
transform 1 0 5304 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1027
timestamp 1581321262
transform 1 0 4284 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1028
timestamp 1581321262
transform 1 0 4080 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1029
timestamp 1581321262
transform 1 0 3468 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1030
timestamp 1581321262
transform 1 0 3060 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1031
timestamp 1581321262
transform 1 0 2856 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1032
timestamp 1581321262
transform 1 0 2448 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1033
timestamp 1581321262
transform 1 0 2040 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1034
timestamp 1581321262
transform 1 0 1836 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1035
timestamp 1581321262
transform 1 0 1224 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1036
timestamp 1581321262
transform 1 0 816 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1037
timestamp 1581321262
transform 1 0 408 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1038
timestamp 1581321262
transform 1 0 204 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_base_zero_cell  sky130_rom_krom_rom_base_zero_cell_1039
timestamp 1581321262
transform 1 0 0 0 1 977
box 0 -51 204 204
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_0
timestamp 1581321262
transform 1 0 9792 0 1 10065
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_1
timestamp 1581321262
transform 1 0 8160 0 1 10065
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_2
timestamp 1581321262
transform 1 0 6528 0 1 10065
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_3
timestamp 1581321262
transform 1 0 4896 0 1 10065
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_4
timestamp 1581321262
transform 1 0 3264 0 1 10065
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_5
timestamp 1581321262
transform 1 0 1632 0 1 10065
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_6
timestamp 1581321262
transform 1 0 0 0 1 10065
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_7
timestamp 1581321262
transform 1 0 9792 0 1 9861
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_8
timestamp 1581321262
transform 1 0 8160 0 1 9861
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_9
timestamp 1581321262
transform 1 0 6528 0 1 9861
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_10
timestamp 1581321262
transform 1 0 4896 0 1 9861
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_11
timestamp 1581321262
transform 1 0 3264 0 1 9861
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_12
timestamp 1581321262
transform 1 0 1632 0 1 9861
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_13
timestamp 1581321262
transform 1 0 0 0 1 9861
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_14
timestamp 1581321262
transform 1 0 9792 0 1 9657
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_15
timestamp 1581321262
transform 1 0 8160 0 1 9657
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_16
timestamp 1581321262
transform 1 0 6528 0 1 9657
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_17
timestamp 1581321262
transform 1 0 4896 0 1 9657
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_18
timestamp 1581321262
transform 1 0 3264 0 1 9657
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_19
timestamp 1581321262
transform 1 0 1632 0 1 9657
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_20
timestamp 1581321262
transform 1 0 0 0 1 9657
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_21
timestamp 1581321262
transform 1 0 9792 0 1 9349
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_22
timestamp 1581321262
transform 1 0 8160 0 1 9349
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_23
timestamp 1581321262
transform 1 0 6528 0 1 9349
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_24
timestamp 1581321262
transform 1 0 4896 0 1 9349
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_25
timestamp 1581321262
transform 1 0 3264 0 1 9349
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_26
timestamp 1581321262
transform 1 0 1632 0 1 9349
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_27
timestamp 1581321262
transform 1 0 0 0 1 9349
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_28
timestamp 1581321262
transform 1 0 9792 0 1 9145
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_29
timestamp 1581321262
transform 1 0 8160 0 1 9145
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_30
timestamp 1581321262
transform 1 0 6528 0 1 9145
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_31
timestamp 1581321262
transform 1 0 4896 0 1 9145
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_32
timestamp 1581321262
transform 1 0 3264 0 1 9145
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_33
timestamp 1581321262
transform 1 0 1632 0 1 9145
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_34
timestamp 1581321262
transform 1 0 0 0 1 9145
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_35
timestamp 1581321262
transform 1 0 9792 0 1 8941
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_36
timestamp 1581321262
transform 1 0 8160 0 1 8941
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_37
timestamp 1581321262
transform 1 0 6528 0 1 8941
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_38
timestamp 1581321262
transform 1 0 4896 0 1 8941
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_39
timestamp 1581321262
transform 1 0 3264 0 1 8941
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_40
timestamp 1581321262
transform 1 0 1632 0 1 8941
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_41
timestamp 1581321262
transform 1 0 0 0 1 8941
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_42
timestamp 1581321262
transform 1 0 9792 0 1 8737
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_43
timestamp 1581321262
transform 1 0 8160 0 1 8737
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_44
timestamp 1581321262
transform 1 0 6528 0 1 8737
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_45
timestamp 1581321262
transform 1 0 4896 0 1 8737
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_46
timestamp 1581321262
transform 1 0 3264 0 1 8737
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_47
timestamp 1581321262
transform 1 0 1632 0 1 8737
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_48
timestamp 1581321262
transform 1 0 0 0 1 8737
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_49
timestamp 1581321262
transform 1 0 9792 0 1 8533
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_50
timestamp 1581321262
transform 1 0 8160 0 1 8533
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_51
timestamp 1581321262
transform 1 0 6528 0 1 8533
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_52
timestamp 1581321262
transform 1 0 4896 0 1 8533
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_53
timestamp 1581321262
transform 1 0 3264 0 1 8533
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_54
timestamp 1581321262
transform 1 0 1632 0 1 8533
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_55
timestamp 1581321262
transform 1 0 0 0 1 8533
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_56
timestamp 1581321262
transform 1 0 9792 0 1 8329
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_57
timestamp 1581321262
transform 1 0 8160 0 1 8329
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_58
timestamp 1581321262
transform 1 0 6528 0 1 8329
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_59
timestamp 1581321262
transform 1 0 4896 0 1 8329
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_60
timestamp 1581321262
transform 1 0 3264 0 1 8329
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_61
timestamp 1581321262
transform 1 0 1632 0 1 8329
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_62
timestamp 1581321262
transform 1 0 0 0 1 8329
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_63
timestamp 1581321262
transform 1 0 9792 0 1 8125
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_64
timestamp 1581321262
transform 1 0 8160 0 1 8125
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_65
timestamp 1581321262
transform 1 0 6528 0 1 8125
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_66
timestamp 1581321262
transform 1 0 4896 0 1 8125
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_67
timestamp 1581321262
transform 1 0 3264 0 1 8125
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_68
timestamp 1581321262
transform 1 0 1632 0 1 8125
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_69
timestamp 1581321262
transform 1 0 0 0 1 8125
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_70
timestamp 1581321262
transform 1 0 9792 0 1 7921
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_71
timestamp 1581321262
transform 1 0 8160 0 1 7921
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_72
timestamp 1581321262
transform 1 0 6528 0 1 7921
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_73
timestamp 1581321262
transform 1 0 4896 0 1 7921
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_74
timestamp 1581321262
transform 1 0 3264 0 1 7921
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_75
timestamp 1581321262
transform 1 0 1632 0 1 7921
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_76
timestamp 1581321262
transform 1 0 0 0 1 7921
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_77
timestamp 1581321262
transform 1 0 9792 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_78
timestamp 1581321262
transform 1 0 8160 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_79
timestamp 1581321262
transform 1 0 6528 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_80
timestamp 1581321262
transform 1 0 4896 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_81
timestamp 1581321262
transform 1 0 3264 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_82
timestamp 1581321262
transform 1 0 1632 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_83
timestamp 1581321262
transform 1 0 0 0 1 7613
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_84
timestamp 1581321262
transform 1 0 9792 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_85
timestamp 1581321262
transform 1 0 8160 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_86
timestamp 1581321262
transform 1 0 6528 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_87
timestamp 1581321262
transform 1 0 4896 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_88
timestamp 1581321262
transform 1 0 3264 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_89
timestamp 1581321262
transform 1 0 1632 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_90
timestamp 1581321262
transform 1 0 0 0 1 7409
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_91
timestamp 1581321262
transform 1 0 9792 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_92
timestamp 1581321262
transform 1 0 8160 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_93
timestamp 1581321262
transform 1 0 6528 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_94
timestamp 1581321262
transform 1 0 4896 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_95
timestamp 1581321262
transform 1 0 3264 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_96
timestamp 1581321262
transform 1 0 1632 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_97
timestamp 1581321262
transform 1 0 0 0 1 7205
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_98
timestamp 1581321262
transform 1 0 9792 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_99
timestamp 1581321262
transform 1 0 8160 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_100
timestamp 1581321262
transform 1 0 6528 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_101
timestamp 1581321262
transform 1 0 4896 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_102
timestamp 1581321262
transform 1 0 3264 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_103
timestamp 1581321262
transform 1 0 1632 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_104
timestamp 1581321262
transform 1 0 0 0 1 7001
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_105
timestamp 1581321262
transform 1 0 9792 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_106
timestamp 1581321262
transform 1 0 8160 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_107
timestamp 1581321262
transform 1 0 6528 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_108
timestamp 1581321262
transform 1 0 4896 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_109
timestamp 1581321262
transform 1 0 3264 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_110
timestamp 1581321262
transform 1 0 1632 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_111
timestamp 1581321262
transform 1 0 0 0 1 6797
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_112
timestamp 1581321262
transform 1 0 9792 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_113
timestamp 1581321262
transform 1 0 8160 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_114
timestamp 1581321262
transform 1 0 6528 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_115
timestamp 1581321262
transform 1 0 4896 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_116
timestamp 1581321262
transform 1 0 3264 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_117
timestamp 1581321262
transform 1 0 1632 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_118
timestamp 1581321262
transform 1 0 0 0 1 6593
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_119
timestamp 1581321262
transform 1 0 9792 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_120
timestamp 1581321262
transform 1 0 8160 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_121
timestamp 1581321262
transform 1 0 6528 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_122
timestamp 1581321262
transform 1 0 4896 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_123
timestamp 1581321262
transform 1 0 3264 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_124
timestamp 1581321262
transform 1 0 1632 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_125
timestamp 1581321262
transform 1 0 0 0 1 6389
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_126
timestamp 1581321262
transform 1 0 9792 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_127
timestamp 1581321262
transform 1 0 8160 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_128
timestamp 1581321262
transform 1 0 6528 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_129
timestamp 1581321262
transform 1 0 4896 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_130
timestamp 1581321262
transform 1 0 3264 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_131
timestamp 1581321262
transform 1 0 1632 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_132
timestamp 1581321262
transform 1 0 0 0 1 6185
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_133
timestamp 1581321262
transform 1 0 9792 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_134
timestamp 1581321262
transform 1 0 8160 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_135
timestamp 1581321262
transform 1 0 6528 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_136
timestamp 1581321262
transform 1 0 4896 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_137
timestamp 1581321262
transform 1 0 3264 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_138
timestamp 1581321262
transform 1 0 1632 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_139
timestamp 1581321262
transform 1 0 0 0 1 5877
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_140
timestamp 1581321262
transform 1 0 9792 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_141
timestamp 1581321262
transform 1 0 8160 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_142
timestamp 1581321262
transform 1 0 6528 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_143
timestamp 1581321262
transform 1 0 4896 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_144
timestamp 1581321262
transform 1 0 3264 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_145
timestamp 1581321262
transform 1 0 1632 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_146
timestamp 1581321262
transform 1 0 0 0 1 5673
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_147
timestamp 1581321262
transform 1 0 9792 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_148
timestamp 1581321262
transform 1 0 8160 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_149
timestamp 1581321262
transform 1 0 6528 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_150
timestamp 1581321262
transform 1 0 4896 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_151
timestamp 1581321262
transform 1 0 3264 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_152
timestamp 1581321262
transform 1 0 1632 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_153
timestamp 1581321262
transform 1 0 0 0 1 5469
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_154
timestamp 1581321262
transform 1 0 9792 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_155
timestamp 1581321262
transform 1 0 8160 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_156
timestamp 1581321262
transform 1 0 6528 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_157
timestamp 1581321262
transform 1 0 4896 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_158
timestamp 1581321262
transform 1 0 3264 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_159
timestamp 1581321262
transform 1 0 1632 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_160
timestamp 1581321262
transform 1 0 0 0 1 5265
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_161
timestamp 1581321262
transform 1 0 9792 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_162
timestamp 1581321262
transform 1 0 8160 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_163
timestamp 1581321262
transform 1 0 6528 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_164
timestamp 1581321262
transform 1 0 4896 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_165
timestamp 1581321262
transform 1 0 3264 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_166
timestamp 1581321262
transform 1 0 1632 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_167
timestamp 1581321262
transform 1 0 0 0 1 5061
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_168
timestamp 1581321262
transform 1 0 9792 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_169
timestamp 1581321262
transform 1 0 8160 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_170
timestamp 1581321262
transform 1 0 6528 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_171
timestamp 1581321262
transform 1 0 4896 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_172
timestamp 1581321262
transform 1 0 3264 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_173
timestamp 1581321262
transform 1 0 1632 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_174
timestamp 1581321262
transform 1 0 0 0 1 4857
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_175
timestamp 1581321262
transform 1 0 9792 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_176
timestamp 1581321262
transform 1 0 8160 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_177
timestamp 1581321262
transform 1 0 6528 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_178
timestamp 1581321262
transform 1 0 4896 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_179
timestamp 1581321262
transform 1 0 3264 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_180
timestamp 1581321262
transform 1 0 1632 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_181
timestamp 1581321262
transform 1 0 0 0 1 4653
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_182
timestamp 1581321262
transform 1 0 9792 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_183
timestamp 1581321262
transform 1 0 8160 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_184
timestamp 1581321262
transform 1 0 6528 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_185
timestamp 1581321262
transform 1 0 4896 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_186
timestamp 1581321262
transform 1 0 3264 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_187
timestamp 1581321262
transform 1 0 1632 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_188
timestamp 1581321262
transform 1 0 0 0 1 4449
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_189
timestamp 1581321262
transform 1 0 9792 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_190
timestamp 1581321262
transform 1 0 8160 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_191
timestamp 1581321262
transform 1 0 6528 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_192
timestamp 1581321262
transform 1 0 4896 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_193
timestamp 1581321262
transform 1 0 3264 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_194
timestamp 1581321262
transform 1 0 1632 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_195
timestamp 1581321262
transform 1 0 0 0 1 4141
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_196
timestamp 1581321262
transform 1 0 9792 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_197
timestamp 1581321262
transform 1 0 8160 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_198
timestamp 1581321262
transform 1 0 6528 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_199
timestamp 1581321262
transform 1 0 4896 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_200
timestamp 1581321262
transform 1 0 3264 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_201
timestamp 1581321262
transform 1 0 1632 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_202
timestamp 1581321262
transform 1 0 0 0 1 3937
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_203
timestamp 1581321262
transform 1 0 9792 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_204
timestamp 1581321262
transform 1 0 8160 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_205
timestamp 1581321262
transform 1 0 6528 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_206
timestamp 1581321262
transform 1 0 4896 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_207
timestamp 1581321262
transform 1 0 3264 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_208
timestamp 1581321262
transform 1 0 1632 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_209
timestamp 1581321262
transform 1 0 0 0 1 3733
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_210
timestamp 1581321262
transform 1 0 9792 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_211
timestamp 1581321262
transform 1 0 8160 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_212
timestamp 1581321262
transform 1 0 6528 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_213
timestamp 1581321262
transform 1 0 4896 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_214
timestamp 1581321262
transform 1 0 3264 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_215
timestamp 1581321262
transform 1 0 1632 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_216
timestamp 1581321262
transform 1 0 0 0 1 3529
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_217
timestamp 1581321262
transform 1 0 9792 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_218
timestamp 1581321262
transform 1 0 8160 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_219
timestamp 1581321262
transform 1 0 6528 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_220
timestamp 1581321262
transform 1 0 4896 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_221
timestamp 1581321262
transform 1 0 3264 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_222
timestamp 1581321262
transform 1 0 1632 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_223
timestamp 1581321262
transform 1 0 0 0 1 3325
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_224
timestamp 1581321262
transform 1 0 9792 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_225
timestamp 1581321262
transform 1 0 8160 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_226
timestamp 1581321262
transform 1 0 6528 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_227
timestamp 1581321262
transform 1 0 4896 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_228
timestamp 1581321262
transform 1 0 3264 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_229
timestamp 1581321262
transform 1 0 1632 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_230
timestamp 1581321262
transform 1 0 0 0 1 3121
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_231
timestamp 1581321262
transform 1 0 9792 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_232
timestamp 1581321262
transform 1 0 8160 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_233
timestamp 1581321262
transform 1 0 6528 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_234
timestamp 1581321262
transform 1 0 4896 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_235
timestamp 1581321262
transform 1 0 3264 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_236
timestamp 1581321262
transform 1 0 1632 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_237
timestamp 1581321262
transform 1 0 0 0 1 2917
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_238
timestamp 1581321262
transform 1 0 9792 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_239
timestamp 1581321262
transform 1 0 8160 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_240
timestamp 1581321262
transform 1 0 6528 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_241
timestamp 1581321262
transform 1 0 4896 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_242
timestamp 1581321262
transform 1 0 3264 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_243
timestamp 1581321262
transform 1 0 1632 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_244
timestamp 1581321262
transform 1 0 0 0 1 2713
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_245
timestamp 1581321262
transform 1 0 9792 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_246
timestamp 1581321262
transform 1 0 8160 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_247
timestamp 1581321262
transform 1 0 6528 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_248
timestamp 1581321262
transform 1 0 4896 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_249
timestamp 1581321262
transform 1 0 3264 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_250
timestamp 1581321262
transform 1 0 1632 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_251
timestamp 1581321262
transform 1 0 0 0 1 2405
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_252
timestamp 1581321262
transform 1 0 9792 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_253
timestamp 1581321262
transform 1 0 8160 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_254
timestamp 1581321262
transform 1 0 6528 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_255
timestamp 1581321262
transform 1 0 4896 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_256
timestamp 1581321262
transform 1 0 3264 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_257
timestamp 1581321262
transform 1 0 1632 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_258
timestamp 1581321262
transform 1 0 0 0 1 2201
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_259
timestamp 1581321262
transform 1 0 9792 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_260
timestamp 1581321262
transform 1 0 8160 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_261
timestamp 1581321262
transform 1 0 6528 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_262
timestamp 1581321262
transform 1 0 4896 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_263
timestamp 1581321262
transform 1 0 3264 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_264
timestamp 1581321262
transform 1 0 1632 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_265
timestamp 1581321262
transform 1 0 0 0 1 1997
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_266
timestamp 1581321262
transform 1 0 9792 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_267
timestamp 1581321262
transform 1 0 8160 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_268
timestamp 1581321262
transform 1 0 6528 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_269
timestamp 1581321262
transform 1 0 4896 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_270
timestamp 1581321262
transform 1 0 3264 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_271
timestamp 1581321262
transform 1 0 1632 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_272
timestamp 1581321262
transform 1 0 0 0 1 1793
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_273
timestamp 1581321262
transform 1 0 9792 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_274
timestamp 1581321262
transform 1 0 8160 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_275
timestamp 1581321262
transform 1 0 6528 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_276
timestamp 1581321262
transform 1 0 4896 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_277
timestamp 1581321262
transform 1 0 3264 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_278
timestamp 1581321262
transform 1 0 1632 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_279
timestamp 1581321262
transform 1 0 0 0 1 1589
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_280
timestamp 1581321262
transform 1 0 9792 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_281
timestamp 1581321262
transform 1 0 8160 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_282
timestamp 1581321262
transform 1 0 6528 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_283
timestamp 1581321262
transform 1 0 4896 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_284
timestamp 1581321262
transform 1 0 3264 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_285
timestamp 1581321262
transform 1 0 1632 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_286
timestamp 1581321262
transform 1 0 0 0 1 1385
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_287
timestamp 1581321262
transform 1 0 9792 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_288
timestamp 1581321262
transform 1 0 8160 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_289
timestamp 1581321262
transform 1 0 6528 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_290
timestamp 1581321262
transform 1 0 4896 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_291
timestamp 1581321262
transform 1 0 3264 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_292
timestamp 1581321262
transform 1 0 1632 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_293
timestamp 1581321262
transform 1 0 0 0 1 1181
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_294
timestamp 1581321262
transform 1 0 9792 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_295
timestamp 1581321262
transform 1 0 8160 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_296
timestamp 1581321262
transform 1 0 6528 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_297
timestamp 1581321262
transform 1 0 4896 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_298
timestamp 1581321262
transform 1 0 3264 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_299
timestamp 1581321262
transform 1 0 1632 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_poly_tap  sky130_rom_krom_rom_poly_tap_300
timestamp 1581321262
transform 1 0 0 0 1 977
box 0 17 66 83
use sky130_rom_krom_rom_precharge_array  sky130_rom_krom_rom_precharge_array_0
timestamp 1581321262
transform 1 0 0 0 1 128
box 0 -212 9900 408
<< labels >>
rlabel metal2 s 61 368 89 396 4 precharge
port 3 nsew
rlabel metal2 s 19 1013 47 1041 4 wl_0_0
port 5 nsew
rlabel metal2 s 19 1217 47 1245 4 wl_0_1
port 7 nsew
rlabel metal2 s 19 1421 47 1449 4 wl_0_2
port 9 nsew
rlabel metal2 s 19 1625 47 1653 4 wl_0_3
port 11 nsew
rlabel metal2 s 19 1829 47 1857 4 wl_0_4
port 13 nsew
rlabel metal2 s 19 2033 47 2061 4 wl_0_5
port 15 nsew
rlabel metal2 s 19 2237 47 2265 4 wl_0_6
port 17 nsew
rlabel metal2 s 19 2441 47 2469 4 wl_0_7
port 19 nsew
rlabel metal2 s 19 2749 47 2777 4 wl_0_8
port 21 nsew
rlabel metal2 s 19 2953 47 2981 4 wl_0_9
port 23 nsew
rlabel metal2 s 19 3157 47 3185 4 wl_0_10
port 25 nsew
rlabel metal2 s 19 3361 47 3389 4 wl_0_11
port 27 nsew
rlabel metal2 s 19 3565 47 3593 4 wl_0_12
port 29 nsew
rlabel metal2 s 19 3769 47 3797 4 wl_0_13
port 31 nsew
rlabel metal2 s 19 3973 47 4001 4 wl_0_14
port 33 nsew
rlabel metal2 s 19 4177 47 4205 4 wl_0_15
port 35 nsew
rlabel metal2 s 19 4485 47 4513 4 wl_0_16
port 37 nsew
rlabel metal2 s 19 4689 47 4717 4 wl_0_17
port 39 nsew
rlabel metal2 s 19 4893 47 4921 4 wl_0_18
port 41 nsew
rlabel metal2 s 19 5097 47 5125 4 wl_0_19
port 43 nsew
rlabel metal2 s 19 5301 47 5329 4 wl_0_20
port 45 nsew
rlabel metal2 s 19 5505 47 5533 4 wl_0_21
port 47 nsew
rlabel metal2 s 19 5709 47 5737 4 wl_0_22
port 49 nsew
rlabel metal2 s 19 5913 47 5941 4 wl_0_23
port 51 nsew
rlabel metal2 s 19 6221 47 6249 4 wl_0_24
port 53 nsew
rlabel metal2 s 19 6425 47 6453 4 wl_0_25
port 55 nsew
rlabel metal2 s 19 6629 47 6657 4 wl_0_26
port 57 nsew
rlabel metal2 s 19 6833 47 6861 4 wl_0_27
port 59 nsew
rlabel metal2 s 19 7037 47 7065 4 wl_0_28
port 61 nsew
rlabel metal2 s 19 7241 47 7269 4 wl_0_29
port 63 nsew
rlabel metal2 s 19 7445 47 7473 4 wl_0_30
port 65 nsew
rlabel metal2 s 19 7649 47 7677 4 wl_0_31
port 67 nsew
rlabel metal2 s 19 7957 47 7985 4 wl_0_32
port 69 nsew
rlabel metal2 s 19 8161 47 8189 4 wl_0_33
port 71 nsew
rlabel metal2 s 19 8365 47 8393 4 wl_0_34
port 73 nsew
rlabel metal2 s 19 8569 47 8597 4 wl_0_35
port 75 nsew
rlabel metal2 s 19 8773 47 8801 4 wl_0_36
port 77 nsew
rlabel metal2 s 19 8977 47 9005 4 wl_0_37
port 79 nsew
rlabel metal2 s 19 9181 47 9209 4 wl_0_38
port 81 nsew
rlabel metal2 s 19 9385 47 9413 4 wl_0_39
port 83 nsew
rlabel metal2 s 19 9693 47 9721 4 wl_0_40
port 85 nsew
rlabel metal2 s 19 9897 47 9925 4 wl_0_41
port 87 nsew
rlabel metal1 s 128 -14 156 14 4 bl_0_0
port 89 nsew
rlabel metal1 s 332 -14 360 14 4 bl_0_1
port 91 nsew
rlabel metal1 s 536 -14 564 14 4 bl_0_2
port 93 nsew
rlabel metal1 s 740 -14 768 14 4 bl_0_3
port 95 nsew
rlabel metal1 s 944 -14 972 14 4 bl_0_4
port 97 nsew
rlabel metal1 s 1148 -14 1176 14 4 bl_0_5
port 99 nsew
rlabel metal1 s 1352 -14 1380 14 4 bl_0_6
port 101 nsew
rlabel metal1 s 1556 -14 1584 14 4 bl_0_7
port 103 nsew
rlabel metal1 s 1760 -14 1788 14 4 bl_0_8
port 105 nsew
rlabel metal1 s 1964 -14 1992 14 4 bl_0_9
port 107 nsew
rlabel metal1 s 2168 -14 2196 14 4 bl_0_10
port 109 nsew
rlabel metal1 s 2372 -14 2400 14 4 bl_0_11
port 111 nsew
rlabel metal1 s 2576 -14 2604 14 4 bl_0_12
port 113 nsew
rlabel metal1 s 2780 -14 2808 14 4 bl_0_13
port 115 nsew
rlabel metal1 s 2984 -14 3012 14 4 bl_0_14
port 117 nsew
rlabel metal1 s 3188 -14 3216 14 4 bl_0_15
port 119 nsew
rlabel metal1 s 3392 -14 3420 14 4 bl_0_16
port 121 nsew
rlabel metal1 s 3596 -14 3624 14 4 bl_0_17
port 123 nsew
rlabel metal1 s 3800 -14 3828 14 4 bl_0_18
port 125 nsew
rlabel metal1 s 4004 -14 4032 14 4 bl_0_19
port 127 nsew
rlabel metal1 s 4208 -14 4236 14 4 bl_0_20
port 129 nsew
rlabel metal1 s 4412 -14 4440 14 4 bl_0_21
port 131 nsew
rlabel metal1 s 4616 -14 4644 14 4 bl_0_22
port 133 nsew
rlabel metal1 s 4820 -14 4848 14 4 bl_0_23
port 135 nsew
rlabel metal1 s 5024 -14 5052 14 4 bl_0_24
port 137 nsew
rlabel metal1 s 5228 -14 5256 14 4 bl_0_25
port 139 nsew
rlabel metal1 s 5432 -14 5460 14 4 bl_0_26
port 141 nsew
rlabel metal1 s 5636 -14 5664 14 4 bl_0_27
port 143 nsew
rlabel metal1 s 5840 -14 5868 14 4 bl_0_28
port 145 nsew
rlabel metal1 s 6044 -14 6072 14 4 bl_0_29
port 147 nsew
rlabel metal1 s 6248 -14 6276 14 4 bl_0_30
port 149 nsew
rlabel metal1 s 6452 -14 6480 14 4 bl_0_31
port 151 nsew
rlabel metal1 s 6656 -14 6684 14 4 bl_0_32
port 153 nsew
rlabel metal1 s 6860 -14 6888 14 4 bl_0_33
port 155 nsew
rlabel metal1 s 7064 -14 7092 14 4 bl_0_34
port 157 nsew
rlabel metal1 s 7268 -14 7296 14 4 bl_0_35
port 159 nsew
rlabel metal1 s 7472 -14 7500 14 4 bl_0_36
port 161 nsew
rlabel metal1 s 7676 -14 7704 14 4 bl_0_37
port 163 nsew
rlabel metal1 s 7880 -14 7908 14 4 bl_0_38
port 165 nsew
rlabel metal1 s 8084 -14 8112 14 4 bl_0_39
port 167 nsew
rlabel metal1 s 8288 -14 8316 14 4 bl_0_40
port 169 nsew
rlabel metal1 s 8492 -14 8520 14 4 bl_0_41
port 171 nsew
rlabel metal1 s 8696 -14 8724 14 4 bl_0_42
port 173 nsew
rlabel metal1 s 8900 -14 8928 14 4 bl_0_43
port 175 nsew
rlabel metal1 s 9104 -14 9132 14 4 bl_0_44
port 177 nsew
rlabel metal1 s 9308 -14 9336 14 4 bl_0_45
port 179 nsew
rlabel metal1 s 9512 -14 9540 14 4 bl_0_46
port 181 nsew
rlabel metal1 s 9716 -14 9744 14 4 bl_0_47
port 183 nsew
rlabel metal1 s 10013 368 10041 396 4 precharge_r
port 185 nsew
rlabel metal2 s 230 7803 9860 7831 4 gnd
port 187 nsew
rlabel metal2 s 230 4331 9860 4359 4 gnd
port 187 nsew
rlabel metal1 s 114 10228 142 10256 4 gnd
port 187 nsew
rlabel metal2 s 230 859 9860 887 4 gnd
port 187 nsew
rlabel metal2 s 230 6067 9860 6095 4 gnd
port 187 nsew
rlabel metal1 s 9730 10228 9758 10256 4 gnd
port 187 nsew
rlabel metal2 s 230 9539 9860 9567 4 gnd
port 187 nsew
rlabel metal2 s 230 2595 9860 2623 4 gnd
port 187 nsew
rlabel metal2 s 12 -32 40 32 4 vdd
port 189 nsew
<< properties >>
string FIXED_BBOX 0 0 10041 974
<< end >>
