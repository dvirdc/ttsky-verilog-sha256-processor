VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_rom_1kbyte
   CLASS BLOCK ;
   SIZE 175.13 BY 122.55 ;
   SYMMETRY X Y R90 ;
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 8.51 -7.1 8.89 ;
      END
   END clk0
   PIN cs0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  15.265 -7.48 15.645 -7.1 ;
      END
   END cs0
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  24.83 -7.48 25.21 -7.1 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  26.87 -7.48 27.25 -7.1 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  28.91 -7.48 29.29 -7.1 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  30.205 -7.48 30.585 -7.1 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 35.7 -7.1 36.08 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 36.445 -7.1 36.825 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 37.135 -7.1 37.515 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 34.23 -7.1 34.61 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 37.825 -7.1 38.205 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 33.54 -7.1 33.92 ;
      END
   END addr0[9]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  51.675 -7.48 52.055 -7.1 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  53.215 -7.48 53.595 -7.1 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  54.755 -7.48 55.135 -7.1 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  56.295 -7.48 56.675 -7.1 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  57.835 -7.48 58.215 -7.1 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  59.375 -7.48 59.755 -7.1 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  60.915 -7.48 61.295 -7.1 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  62.455 -7.48 62.835 -7.1 ;
      END
   END dout0[7]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  180.87 -7.48 182.61 130.03 ;
         LAYER met3 ;
         RECT  -7.48 128.29 182.61 130.03 ;
         LAYER met4 ;
         RECT  -7.48 -7.48 -5.74 130.03 ;
         LAYER met3 ;
         RECT  -7.48 -7.48 182.61 -5.74 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  177.39 -4.0 179.13 126.55 ;
         LAYER met4 ;
         RECT  -4.0 -4.0 -2.26 126.55 ;
         LAYER met3 ;
         RECT  -4.0 124.81 179.13 126.55 ;
         LAYER met3 ;
         RECT  -4.0 -4.0 179.13 -2.26 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 174.51 121.93 ;
   LAYER  met2 ;
      RECT  0.62 0.62 174.51 121.93 ;
   LAYER  met3 ;
      RECT  0.62 0.62 174.51 121.93 ;
   LAYER  met4 ;
      RECT  0.62 0.62 174.51 121.93 ;
   END
END    sky130_rom_1kbyte
END    LIBRARY
